module HasDeadCode(
  input   i,
  output  o
);
  assign o = i;
endmodule
