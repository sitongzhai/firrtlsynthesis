module Console(
    input clock,
    input reset,
    input io_toggle,
    output [7:0] io_character,
    output [7:0] io_characterAvailable
);
    wire [7:0] helloWorld_0;
    wire [7:0] helloWorld_1;
    wire [7:0] helloWorld_2;
    wire [7:0] helloWorld_3;
    wire [7:0] helloWorld_4;
    wire [7:0] helloWorld_5;
    wire [7:0] helloWorld_6;
    wire [7:0] helloWorld_7;
    wire [7:0] helloWorld_8;
    wire [7:0] helloWorld_9;
    wire [7:0] helloWorld_10;
    wire [7:0] helloWorld_11;
    wire [7:0] helloWorld_12;
    wire [7:0] helloWorld_13;
    wire [7:0] helloWorld_14;
    wire [7:0] helloWorld_15;
    wire [7:0] helloWorld_16;
    wire [7:0] helloWorld_17;
    wire [7:0] helloWorld_18;
    wire [7:0] helloWorld_19;
    wire [7:0] helloWorld_20;
    wire [7:0] helloWorld_21;
    wire [7:0] helloWorld_22;
    wire [7:0] helloWorld_23;
    wire [7:0] helloWorld_24;
    wire [7:0] helloWorld_25;
    wire [7:0] helloWorld_26;
    wire [7:0] helloWorld_27;
    wire [7:0] helloWorld_28;
    wire [7:0] helloWorld_29;
    wire [7:0] helloWorld_30;
    wire [7:0] helloWorld_31;
    wire [7:0] helloWorld_32;
    wire [7:0] helloWorld_33;
    wire [7:0] helloWorld_34;
    wire [7:0] helloWorld_35;
    wire [7:0] helloWorld_36;
    wire [7:0] helloWorld_37;
    wire [7:0] helloWorld_38;
    wire [7:0] helloWorld_39;
    wire [7:0] helloWorld_40;
    wire [7:0] helloWorld_41;
    wire [7:0] helloWorld_42;
    wire [7:0] helloWorld_43;
    wire [7:0] helloWorld_44;
    wire [7:0] helloWorld_45;
    wire [7:0] helloWorld_46;
    wire [7:0] helloWorld_47;
    wire [7:0] helloWorld_48;
    wire [7:0] helloWorld_49;
    wire [7:0] helloWorld_50;
    wire [7:0] helloWorld_51;
    wire [7:0] helloWorld_52;
    wire [7:0] helloWorld_53;
    wire [7:0] helloWorld_54;
    wire [7:0] helloWorld_55;
    wire [7:0] helloWorld_56;
    wire [7:0] helloWorld_57;
    wire [7:0] helloWorld_58;
    wire [7:0] helloWorld_59;
    wire [7:0] helloWorld_60;
    wire [7:0] helloWorld_61;
    wire [7:0] helloWorld_62;
    wire [7:0] helloWorld_63;
    wire [7:0] helloWorld_64;
    wire [7:0] helloWorld_65;
    wire [7:0] helloWorld_66;
    wire [7:0] helloWorld_67;
    wire [7:0] helloWorld_68;
    wire [7:0] helloWorld_69;
    wire [7:0] helloWorld_70;
    wire [7:0] helloWorld_71;
    wire [7:0] helloWorld_72;
    wire [7:0] helloWorld_73;
    wire [7:0] helloWorld_74;
    wire [7:0] helloWorld_75;
    wire [7:0] helloWorld_76;
    wire [7:0] helloWorld_77;
    wire [7:0] helloWorld_78;
    wire [7:0] helloWorld_79;
    wire [7:0] helloWorld_80;
    wire [7:0] helloWorld_81;
    wire [7:0] helloWorld_82;
    wire [7:0] helloWorld_83;
    wire [7:0] helloWorld_84;
    wire [7:0] helloWorld_85;
    wire [7:0] helloWorld_86;
    wire [7:0] helloWorld_87;
    wire [7:0] helloWorld_88;
    wire [7:0] helloWorld_89;
    wire [7:0] helloWorld_90;
    wire [7:0] helloWorld_91;
    wire [7:0] helloWorld_92;
    wire [7:0] helloWorld_93;
    wire [7:0] helloWorld_94;
    wire [7:0] helloWorld_95;
    wire [7:0] helloWorld_96;
    wire [7:0] helloWorld_97;
    wire [7:0] helloWorld_98;
    wire [7:0] helloWorld_99;
    wire [7:0] helloWorld_100;
    wire [7:0] helloWorld_101;
    wire [7:0] helloWorld_102;
    wire [7:0] helloWorld_103;
    wire [7:0] helloWorld_104;
    wire [7:0] helloWorld_105;
    wire [7:0] helloWorld_106;
    wire [7:0] helloWorld_107;
    wire [7:0] helloWorld_108;
    wire [7:0] helloWorld_109;
    wire [7:0] helloWorld_110;
    wire [7:0] helloWorld_111;
    wire [7:0] helloWorld_112;
    wire [7:0] helloWorld_113;
    wire [7:0] helloWorld_114;
    wire [7:0] helloWorld_115;
    wire [7:0] helloWorld_116;
    wire [7:0] helloWorld_117;
    wire [7:0] helloWorld_118;
    wire [7:0] helloWorld_119;
    wire [7:0] helloWorld_120;
    wire [7:0] helloWorld_121;
    wire [7:0] helloWorld_122;
    wire [7:0] helloWorld_123;
    wire [7:0] helloWorld_124;
    wire [7:0] helloWorld_125;
    wire [7:0] helloWorld_126;
    wire [7:0] helloWorld_127;
    wire [7:0] helloWorld_128;
    wire [7:0] helloWorld_129;
    wire [7:0] helloWorld_130;
    wire [7:0] helloWorld_131;
    wire [7:0] helloWorld_132;
    wire [7:0] helloWorld_133;
    wire [7:0] helloWorld_134;
    wire [7:0] helloWorld_135;
    wire [7:0] helloWorld_136;
    wire [7:0] helloWorld_137;
    wire [7:0] helloWorld_138;
    wire [7:0] helloWorld_139;
    wire [7:0] helloWorld_140;
    wire [7:0] helloWorld_141;
    wire [7:0] helloWorld_142;
    wire [7:0] helloWorld_143;
    wire [7:0] helloWorld_144;
    wire [7:0] helloWorld_145;
    wire [7:0] helloWorld_146;
    wire [7:0] helloWorld_147;
    wire [7:0] helloWorld_148;
    wire [7:0] helloWorld_149;
    wire [7:0] helloWorld_150;
    wire [7:0] helloWorld_151;
    wire [7:0] helloWorld_152;
    wire [7:0] helloWorld_153;
    wire [7:0] helloWorld_154;
    wire [7:0] helloWorld_155;
    wire [7:0] helloWorld_156;
    wire [7:0] helloWorld_157;
    wire [7:0] helloWorld_158;
    wire [7:0] helloWorld_159;
    wire [7:0] helloWorld_160;
    wire [7:0] helloWorld_161;
    wire [7:0] helloWorld_162;
    wire [7:0] helloWorld_163;
    wire [7:0] helloWorld_164;
    wire [7:0] helloWorld_165;
    wire [7:0] helloWorld_166;
    wire [7:0] helloWorld_167;
    wire [7:0] helloWorld_168;
    wire [7:0] helloWorld_169;
    wire [7:0] helloWorld_170;
    wire [7:0] helloWorld_171;
    wire [7:0] helloWorld_172;
    wire [7:0] helloWorld_173;
    wire [7:0] helloWorld_174;
    wire [7:0] helloWorld_175;
    wire [7:0] helloWorld_176;
    wire [7:0] helloWorld_177;
    wire [7:0] helloWorld_178;
    wire [7:0] helloWorld_179;
    wire [7:0] helloWorld_180;
    wire [7:0] helloWorld_181;
    wire [7:0] helloWorld_182;
    wire [7:0] helloWorld_183;
    wire [7:0] helloWorld_184;
    wire [7:0] helloWorld_185;
    wire [7:0] helloWorld_186;
    wire [7:0] helloWorld_187;
    wire [7:0] helloWorld_188;
    wire [7:0] helloWorld_189;
    wire [7:0] helloWorld_190;
    wire [7:0] helloWorld_191;
    wire [7:0] helloWorld_192;
    wire [7:0] helloWorld_193;
    wire [7:0] helloWorld_194;
    wire [7:0] helloWorld_195;
    wire [7:0] helloWorld_196;
    wire [7:0] helloWorld_197;
    wire [7:0] helloWorld_198;
    wire [7:0] helloWorld_199;
    wire [7:0] helloWorld_200;
    wire [7:0] helloWorld_201;
    wire [7:0] helloWorld_202;
    wire [7:0] helloWorld_203;
    wire [7:0] helloWorld_204;
    wire [7:0] helloWorld_205;
    wire [7:0] helloWorld_206;
    wire [7:0] helloWorld_207;
    wire [7:0] helloWorld_208;
    wire [7:0] helloWorld_209;
    wire [7:0] helloWorld_210;
    wire [7:0] helloWorld_211;
    wire [7:0] helloWorld_212;
    wire [7:0] helloWorld_213;
    wire [7:0] helloWorld_214;
    wire [7:0] helloWorld_215;
    wire [7:0] helloWorld_216;
    wire [7:0] helloWorld_217;
    wire [7:0] helloWorld_218;
    wire [7:0] helloWorld_219;
    wire [7:0] helloWorld_220;
    wire [7:0] helloWorld_221;
    wire [7:0] helloWorld_222;
    wire [7:0] helloWorld_223;
    wire [7:0] helloWorld_224;
    wire [7:0] helloWorld_225;
    wire [7:0] helloWorld_226;
    wire [7:0] helloWorld_227;
    wire [7:0] helloWorld_228;
    wire [7:0] helloWorld_229;
    wire [7:0] helloWorld_230;
    wire [7:0] helloWorld_231;
    wire [7:0] helloWorld_232;
    wire [7:0] helloWorld_233;
    wire [7:0] helloWorld_234;
    wire [7:0] helloWorld_235;
    wire [7:0] helloWorld_236;
    wire [7:0] helloWorld_237;
    wire [7:0] helloWorld_238;
    wire [7:0] helloWorld_239;
    wire [7:0] helloWorld_240;
    wire [7:0] helloWorld_241;
    wire [7:0] helloWorld_242;
    wire [7:0] helloWorld_243;
    wire [7:0] helloWorld_244;
    wire [7:0] helloWorld_245;
    wire [7:0] helloWorld_246;
    wire [7:0] helloWorld_247;
    wire [7:0] helloWorld_248;
    wire [7:0] helloWorld_249;
    wire [7:0] helloWorld_250;
    wire [7:0] helloWorld_251;
    wire [7:0] helloWorld_252;
    wire [7:0] helloWorld_253;
    wire [7:0] helloWorld_254;
    wire [7:0] helloWorld_255;
    wire [7:0] helloWorld_256;
    wire [7:0] helloWorld_257;
    wire [7:0] helloWorld_258;
    wire [7:0] helloWorld_259;
    wire [7:0] helloWorld_260;
    wire [7:0] helloWorld_261;
    wire [7:0] helloWorld_262;
    wire [7:0] helloWorld_263;
    wire [7:0] helloWorld_264;
    wire [7:0] helloWorld_265;
    wire [7:0] helloWorld_266;
    wire [7:0] helloWorld_267;
    wire [7:0] helloWorld_268;
    wire [7:0] helloWorld_269;
    wire [7:0] helloWorld_270;
    wire [7:0] helloWorld_271;
    wire [7:0] helloWorld_272;
    wire [7:0] helloWorld_273;
    wire [7:0] helloWorld_274;
    wire [7:0] helloWorld_275;
    wire [7:0] helloWorld_276;
    wire [7:0] helloWorld_277;
    wire [7:0] helloWorld_278;
    wire [7:0] helloWorld_279;
    wire [7:0] helloWorld_280;
    wire [7:0] helloWorld_281;
    wire [7:0] helloWorld_282;
    wire [7:0] helloWorld_283;
    wire [7:0] helloWorld_284;
    wire [7:0] helloWorld_285;
    wire [7:0] helloWorld_286;
    wire [7:0] helloWorld_287;
    wire [7:0] helloWorld_288;
    wire [7:0] helloWorld_289;
    wire [7:0] helloWorld_290;
    wire [7:0] helloWorld_291;
    wire [7:0] helloWorld_292;
    wire [7:0] helloWorld_293;
    wire [7:0] helloWorld_294;
    wire [7:0] helloWorld_295;
    wire [7:0] helloWorld_296;
    wire [7:0] helloWorld_297;
    wire [7:0] helloWorld_298;
    wire [7:0] helloWorld_299;
    wire [7:0] helloWorld_300;
    wire [7:0] helloWorld_301;
    wire [7:0] helloWorld_302;
    wire [7:0] helloWorld_303;
    wire [7:0] helloWorld_304;
    wire [7:0] helloWorld_305;
    wire [7:0] helloWorld_306;
    wire [7:0] helloWorld_307;
    wire [7:0] helloWorld_308;
    wire [7:0] helloWorld_309;
    wire [7:0] helloWorld_310;
    wire [7:0] helloWorld_311;
    wire [7:0] helloWorld_312;
    wire [7:0] helloWorld_313;
    wire [7:0] helloWorld_314;
    wire [7:0] helloWorld_315;
    wire [7:0] helloWorld_316;
    wire [7:0] helloWorld_317;
    wire [7:0] helloWorld_318;
    wire [7:0] helloWorld_319;
    wire [7:0] helloWorld_320;
    wire [7:0] helloWorld_321;
    wire [7:0] helloWorld_322;
    wire [7:0] helloWorld_323;
    wire [7:0] helloWorld_324;
    wire [7:0] helloWorld_325;
    wire [7:0] helloWorld_326;
    wire [7:0] helloWorld_327;
    wire [7:0] helloWorld_328;
    wire [7:0] helloWorld_329;
    wire [7:0] helloWorld_330;
    wire [7:0] helloWorld_331;
    wire [7:0] helloWorld_332;
    wire [7:0] helloWorld_333;
    wire [7:0] helloWorld_334;
    wire [7:0] helloWorld_335;
    wire [7:0] helloWorld_336;
    wire [7:0] helloWorld_337;
    wire [7:0] helloWorld_338;
    wire [7:0] helloWorld_339;
    wire [7:0] helloWorld_340;
    wire [7:0] helloWorld_341;
    wire [7:0] helloWorld_342;
    wire [7:0] helloWorld_343;
    wire [7:0] helloWorld_344;
    wire [7:0] helloWorld_345;
    wire [7:0] helloWorld_346;
    wire [7:0] helloWorld_347;
    wire [7:0] helloWorld_348;
    wire [7:0] helloWorld_349;
    wire [7:0] helloWorld_350;
    wire [7:0] helloWorld_351;
    wire [7:0] helloWorld_352;
    wire [7:0] helloWorld_353;
    wire [7:0] helloWorld_354;
    wire [7:0] helloWorld_355;
    wire [7:0] helloWorld_356;
    wire [7:0] helloWorld_357;
    wire [7:0] helloWorld_358;
    wire [7:0] helloWorld_359;
    wire [7:0] helloWorld_360;
    wire [7:0] helloWorld_361;
    wire [7:0] helloWorld_362;
    wire [7:0] helloWorld_363;
    wire [7:0] helloWorld_364;
    wire [7:0] helloWorld_365;
    wire [7:0] helloWorld_366;
    wire [7:0] helloWorld_367;
    wire [7:0] helloWorld_368;
    wire [7:0] helloWorld_369;
    wire [7:0] helloWorld_370;
    wire [7:0] helloWorld_371;
    wire [7:0] helloWorld_372;
    wire [7:0] helloWorld_373;
    wire [7:0] helloWorld_374;
    wire [7:0] helloWorld_375;
    wire [7:0] helloWorld_376;
    wire [7:0] helloWorld_377;
    wire [7:0] helloWorld_378;
    wire [7:0] helloWorld_379;
    wire [7:0] helloWorld_380;
    wire [7:0] helloWorld_381;
    wire [7:0] helloWorld_382;
    wire [7:0] helloWorld_383;
    wire [7:0] helloWorld_384;
    wire [7:0] helloWorld_385;
    wire [7:0] helloWorld_386;
    wire [7:0] helloWorld_387;
    wire [8:0] _pointer__q;
    wire [8:0] _pointer__d;
    DFF_POSCLK #(.width(9)) pointer (
        .q(_pointer__q),
        .d(_pointer__d),
        .clk(clock)
    );
    wire [8:0] _arrivedPointer__q;
    wire [8:0] _arrivedPointer__d;
    DFF_POSCLK #(.width(9)) arrivedPointer (
        .q(_arrivedPointer__q),
        .d(_arrivedPointer__d),
        .clk(clock)
    );
    wire _lastToggle__q;
    wire _lastToggle__d;
    DFF_POSCLK #(.width(1)) lastToggle (
        .q(_lastToggle__q),
        .d(_lastToggle__d),
        .clk(clock)
    );
    wire _characterArrived__q;
    wire _characterArrived__d;
    DFF_POSCLK #(.width(1)) characterArrived (
        .q(_characterArrived__q),
        .d(_characterArrived__d),
        .clk(clock)
    );
    wire gotToggle;
    NEQ_UNSIGNED #(.width(1)) u_neq_1 (
        .y(gotToggle),
        .a(io_toggle),
        .b(_lastToggle__q)
    );
    wire [9:0] _T_796;
    assign _T_796 = 10'h183;
    wire [9:0] _T_797;
    assign _T_797 = 10'h183;
    wire [8:0] _T_798;
    assign _T_798 = 9'h183;
    wire _T_799;
    EQ_UNSIGNED #(.width(9)) u_eq_2 (
        .y(_T_799),
        .a(_pointer__q),
        .b(_T_798)
    );
    wire [9:0] _T_802;
    wire [8:0] _WTEMP_0;
    PAD_UNSIGNED #(.width(1), .n(9)) u_pad_3 (
        .y(_WTEMP_0),
        .in(1'h1)
    );
    ADD_UNSIGNED #(.width(9)) u_add_4 (
        .y(_T_802),
        .a(_pointer__q),
        .b(_WTEMP_0)
    );
    wire [8:0] _T_803;
    TAIL #(.width(10), .n(1)) tail_5 (
        .y(_T_803),
        .in(_T_802)
    );
    wire [8:0] _T_804;
    wire [8:0] _WTEMP_1;
    PAD_UNSIGNED #(.width(1), .n(9)) u_pad_6 (
        .y(_WTEMP_1),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(9)) u_mux_7 (
        .y(_T_804),
        .sel(_T_799),
        .a(_WTEMP_1),
        .b(_T_803)
    );
    wire _GEN_1;
    MUX_UNSIGNED #(.width(1)) u_mux_8 (
        .y(_GEN_1),
        .sel(gotToggle),
        .a(io_toggle),
        .b(_lastToggle__q)
    );
    wire _GEN_2;
    MUX_UNSIGNED #(.width(1)) u_mux_9 (
        .y(_GEN_2),
        .sel(gotToggle),
        .a(1'h0),
        .b(_characterArrived__q)
    );
    wire [8:0] _GEN_3;
    MUX_UNSIGNED #(.width(9)) u_mux_10 (
        .y(_GEN_3),
        .sel(gotToggle),
        .a(_T_804),
        .b(_pointer__q)
    );
    wire [8:0] _GEN_4;
    MUX_UNSIGNED #(.width(9)) u_mux_11 (
        .y(_GEN_4),
        .sel(gotToggle),
        .a(_pointer__q),
        .b(_arrivedPointer__q)
    );
    wire __T_807__q;
    wire __T_807__d;
    DFF_POSCLK #(.width(1)) _T_807 (
        .q(__T_807__q),
        .d(__T_807__d),
        .clk(clock)
    );
    wire _GEN_5;
    assign _GEN_5 = gotToggle;
    wire __T_809__q;
    wire __T_809__d;
    DFF_POSCLK #(.width(1)) _T_809 (
        .q(__T_809__q),
        .d(__T_809__d),
        .clk(clock)
    );
    wire _GEN_6;
    assign _GEN_6 = __T_807__q;
    wire __T_811__q;
    wire __T_811__d;
    DFF_POSCLK #(.width(1)) _T_811 (
        .q(__T_811__q),
        .d(__T_811__d),
        .clk(clock)
    );
    wire _GEN_7;
    assign _GEN_7 = __T_809__q;
    wire __T_813__q;
    wire __T_813__d;
    DFF_POSCLK #(.width(1)) _T_813 (
        .q(__T_813__q),
        .d(__T_813__d),
        .clk(clock)
    );
    wire _GEN_8;
    assign _GEN_8 = __T_811__q;
    wire __T_815__q;
    wire __T_815__d;
    DFF_POSCLK #(.width(1)) _T_815 (
        .q(__T_815__q),
        .d(__T_815__d),
        .clk(clock)
    );
    wire _GEN_9;
    assign _GEN_9 = __T_813__q;
    wire _GEN_10;
    MUX_UNSIGNED #(.width(1)) u_mux_12 (
        .y(_GEN_10),
        .sel(__T_815__q),
        .a(1'h1),
        .b(_GEN_2)
    );
    wire [7:0] _GEN_0;
    wire _node_0;
    wire [8:0] _WTEMP_2;
    PAD_UNSIGNED #(.width(1), .n(9)) u_pad_13 (
        .y(_WTEMP_2),
        .in(1'h1)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_14 (
        .y(_node_0),
        .a(_WTEMP_2),
        .b(_arrivedPointer__q)
    );
    wire _node_1;
    BITWISEAND #(.width(1)) bitwiseand_15 (
        .y(_node_1),
        .a(1'h1),
        .b(_node_0)
    );
    wire [7:0] _GEN_11;
    MUX_UNSIGNED #(.width(8)) u_mux_16 (
        .y(_GEN_11),
        .sel(_node_1),
        .a(helloWorld_1),
        .b(helloWorld_0)
    );
    wire _node_2;
    wire [8:0] _WTEMP_3;
    PAD_UNSIGNED #(.width(2), .n(9)) u_pad_17 (
        .y(_WTEMP_3),
        .in(2'h2)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_18 (
        .y(_node_2),
        .a(_WTEMP_3),
        .b(_arrivedPointer__q)
    );
    wire _node_3;
    BITWISEAND #(.width(1)) bitwiseand_19 (
        .y(_node_3),
        .a(1'h1),
        .b(_node_2)
    );
    wire [7:0] _GEN_12;
    MUX_UNSIGNED #(.width(8)) u_mux_20 (
        .y(_GEN_12),
        .sel(_node_3),
        .a(helloWorld_2),
        .b(_GEN_11)
    );
    wire _node_4;
    wire [8:0] _WTEMP_4;
    PAD_UNSIGNED #(.width(2), .n(9)) u_pad_21 (
        .y(_WTEMP_4),
        .in(2'h3)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_22 (
        .y(_node_4),
        .a(_WTEMP_4),
        .b(_arrivedPointer__q)
    );
    wire _node_5;
    BITWISEAND #(.width(1)) bitwiseand_23 (
        .y(_node_5),
        .a(1'h1),
        .b(_node_4)
    );
    wire [7:0] _GEN_13;
    MUX_UNSIGNED #(.width(8)) u_mux_24 (
        .y(_GEN_13),
        .sel(_node_5),
        .a(helloWorld_3),
        .b(_GEN_12)
    );
    wire _node_6;
    wire [8:0] _WTEMP_5;
    PAD_UNSIGNED #(.width(3), .n(9)) u_pad_25 (
        .y(_WTEMP_5),
        .in(3'h4)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_26 (
        .y(_node_6),
        .a(_WTEMP_5),
        .b(_arrivedPointer__q)
    );
    wire _node_7;
    BITWISEAND #(.width(1)) bitwiseand_27 (
        .y(_node_7),
        .a(1'h1),
        .b(_node_6)
    );
    wire [7:0] _GEN_14;
    MUX_UNSIGNED #(.width(8)) u_mux_28 (
        .y(_GEN_14),
        .sel(_node_7),
        .a(helloWorld_4),
        .b(_GEN_13)
    );
    wire _node_8;
    wire [8:0] _WTEMP_6;
    PAD_UNSIGNED #(.width(3), .n(9)) u_pad_29 (
        .y(_WTEMP_6),
        .in(3'h5)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_30 (
        .y(_node_8),
        .a(_WTEMP_6),
        .b(_arrivedPointer__q)
    );
    wire _node_9;
    BITWISEAND #(.width(1)) bitwiseand_31 (
        .y(_node_9),
        .a(1'h1),
        .b(_node_8)
    );
    wire [7:0] _GEN_15;
    MUX_UNSIGNED #(.width(8)) u_mux_32 (
        .y(_GEN_15),
        .sel(_node_9),
        .a(helloWorld_5),
        .b(_GEN_14)
    );
    wire _node_10;
    wire [8:0] _WTEMP_7;
    PAD_UNSIGNED #(.width(3), .n(9)) u_pad_33 (
        .y(_WTEMP_7),
        .in(3'h6)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_34 (
        .y(_node_10),
        .a(_WTEMP_7),
        .b(_arrivedPointer__q)
    );
    wire _node_11;
    BITWISEAND #(.width(1)) bitwiseand_35 (
        .y(_node_11),
        .a(1'h1),
        .b(_node_10)
    );
    wire [7:0] _GEN_16;
    MUX_UNSIGNED #(.width(8)) u_mux_36 (
        .y(_GEN_16),
        .sel(_node_11),
        .a(helloWorld_6),
        .b(_GEN_15)
    );
    wire _node_12;
    wire [8:0] _WTEMP_8;
    PAD_UNSIGNED #(.width(3), .n(9)) u_pad_37 (
        .y(_WTEMP_8),
        .in(3'h7)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_38 (
        .y(_node_12),
        .a(_WTEMP_8),
        .b(_arrivedPointer__q)
    );
    wire _node_13;
    BITWISEAND #(.width(1)) bitwiseand_39 (
        .y(_node_13),
        .a(1'h1),
        .b(_node_12)
    );
    wire [7:0] _GEN_17;
    MUX_UNSIGNED #(.width(8)) u_mux_40 (
        .y(_GEN_17),
        .sel(_node_13),
        .a(helloWorld_7),
        .b(_GEN_16)
    );
    wire _node_14;
    wire [8:0] _WTEMP_9;
    PAD_UNSIGNED #(.width(4), .n(9)) u_pad_41 (
        .y(_WTEMP_9),
        .in(4'h8)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_42 (
        .y(_node_14),
        .a(_WTEMP_9),
        .b(_arrivedPointer__q)
    );
    wire _node_15;
    BITWISEAND #(.width(1)) bitwiseand_43 (
        .y(_node_15),
        .a(1'h1),
        .b(_node_14)
    );
    wire [7:0] _GEN_18;
    MUX_UNSIGNED #(.width(8)) u_mux_44 (
        .y(_GEN_18),
        .sel(_node_15),
        .a(helloWorld_8),
        .b(_GEN_17)
    );
    wire _node_16;
    wire [8:0] _WTEMP_10;
    PAD_UNSIGNED #(.width(4), .n(9)) u_pad_45 (
        .y(_WTEMP_10),
        .in(4'h9)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_46 (
        .y(_node_16),
        .a(_WTEMP_10),
        .b(_arrivedPointer__q)
    );
    wire _node_17;
    BITWISEAND #(.width(1)) bitwiseand_47 (
        .y(_node_17),
        .a(1'h1),
        .b(_node_16)
    );
    wire [7:0] _GEN_19;
    MUX_UNSIGNED #(.width(8)) u_mux_48 (
        .y(_GEN_19),
        .sel(_node_17),
        .a(helloWorld_9),
        .b(_GEN_18)
    );
    wire _node_18;
    wire [8:0] _WTEMP_11;
    PAD_UNSIGNED #(.width(4), .n(9)) u_pad_49 (
        .y(_WTEMP_11),
        .in(4'hA)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_50 (
        .y(_node_18),
        .a(_WTEMP_11),
        .b(_arrivedPointer__q)
    );
    wire _node_19;
    BITWISEAND #(.width(1)) bitwiseand_51 (
        .y(_node_19),
        .a(1'h1),
        .b(_node_18)
    );
    wire [7:0] _GEN_20;
    MUX_UNSIGNED #(.width(8)) u_mux_52 (
        .y(_GEN_20),
        .sel(_node_19),
        .a(helloWorld_10),
        .b(_GEN_19)
    );
    wire _node_20;
    wire [8:0] _WTEMP_12;
    PAD_UNSIGNED #(.width(4), .n(9)) u_pad_53 (
        .y(_WTEMP_12),
        .in(4'hB)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_54 (
        .y(_node_20),
        .a(_WTEMP_12),
        .b(_arrivedPointer__q)
    );
    wire _node_21;
    BITWISEAND #(.width(1)) bitwiseand_55 (
        .y(_node_21),
        .a(1'h1),
        .b(_node_20)
    );
    wire [7:0] _GEN_21;
    MUX_UNSIGNED #(.width(8)) u_mux_56 (
        .y(_GEN_21),
        .sel(_node_21),
        .a(helloWorld_11),
        .b(_GEN_20)
    );
    wire _node_22;
    wire [8:0] _WTEMP_13;
    PAD_UNSIGNED #(.width(4), .n(9)) u_pad_57 (
        .y(_WTEMP_13),
        .in(4'hC)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_58 (
        .y(_node_22),
        .a(_WTEMP_13),
        .b(_arrivedPointer__q)
    );
    wire _node_23;
    BITWISEAND #(.width(1)) bitwiseand_59 (
        .y(_node_23),
        .a(1'h1),
        .b(_node_22)
    );
    wire [7:0] _GEN_22;
    MUX_UNSIGNED #(.width(8)) u_mux_60 (
        .y(_GEN_22),
        .sel(_node_23),
        .a(helloWorld_12),
        .b(_GEN_21)
    );
    wire _node_24;
    wire [8:0] _WTEMP_14;
    PAD_UNSIGNED #(.width(4), .n(9)) u_pad_61 (
        .y(_WTEMP_14),
        .in(4'hD)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_62 (
        .y(_node_24),
        .a(_WTEMP_14),
        .b(_arrivedPointer__q)
    );
    wire _node_25;
    BITWISEAND #(.width(1)) bitwiseand_63 (
        .y(_node_25),
        .a(1'h1),
        .b(_node_24)
    );
    wire [7:0] _GEN_23;
    MUX_UNSIGNED #(.width(8)) u_mux_64 (
        .y(_GEN_23),
        .sel(_node_25),
        .a(helloWorld_13),
        .b(_GEN_22)
    );
    wire _node_26;
    wire [8:0] _WTEMP_15;
    PAD_UNSIGNED #(.width(4), .n(9)) u_pad_65 (
        .y(_WTEMP_15),
        .in(4'hE)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_66 (
        .y(_node_26),
        .a(_WTEMP_15),
        .b(_arrivedPointer__q)
    );
    wire _node_27;
    BITWISEAND #(.width(1)) bitwiseand_67 (
        .y(_node_27),
        .a(1'h1),
        .b(_node_26)
    );
    wire [7:0] _GEN_24;
    MUX_UNSIGNED #(.width(8)) u_mux_68 (
        .y(_GEN_24),
        .sel(_node_27),
        .a(helloWorld_14),
        .b(_GEN_23)
    );
    wire _node_28;
    wire [8:0] _WTEMP_16;
    PAD_UNSIGNED #(.width(4), .n(9)) u_pad_69 (
        .y(_WTEMP_16),
        .in(4'hF)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_70 (
        .y(_node_28),
        .a(_WTEMP_16),
        .b(_arrivedPointer__q)
    );
    wire _node_29;
    BITWISEAND #(.width(1)) bitwiseand_71 (
        .y(_node_29),
        .a(1'h1),
        .b(_node_28)
    );
    wire [7:0] _GEN_25;
    MUX_UNSIGNED #(.width(8)) u_mux_72 (
        .y(_GEN_25),
        .sel(_node_29),
        .a(helloWorld_15),
        .b(_GEN_24)
    );
    wire _node_30;
    wire [8:0] _WTEMP_17;
    PAD_UNSIGNED #(.width(5), .n(9)) u_pad_73 (
        .y(_WTEMP_17),
        .in(5'h10)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_74 (
        .y(_node_30),
        .a(_WTEMP_17),
        .b(_arrivedPointer__q)
    );
    wire _node_31;
    BITWISEAND #(.width(1)) bitwiseand_75 (
        .y(_node_31),
        .a(1'h1),
        .b(_node_30)
    );
    wire [7:0] _GEN_26;
    MUX_UNSIGNED #(.width(8)) u_mux_76 (
        .y(_GEN_26),
        .sel(_node_31),
        .a(helloWorld_16),
        .b(_GEN_25)
    );
    wire _node_32;
    wire [8:0] _WTEMP_18;
    PAD_UNSIGNED #(.width(5), .n(9)) u_pad_77 (
        .y(_WTEMP_18),
        .in(5'h11)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_78 (
        .y(_node_32),
        .a(_WTEMP_18),
        .b(_arrivedPointer__q)
    );
    wire _node_33;
    BITWISEAND #(.width(1)) bitwiseand_79 (
        .y(_node_33),
        .a(1'h1),
        .b(_node_32)
    );
    wire [7:0] _GEN_27;
    MUX_UNSIGNED #(.width(8)) u_mux_80 (
        .y(_GEN_27),
        .sel(_node_33),
        .a(helloWorld_17),
        .b(_GEN_26)
    );
    wire _node_34;
    wire [8:0] _WTEMP_19;
    PAD_UNSIGNED #(.width(5), .n(9)) u_pad_81 (
        .y(_WTEMP_19),
        .in(5'h12)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_82 (
        .y(_node_34),
        .a(_WTEMP_19),
        .b(_arrivedPointer__q)
    );
    wire _node_35;
    BITWISEAND #(.width(1)) bitwiseand_83 (
        .y(_node_35),
        .a(1'h1),
        .b(_node_34)
    );
    wire [7:0] _GEN_28;
    MUX_UNSIGNED #(.width(8)) u_mux_84 (
        .y(_GEN_28),
        .sel(_node_35),
        .a(helloWorld_18),
        .b(_GEN_27)
    );
    wire _node_36;
    wire [8:0] _WTEMP_20;
    PAD_UNSIGNED #(.width(5), .n(9)) u_pad_85 (
        .y(_WTEMP_20),
        .in(5'h13)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_86 (
        .y(_node_36),
        .a(_WTEMP_20),
        .b(_arrivedPointer__q)
    );
    wire _node_37;
    BITWISEAND #(.width(1)) bitwiseand_87 (
        .y(_node_37),
        .a(1'h1),
        .b(_node_36)
    );
    wire [7:0] _GEN_29;
    MUX_UNSIGNED #(.width(8)) u_mux_88 (
        .y(_GEN_29),
        .sel(_node_37),
        .a(helloWorld_19),
        .b(_GEN_28)
    );
    wire _node_38;
    wire [8:0] _WTEMP_21;
    PAD_UNSIGNED #(.width(5), .n(9)) u_pad_89 (
        .y(_WTEMP_21),
        .in(5'h14)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_90 (
        .y(_node_38),
        .a(_WTEMP_21),
        .b(_arrivedPointer__q)
    );
    wire _node_39;
    BITWISEAND #(.width(1)) bitwiseand_91 (
        .y(_node_39),
        .a(1'h1),
        .b(_node_38)
    );
    wire [7:0] _GEN_30;
    MUX_UNSIGNED #(.width(8)) u_mux_92 (
        .y(_GEN_30),
        .sel(_node_39),
        .a(helloWorld_20),
        .b(_GEN_29)
    );
    wire _node_40;
    wire [8:0] _WTEMP_22;
    PAD_UNSIGNED #(.width(5), .n(9)) u_pad_93 (
        .y(_WTEMP_22),
        .in(5'h15)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_94 (
        .y(_node_40),
        .a(_WTEMP_22),
        .b(_arrivedPointer__q)
    );
    wire _node_41;
    BITWISEAND #(.width(1)) bitwiseand_95 (
        .y(_node_41),
        .a(1'h1),
        .b(_node_40)
    );
    wire [7:0] _GEN_31;
    MUX_UNSIGNED #(.width(8)) u_mux_96 (
        .y(_GEN_31),
        .sel(_node_41),
        .a(helloWorld_21),
        .b(_GEN_30)
    );
    wire _node_42;
    wire [8:0] _WTEMP_23;
    PAD_UNSIGNED #(.width(5), .n(9)) u_pad_97 (
        .y(_WTEMP_23),
        .in(5'h16)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_98 (
        .y(_node_42),
        .a(_WTEMP_23),
        .b(_arrivedPointer__q)
    );
    wire _node_43;
    BITWISEAND #(.width(1)) bitwiseand_99 (
        .y(_node_43),
        .a(1'h1),
        .b(_node_42)
    );
    wire [7:0] _GEN_32;
    MUX_UNSIGNED #(.width(8)) u_mux_100 (
        .y(_GEN_32),
        .sel(_node_43),
        .a(helloWorld_22),
        .b(_GEN_31)
    );
    wire _node_44;
    wire [8:0] _WTEMP_24;
    PAD_UNSIGNED #(.width(5), .n(9)) u_pad_101 (
        .y(_WTEMP_24),
        .in(5'h17)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_102 (
        .y(_node_44),
        .a(_WTEMP_24),
        .b(_arrivedPointer__q)
    );
    wire _node_45;
    BITWISEAND #(.width(1)) bitwiseand_103 (
        .y(_node_45),
        .a(1'h1),
        .b(_node_44)
    );
    wire [7:0] _GEN_33;
    MUX_UNSIGNED #(.width(8)) u_mux_104 (
        .y(_GEN_33),
        .sel(_node_45),
        .a(helloWorld_23),
        .b(_GEN_32)
    );
    wire _node_46;
    wire [8:0] _WTEMP_25;
    PAD_UNSIGNED #(.width(5), .n(9)) u_pad_105 (
        .y(_WTEMP_25),
        .in(5'h18)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_106 (
        .y(_node_46),
        .a(_WTEMP_25),
        .b(_arrivedPointer__q)
    );
    wire _node_47;
    BITWISEAND #(.width(1)) bitwiseand_107 (
        .y(_node_47),
        .a(1'h1),
        .b(_node_46)
    );
    wire [7:0] _GEN_34;
    MUX_UNSIGNED #(.width(8)) u_mux_108 (
        .y(_GEN_34),
        .sel(_node_47),
        .a(helloWorld_24),
        .b(_GEN_33)
    );
    wire _node_48;
    wire [8:0] _WTEMP_26;
    PAD_UNSIGNED #(.width(5), .n(9)) u_pad_109 (
        .y(_WTEMP_26),
        .in(5'h19)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_110 (
        .y(_node_48),
        .a(_WTEMP_26),
        .b(_arrivedPointer__q)
    );
    wire _node_49;
    BITWISEAND #(.width(1)) bitwiseand_111 (
        .y(_node_49),
        .a(1'h1),
        .b(_node_48)
    );
    wire [7:0] _GEN_35;
    MUX_UNSIGNED #(.width(8)) u_mux_112 (
        .y(_GEN_35),
        .sel(_node_49),
        .a(helloWorld_25),
        .b(_GEN_34)
    );
    wire _node_50;
    wire [8:0] _WTEMP_27;
    PAD_UNSIGNED #(.width(5), .n(9)) u_pad_113 (
        .y(_WTEMP_27),
        .in(5'h1A)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_114 (
        .y(_node_50),
        .a(_WTEMP_27),
        .b(_arrivedPointer__q)
    );
    wire _node_51;
    BITWISEAND #(.width(1)) bitwiseand_115 (
        .y(_node_51),
        .a(1'h1),
        .b(_node_50)
    );
    wire [7:0] _GEN_36;
    MUX_UNSIGNED #(.width(8)) u_mux_116 (
        .y(_GEN_36),
        .sel(_node_51),
        .a(helloWorld_26),
        .b(_GEN_35)
    );
    wire _node_52;
    wire [8:0] _WTEMP_28;
    PAD_UNSIGNED #(.width(5), .n(9)) u_pad_117 (
        .y(_WTEMP_28),
        .in(5'h1B)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_118 (
        .y(_node_52),
        .a(_WTEMP_28),
        .b(_arrivedPointer__q)
    );
    wire _node_53;
    BITWISEAND #(.width(1)) bitwiseand_119 (
        .y(_node_53),
        .a(1'h1),
        .b(_node_52)
    );
    wire [7:0] _GEN_37;
    MUX_UNSIGNED #(.width(8)) u_mux_120 (
        .y(_GEN_37),
        .sel(_node_53),
        .a(helloWorld_27),
        .b(_GEN_36)
    );
    wire _node_54;
    wire [8:0] _WTEMP_29;
    PAD_UNSIGNED #(.width(5), .n(9)) u_pad_121 (
        .y(_WTEMP_29),
        .in(5'h1C)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_122 (
        .y(_node_54),
        .a(_WTEMP_29),
        .b(_arrivedPointer__q)
    );
    wire _node_55;
    BITWISEAND #(.width(1)) bitwiseand_123 (
        .y(_node_55),
        .a(1'h1),
        .b(_node_54)
    );
    wire [7:0] _GEN_38;
    MUX_UNSIGNED #(.width(8)) u_mux_124 (
        .y(_GEN_38),
        .sel(_node_55),
        .a(helloWorld_28),
        .b(_GEN_37)
    );
    wire _node_56;
    wire [8:0] _WTEMP_30;
    PAD_UNSIGNED #(.width(5), .n(9)) u_pad_125 (
        .y(_WTEMP_30),
        .in(5'h1D)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_126 (
        .y(_node_56),
        .a(_WTEMP_30),
        .b(_arrivedPointer__q)
    );
    wire _node_57;
    BITWISEAND #(.width(1)) bitwiseand_127 (
        .y(_node_57),
        .a(1'h1),
        .b(_node_56)
    );
    wire [7:0] _GEN_39;
    MUX_UNSIGNED #(.width(8)) u_mux_128 (
        .y(_GEN_39),
        .sel(_node_57),
        .a(helloWorld_29),
        .b(_GEN_38)
    );
    wire _node_58;
    wire [8:0] _WTEMP_31;
    PAD_UNSIGNED #(.width(5), .n(9)) u_pad_129 (
        .y(_WTEMP_31),
        .in(5'h1E)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_130 (
        .y(_node_58),
        .a(_WTEMP_31),
        .b(_arrivedPointer__q)
    );
    wire _node_59;
    BITWISEAND #(.width(1)) bitwiseand_131 (
        .y(_node_59),
        .a(1'h1),
        .b(_node_58)
    );
    wire [7:0] _GEN_40;
    MUX_UNSIGNED #(.width(8)) u_mux_132 (
        .y(_GEN_40),
        .sel(_node_59),
        .a(helloWorld_30),
        .b(_GEN_39)
    );
    wire _node_60;
    wire [8:0] _WTEMP_32;
    PAD_UNSIGNED #(.width(5), .n(9)) u_pad_133 (
        .y(_WTEMP_32),
        .in(5'h1F)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_134 (
        .y(_node_60),
        .a(_WTEMP_32),
        .b(_arrivedPointer__q)
    );
    wire _node_61;
    BITWISEAND #(.width(1)) bitwiseand_135 (
        .y(_node_61),
        .a(1'h1),
        .b(_node_60)
    );
    wire [7:0] _GEN_41;
    MUX_UNSIGNED #(.width(8)) u_mux_136 (
        .y(_GEN_41),
        .sel(_node_61),
        .a(helloWorld_31),
        .b(_GEN_40)
    );
    wire _node_62;
    wire [8:0] _WTEMP_33;
    PAD_UNSIGNED #(.width(6), .n(9)) u_pad_137 (
        .y(_WTEMP_33),
        .in(6'h20)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_138 (
        .y(_node_62),
        .a(_WTEMP_33),
        .b(_arrivedPointer__q)
    );
    wire _node_63;
    BITWISEAND #(.width(1)) bitwiseand_139 (
        .y(_node_63),
        .a(1'h1),
        .b(_node_62)
    );
    wire [7:0] _GEN_42;
    MUX_UNSIGNED #(.width(8)) u_mux_140 (
        .y(_GEN_42),
        .sel(_node_63),
        .a(helloWorld_32),
        .b(_GEN_41)
    );
    wire _node_64;
    wire [8:0] _WTEMP_34;
    PAD_UNSIGNED #(.width(6), .n(9)) u_pad_141 (
        .y(_WTEMP_34),
        .in(6'h21)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_142 (
        .y(_node_64),
        .a(_WTEMP_34),
        .b(_arrivedPointer__q)
    );
    wire _node_65;
    BITWISEAND #(.width(1)) bitwiseand_143 (
        .y(_node_65),
        .a(1'h1),
        .b(_node_64)
    );
    wire [7:0] _GEN_43;
    MUX_UNSIGNED #(.width(8)) u_mux_144 (
        .y(_GEN_43),
        .sel(_node_65),
        .a(helloWorld_33),
        .b(_GEN_42)
    );
    wire _node_66;
    wire [8:0] _WTEMP_35;
    PAD_UNSIGNED #(.width(6), .n(9)) u_pad_145 (
        .y(_WTEMP_35),
        .in(6'h22)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_146 (
        .y(_node_66),
        .a(_WTEMP_35),
        .b(_arrivedPointer__q)
    );
    wire _node_67;
    BITWISEAND #(.width(1)) bitwiseand_147 (
        .y(_node_67),
        .a(1'h1),
        .b(_node_66)
    );
    wire [7:0] _GEN_44;
    MUX_UNSIGNED #(.width(8)) u_mux_148 (
        .y(_GEN_44),
        .sel(_node_67),
        .a(helloWorld_34),
        .b(_GEN_43)
    );
    wire _node_68;
    wire [8:0] _WTEMP_36;
    PAD_UNSIGNED #(.width(6), .n(9)) u_pad_149 (
        .y(_WTEMP_36),
        .in(6'h23)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_150 (
        .y(_node_68),
        .a(_WTEMP_36),
        .b(_arrivedPointer__q)
    );
    wire _node_69;
    BITWISEAND #(.width(1)) bitwiseand_151 (
        .y(_node_69),
        .a(1'h1),
        .b(_node_68)
    );
    wire [7:0] _GEN_45;
    MUX_UNSIGNED #(.width(8)) u_mux_152 (
        .y(_GEN_45),
        .sel(_node_69),
        .a(helloWorld_35),
        .b(_GEN_44)
    );
    wire _node_70;
    wire [8:0] _WTEMP_37;
    PAD_UNSIGNED #(.width(6), .n(9)) u_pad_153 (
        .y(_WTEMP_37),
        .in(6'h24)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_154 (
        .y(_node_70),
        .a(_WTEMP_37),
        .b(_arrivedPointer__q)
    );
    wire _node_71;
    BITWISEAND #(.width(1)) bitwiseand_155 (
        .y(_node_71),
        .a(1'h1),
        .b(_node_70)
    );
    wire [7:0] _GEN_46;
    MUX_UNSIGNED #(.width(8)) u_mux_156 (
        .y(_GEN_46),
        .sel(_node_71),
        .a(helloWorld_36),
        .b(_GEN_45)
    );
    wire _node_72;
    wire [8:0] _WTEMP_38;
    PAD_UNSIGNED #(.width(6), .n(9)) u_pad_157 (
        .y(_WTEMP_38),
        .in(6'h25)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_158 (
        .y(_node_72),
        .a(_WTEMP_38),
        .b(_arrivedPointer__q)
    );
    wire _node_73;
    BITWISEAND #(.width(1)) bitwiseand_159 (
        .y(_node_73),
        .a(1'h1),
        .b(_node_72)
    );
    wire [7:0] _GEN_47;
    MUX_UNSIGNED #(.width(8)) u_mux_160 (
        .y(_GEN_47),
        .sel(_node_73),
        .a(helloWorld_37),
        .b(_GEN_46)
    );
    wire _node_74;
    wire [8:0] _WTEMP_39;
    PAD_UNSIGNED #(.width(6), .n(9)) u_pad_161 (
        .y(_WTEMP_39),
        .in(6'h26)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_162 (
        .y(_node_74),
        .a(_WTEMP_39),
        .b(_arrivedPointer__q)
    );
    wire _node_75;
    BITWISEAND #(.width(1)) bitwiseand_163 (
        .y(_node_75),
        .a(1'h1),
        .b(_node_74)
    );
    wire [7:0] _GEN_48;
    MUX_UNSIGNED #(.width(8)) u_mux_164 (
        .y(_GEN_48),
        .sel(_node_75),
        .a(helloWorld_38),
        .b(_GEN_47)
    );
    wire _node_76;
    wire [8:0] _WTEMP_40;
    PAD_UNSIGNED #(.width(6), .n(9)) u_pad_165 (
        .y(_WTEMP_40),
        .in(6'h27)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_166 (
        .y(_node_76),
        .a(_WTEMP_40),
        .b(_arrivedPointer__q)
    );
    wire _node_77;
    BITWISEAND #(.width(1)) bitwiseand_167 (
        .y(_node_77),
        .a(1'h1),
        .b(_node_76)
    );
    wire [7:0] _GEN_49;
    MUX_UNSIGNED #(.width(8)) u_mux_168 (
        .y(_GEN_49),
        .sel(_node_77),
        .a(helloWorld_39),
        .b(_GEN_48)
    );
    wire _node_78;
    wire [8:0] _WTEMP_41;
    PAD_UNSIGNED #(.width(6), .n(9)) u_pad_169 (
        .y(_WTEMP_41),
        .in(6'h28)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_170 (
        .y(_node_78),
        .a(_WTEMP_41),
        .b(_arrivedPointer__q)
    );
    wire _node_79;
    BITWISEAND #(.width(1)) bitwiseand_171 (
        .y(_node_79),
        .a(1'h1),
        .b(_node_78)
    );
    wire [7:0] _GEN_50;
    MUX_UNSIGNED #(.width(8)) u_mux_172 (
        .y(_GEN_50),
        .sel(_node_79),
        .a(helloWorld_40),
        .b(_GEN_49)
    );
    wire _node_80;
    wire [8:0] _WTEMP_42;
    PAD_UNSIGNED #(.width(6), .n(9)) u_pad_173 (
        .y(_WTEMP_42),
        .in(6'h29)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_174 (
        .y(_node_80),
        .a(_WTEMP_42),
        .b(_arrivedPointer__q)
    );
    wire _node_81;
    BITWISEAND #(.width(1)) bitwiseand_175 (
        .y(_node_81),
        .a(1'h1),
        .b(_node_80)
    );
    wire [7:0] _GEN_51;
    MUX_UNSIGNED #(.width(8)) u_mux_176 (
        .y(_GEN_51),
        .sel(_node_81),
        .a(helloWorld_41),
        .b(_GEN_50)
    );
    wire _node_82;
    wire [8:0] _WTEMP_43;
    PAD_UNSIGNED #(.width(6), .n(9)) u_pad_177 (
        .y(_WTEMP_43),
        .in(6'h2A)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_178 (
        .y(_node_82),
        .a(_WTEMP_43),
        .b(_arrivedPointer__q)
    );
    wire _node_83;
    BITWISEAND #(.width(1)) bitwiseand_179 (
        .y(_node_83),
        .a(1'h1),
        .b(_node_82)
    );
    wire [7:0] _GEN_52;
    MUX_UNSIGNED #(.width(8)) u_mux_180 (
        .y(_GEN_52),
        .sel(_node_83),
        .a(helloWorld_42),
        .b(_GEN_51)
    );
    wire _node_84;
    wire [8:0] _WTEMP_44;
    PAD_UNSIGNED #(.width(6), .n(9)) u_pad_181 (
        .y(_WTEMP_44),
        .in(6'h2B)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_182 (
        .y(_node_84),
        .a(_WTEMP_44),
        .b(_arrivedPointer__q)
    );
    wire _node_85;
    BITWISEAND #(.width(1)) bitwiseand_183 (
        .y(_node_85),
        .a(1'h1),
        .b(_node_84)
    );
    wire [7:0] _GEN_53;
    MUX_UNSIGNED #(.width(8)) u_mux_184 (
        .y(_GEN_53),
        .sel(_node_85),
        .a(helloWorld_43),
        .b(_GEN_52)
    );
    wire _node_86;
    wire [8:0] _WTEMP_45;
    PAD_UNSIGNED #(.width(6), .n(9)) u_pad_185 (
        .y(_WTEMP_45),
        .in(6'h2C)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_186 (
        .y(_node_86),
        .a(_WTEMP_45),
        .b(_arrivedPointer__q)
    );
    wire _node_87;
    BITWISEAND #(.width(1)) bitwiseand_187 (
        .y(_node_87),
        .a(1'h1),
        .b(_node_86)
    );
    wire [7:0] _GEN_54;
    MUX_UNSIGNED #(.width(8)) u_mux_188 (
        .y(_GEN_54),
        .sel(_node_87),
        .a(helloWorld_44),
        .b(_GEN_53)
    );
    wire _node_88;
    wire [8:0] _WTEMP_46;
    PAD_UNSIGNED #(.width(6), .n(9)) u_pad_189 (
        .y(_WTEMP_46),
        .in(6'h2D)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_190 (
        .y(_node_88),
        .a(_WTEMP_46),
        .b(_arrivedPointer__q)
    );
    wire _node_89;
    BITWISEAND #(.width(1)) bitwiseand_191 (
        .y(_node_89),
        .a(1'h1),
        .b(_node_88)
    );
    wire [7:0] _GEN_55;
    MUX_UNSIGNED #(.width(8)) u_mux_192 (
        .y(_GEN_55),
        .sel(_node_89),
        .a(helloWorld_45),
        .b(_GEN_54)
    );
    wire _node_90;
    wire [8:0] _WTEMP_47;
    PAD_UNSIGNED #(.width(6), .n(9)) u_pad_193 (
        .y(_WTEMP_47),
        .in(6'h2E)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_194 (
        .y(_node_90),
        .a(_WTEMP_47),
        .b(_arrivedPointer__q)
    );
    wire _node_91;
    BITWISEAND #(.width(1)) bitwiseand_195 (
        .y(_node_91),
        .a(1'h1),
        .b(_node_90)
    );
    wire [7:0] _GEN_56;
    MUX_UNSIGNED #(.width(8)) u_mux_196 (
        .y(_GEN_56),
        .sel(_node_91),
        .a(helloWorld_46),
        .b(_GEN_55)
    );
    wire _node_92;
    wire [8:0] _WTEMP_48;
    PAD_UNSIGNED #(.width(6), .n(9)) u_pad_197 (
        .y(_WTEMP_48),
        .in(6'h2F)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_198 (
        .y(_node_92),
        .a(_WTEMP_48),
        .b(_arrivedPointer__q)
    );
    wire _node_93;
    BITWISEAND #(.width(1)) bitwiseand_199 (
        .y(_node_93),
        .a(1'h1),
        .b(_node_92)
    );
    wire [7:0] _GEN_57;
    MUX_UNSIGNED #(.width(8)) u_mux_200 (
        .y(_GEN_57),
        .sel(_node_93),
        .a(helloWorld_47),
        .b(_GEN_56)
    );
    wire _node_94;
    wire [8:0] _WTEMP_49;
    PAD_UNSIGNED #(.width(6), .n(9)) u_pad_201 (
        .y(_WTEMP_49),
        .in(6'h30)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_202 (
        .y(_node_94),
        .a(_WTEMP_49),
        .b(_arrivedPointer__q)
    );
    wire _node_95;
    BITWISEAND #(.width(1)) bitwiseand_203 (
        .y(_node_95),
        .a(1'h1),
        .b(_node_94)
    );
    wire [7:0] _GEN_58;
    MUX_UNSIGNED #(.width(8)) u_mux_204 (
        .y(_GEN_58),
        .sel(_node_95),
        .a(helloWorld_48),
        .b(_GEN_57)
    );
    wire _node_96;
    wire [8:0] _WTEMP_50;
    PAD_UNSIGNED #(.width(6), .n(9)) u_pad_205 (
        .y(_WTEMP_50),
        .in(6'h31)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_206 (
        .y(_node_96),
        .a(_WTEMP_50),
        .b(_arrivedPointer__q)
    );
    wire _node_97;
    BITWISEAND #(.width(1)) bitwiseand_207 (
        .y(_node_97),
        .a(1'h1),
        .b(_node_96)
    );
    wire [7:0] _GEN_59;
    MUX_UNSIGNED #(.width(8)) u_mux_208 (
        .y(_GEN_59),
        .sel(_node_97),
        .a(helloWorld_49),
        .b(_GEN_58)
    );
    wire _node_98;
    wire [8:0] _WTEMP_51;
    PAD_UNSIGNED #(.width(6), .n(9)) u_pad_209 (
        .y(_WTEMP_51),
        .in(6'h32)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_210 (
        .y(_node_98),
        .a(_WTEMP_51),
        .b(_arrivedPointer__q)
    );
    wire _node_99;
    BITWISEAND #(.width(1)) bitwiseand_211 (
        .y(_node_99),
        .a(1'h1),
        .b(_node_98)
    );
    wire [7:0] _GEN_60;
    MUX_UNSIGNED #(.width(8)) u_mux_212 (
        .y(_GEN_60),
        .sel(_node_99),
        .a(helloWorld_50),
        .b(_GEN_59)
    );
    wire _node_100;
    wire [8:0] _WTEMP_52;
    PAD_UNSIGNED #(.width(6), .n(9)) u_pad_213 (
        .y(_WTEMP_52),
        .in(6'h33)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_214 (
        .y(_node_100),
        .a(_WTEMP_52),
        .b(_arrivedPointer__q)
    );
    wire _node_101;
    BITWISEAND #(.width(1)) bitwiseand_215 (
        .y(_node_101),
        .a(1'h1),
        .b(_node_100)
    );
    wire [7:0] _GEN_61;
    MUX_UNSIGNED #(.width(8)) u_mux_216 (
        .y(_GEN_61),
        .sel(_node_101),
        .a(helloWorld_51),
        .b(_GEN_60)
    );
    wire _node_102;
    wire [8:0] _WTEMP_53;
    PAD_UNSIGNED #(.width(6), .n(9)) u_pad_217 (
        .y(_WTEMP_53),
        .in(6'h34)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_218 (
        .y(_node_102),
        .a(_WTEMP_53),
        .b(_arrivedPointer__q)
    );
    wire _node_103;
    BITWISEAND #(.width(1)) bitwiseand_219 (
        .y(_node_103),
        .a(1'h1),
        .b(_node_102)
    );
    wire [7:0] _GEN_62;
    MUX_UNSIGNED #(.width(8)) u_mux_220 (
        .y(_GEN_62),
        .sel(_node_103),
        .a(helloWorld_52),
        .b(_GEN_61)
    );
    wire _node_104;
    wire [8:0] _WTEMP_54;
    PAD_UNSIGNED #(.width(6), .n(9)) u_pad_221 (
        .y(_WTEMP_54),
        .in(6'h35)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_222 (
        .y(_node_104),
        .a(_WTEMP_54),
        .b(_arrivedPointer__q)
    );
    wire _node_105;
    BITWISEAND #(.width(1)) bitwiseand_223 (
        .y(_node_105),
        .a(1'h1),
        .b(_node_104)
    );
    wire [7:0] _GEN_63;
    MUX_UNSIGNED #(.width(8)) u_mux_224 (
        .y(_GEN_63),
        .sel(_node_105),
        .a(helloWorld_53),
        .b(_GEN_62)
    );
    wire _node_106;
    wire [8:0] _WTEMP_55;
    PAD_UNSIGNED #(.width(6), .n(9)) u_pad_225 (
        .y(_WTEMP_55),
        .in(6'h36)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_226 (
        .y(_node_106),
        .a(_WTEMP_55),
        .b(_arrivedPointer__q)
    );
    wire _node_107;
    BITWISEAND #(.width(1)) bitwiseand_227 (
        .y(_node_107),
        .a(1'h1),
        .b(_node_106)
    );
    wire [7:0] _GEN_64;
    MUX_UNSIGNED #(.width(8)) u_mux_228 (
        .y(_GEN_64),
        .sel(_node_107),
        .a(helloWorld_54),
        .b(_GEN_63)
    );
    wire _node_108;
    wire [8:0] _WTEMP_56;
    PAD_UNSIGNED #(.width(6), .n(9)) u_pad_229 (
        .y(_WTEMP_56),
        .in(6'h37)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_230 (
        .y(_node_108),
        .a(_WTEMP_56),
        .b(_arrivedPointer__q)
    );
    wire _node_109;
    BITWISEAND #(.width(1)) bitwiseand_231 (
        .y(_node_109),
        .a(1'h1),
        .b(_node_108)
    );
    wire [7:0] _GEN_65;
    MUX_UNSIGNED #(.width(8)) u_mux_232 (
        .y(_GEN_65),
        .sel(_node_109),
        .a(helloWorld_55),
        .b(_GEN_64)
    );
    wire _node_110;
    wire [8:0] _WTEMP_57;
    PAD_UNSIGNED #(.width(6), .n(9)) u_pad_233 (
        .y(_WTEMP_57),
        .in(6'h38)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_234 (
        .y(_node_110),
        .a(_WTEMP_57),
        .b(_arrivedPointer__q)
    );
    wire _node_111;
    BITWISEAND #(.width(1)) bitwiseand_235 (
        .y(_node_111),
        .a(1'h1),
        .b(_node_110)
    );
    wire [7:0] _GEN_66;
    MUX_UNSIGNED #(.width(8)) u_mux_236 (
        .y(_GEN_66),
        .sel(_node_111),
        .a(helloWorld_56),
        .b(_GEN_65)
    );
    wire _node_112;
    wire [8:0] _WTEMP_58;
    PAD_UNSIGNED #(.width(6), .n(9)) u_pad_237 (
        .y(_WTEMP_58),
        .in(6'h39)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_238 (
        .y(_node_112),
        .a(_WTEMP_58),
        .b(_arrivedPointer__q)
    );
    wire _node_113;
    BITWISEAND #(.width(1)) bitwiseand_239 (
        .y(_node_113),
        .a(1'h1),
        .b(_node_112)
    );
    wire [7:0] _GEN_67;
    MUX_UNSIGNED #(.width(8)) u_mux_240 (
        .y(_GEN_67),
        .sel(_node_113),
        .a(helloWorld_57),
        .b(_GEN_66)
    );
    wire _node_114;
    wire [8:0] _WTEMP_59;
    PAD_UNSIGNED #(.width(6), .n(9)) u_pad_241 (
        .y(_WTEMP_59),
        .in(6'h3A)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_242 (
        .y(_node_114),
        .a(_WTEMP_59),
        .b(_arrivedPointer__q)
    );
    wire _node_115;
    BITWISEAND #(.width(1)) bitwiseand_243 (
        .y(_node_115),
        .a(1'h1),
        .b(_node_114)
    );
    wire [7:0] _GEN_68;
    MUX_UNSIGNED #(.width(8)) u_mux_244 (
        .y(_GEN_68),
        .sel(_node_115),
        .a(helloWorld_58),
        .b(_GEN_67)
    );
    wire _node_116;
    wire [8:0] _WTEMP_60;
    PAD_UNSIGNED #(.width(6), .n(9)) u_pad_245 (
        .y(_WTEMP_60),
        .in(6'h3B)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_246 (
        .y(_node_116),
        .a(_WTEMP_60),
        .b(_arrivedPointer__q)
    );
    wire _node_117;
    BITWISEAND #(.width(1)) bitwiseand_247 (
        .y(_node_117),
        .a(1'h1),
        .b(_node_116)
    );
    wire [7:0] _GEN_69;
    MUX_UNSIGNED #(.width(8)) u_mux_248 (
        .y(_GEN_69),
        .sel(_node_117),
        .a(helloWorld_59),
        .b(_GEN_68)
    );
    wire _node_118;
    wire [8:0] _WTEMP_61;
    PAD_UNSIGNED #(.width(6), .n(9)) u_pad_249 (
        .y(_WTEMP_61),
        .in(6'h3C)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_250 (
        .y(_node_118),
        .a(_WTEMP_61),
        .b(_arrivedPointer__q)
    );
    wire _node_119;
    BITWISEAND #(.width(1)) bitwiseand_251 (
        .y(_node_119),
        .a(1'h1),
        .b(_node_118)
    );
    wire [7:0] _GEN_70;
    MUX_UNSIGNED #(.width(8)) u_mux_252 (
        .y(_GEN_70),
        .sel(_node_119),
        .a(helloWorld_60),
        .b(_GEN_69)
    );
    wire _node_120;
    wire [8:0] _WTEMP_62;
    PAD_UNSIGNED #(.width(6), .n(9)) u_pad_253 (
        .y(_WTEMP_62),
        .in(6'h3D)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_254 (
        .y(_node_120),
        .a(_WTEMP_62),
        .b(_arrivedPointer__q)
    );
    wire _node_121;
    BITWISEAND #(.width(1)) bitwiseand_255 (
        .y(_node_121),
        .a(1'h1),
        .b(_node_120)
    );
    wire [7:0] _GEN_71;
    MUX_UNSIGNED #(.width(8)) u_mux_256 (
        .y(_GEN_71),
        .sel(_node_121),
        .a(helloWorld_61),
        .b(_GEN_70)
    );
    wire _node_122;
    wire [8:0] _WTEMP_63;
    PAD_UNSIGNED #(.width(6), .n(9)) u_pad_257 (
        .y(_WTEMP_63),
        .in(6'h3E)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_258 (
        .y(_node_122),
        .a(_WTEMP_63),
        .b(_arrivedPointer__q)
    );
    wire _node_123;
    BITWISEAND #(.width(1)) bitwiseand_259 (
        .y(_node_123),
        .a(1'h1),
        .b(_node_122)
    );
    wire [7:0] _GEN_72;
    MUX_UNSIGNED #(.width(8)) u_mux_260 (
        .y(_GEN_72),
        .sel(_node_123),
        .a(helloWorld_62),
        .b(_GEN_71)
    );
    wire _node_124;
    wire [8:0] _WTEMP_64;
    PAD_UNSIGNED #(.width(6), .n(9)) u_pad_261 (
        .y(_WTEMP_64),
        .in(6'h3F)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_262 (
        .y(_node_124),
        .a(_WTEMP_64),
        .b(_arrivedPointer__q)
    );
    wire _node_125;
    BITWISEAND #(.width(1)) bitwiseand_263 (
        .y(_node_125),
        .a(1'h1),
        .b(_node_124)
    );
    wire [7:0] _GEN_73;
    MUX_UNSIGNED #(.width(8)) u_mux_264 (
        .y(_GEN_73),
        .sel(_node_125),
        .a(helloWorld_63),
        .b(_GEN_72)
    );
    wire _node_126;
    wire [8:0] _WTEMP_65;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_265 (
        .y(_WTEMP_65),
        .in(7'h40)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_266 (
        .y(_node_126),
        .a(_WTEMP_65),
        .b(_arrivedPointer__q)
    );
    wire _node_127;
    BITWISEAND #(.width(1)) bitwiseand_267 (
        .y(_node_127),
        .a(1'h1),
        .b(_node_126)
    );
    wire [7:0] _GEN_74;
    MUX_UNSIGNED #(.width(8)) u_mux_268 (
        .y(_GEN_74),
        .sel(_node_127),
        .a(helloWorld_64),
        .b(_GEN_73)
    );
    wire _node_128;
    wire [8:0] _WTEMP_66;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_269 (
        .y(_WTEMP_66),
        .in(7'h41)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_270 (
        .y(_node_128),
        .a(_WTEMP_66),
        .b(_arrivedPointer__q)
    );
    wire _node_129;
    BITWISEAND #(.width(1)) bitwiseand_271 (
        .y(_node_129),
        .a(1'h1),
        .b(_node_128)
    );
    wire [7:0] _GEN_75;
    MUX_UNSIGNED #(.width(8)) u_mux_272 (
        .y(_GEN_75),
        .sel(_node_129),
        .a(helloWorld_65),
        .b(_GEN_74)
    );
    wire _node_130;
    wire [8:0] _WTEMP_67;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_273 (
        .y(_WTEMP_67),
        .in(7'h42)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_274 (
        .y(_node_130),
        .a(_WTEMP_67),
        .b(_arrivedPointer__q)
    );
    wire _node_131;
    BITWISEAND #(.width(1)) bitwiseand_275 (
        .y(_node_131),
        .a(1'h1),
        .b(_node_130)
    );
    wire [7:0] _GEN_76;
    MUX_UNSIGNED #(.width(8)) u_mux_276 (
        .y(_GEN_76),
        .sel(_node_131),
        .a(helloWorld_66),
        .b(_GEN_75)
    );
    wire _node_132;
    wire [8:0] _WTEMP_68;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_277 (
        .y(_WTEMP_68),
        .in(7'h43)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_278 (
        .y(_node_132),
        .a(_WTEMP_68),
        .b(_arrivedPointer__q)
    );
    wire _node_133;
    BITWISEAND #(.width(1)) bitwiseand_279 (
        .y(_node_133),
        .a(1'h1),
        .b(_node_132)
    );
    wire [7:0] _GEN_77;
    MUX_UNSIGNED #(.width(8)) u_mux_280 (
        .y(_GEN_77),
        .sel(_node_133),
        .a(helloWorld_67),
        .b(_GEN_76)
    );
    wire _node_134;
    wire [8:0] _WTEMP_69;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_281 (
        .y(_WTEMP_69),
        .in(7'h44)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_282 (
        .y(_node_134),
        .a(_WTEMP_69),
        .b(_arrivedPointer__q)
    );
    wire _node_135;
    BITWISEAND #(.width(1)) bitwiseand_283 (
        .y(_node_135),
        .a(1'h1),
        .b(_node_134)
    );
    wire [7:0] _GEN_78;
    MUX_UNSIGNED #(.width(8)) u_mux_284 (
        .y(_GEN_78),
        .sel(_node_135),
        .a(helloWorld_68),
        .b(_GEN_77)
    );
    wire _node_136;
    wire [8:0] _WTEMP_70;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_285 (
        .y(_WTEMP_70),
        .in(7'h45)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_286 (
        .y(_node_136),
        .a(_WTEMP_70),
        .b(_arrivedPointer__q)
    );
    wire _node_137;
    BITWISEAND #(.width(1)) bitwiseand_287 (
        .y(_node_137),
        .a(1'h1),
        .b(_node_136)
    );
    wire [7:0] _GEN_79;
    MUX_UNSIGNED #(.width(8)) u_mux_288 (
        .y(_GEN_79),
        .sel(_node_137),
        .a(helloWorld_69),
        .b(_GEN_78)
    );
    wire _node_138;
    wire [8:0] _WTEMP_71;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_289 (
        .y(_WTEMP_71),
        .in(7'h46)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_290 (
        .y(_node_138),
        .a(_WTEMP_71),
        .b(_arrivedPointer__q)
    );
    wire _node_139;
    BITWISEAND #(.width(1)) bitwiseand_291 (
        .y(_node_139),
        .a(1'h1),
        .b(_node_138)
    );
    wire [7:0] _GEN_80;
    MUX_UNSIGNED #(.width(8)) u_mux_292 (
        .y(_GEN_80),
        .sel(_node_139),
        .a(helloWorld_70),
        .b(_GEN_79)
    );
    wire _node_140;
    wire [8:0] _WTEMP_72;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_293 (
        .y(_WTEMP_72),
        .in(7'h47)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_294 (
        .y(_node_140),
        .a(_WTEMP_72),
        .b(_arrivedPointer__q)
    );
    wire _node_141;
    BITWISEAND #(.width(1)) bitwiseand_295 (
        .y(_node_141),
        .a(1'h1),
        .b(_node_140)
    );
    wire [7:0] _GEN_81;
    MUX_UNSIGNED #(.width(8)) u_mux_296 (
        .y(_GEN_81),
        .sel(_node_141),
        .a(helloWorld_71),
        .b(_GEN_80)
    );
    wire _node_142;
    wire [8:0] _WTEMP_73;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_297 (
        .y(_WTEMP_73),
        .in(7'h48)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_298 (
        .y(_node_142),
        .a(_WTEMP_73),
        .b(_arrivedPointer__q)
    );
    wire _node_143;
    BITWISEAND #(.width(1)) bitwiseand_299 (
        .y(_node_143),
        .a(1'h1),
        .b(_node_142)
    );
    wire [7:0] _GEN_82;
    MUX_UNSIGNED #(.width(8)) u_mux_300 (
        .y(_GEN_82),
        .sel(_node_143),
        .a(helloWorld_72),
        .b(_GEN_81)
    );
    wire _node_144;
    wire [8:0] _WTEMP_74;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_301 (
        .y(_WTEMP_74),
        .in(7'h49)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_302 (
        .y(_node_144),
        .a(_WTEMP_74),
        .b(_arrivedPointer__q)
    );
    wire _node_145;
    BITWISEAND #(.width(1)) bitwiseand_303 (
        .y(_node_145),
        .a(1'h1),
        .b(_node_144)
    );
    wire [7:0] _GEN_83;
    MUX_UNSIGNED #(.width(8)) u_mux_304 (
        .y(_GEN_83),
        .sel(_node_145),
        .a(helloWorld_73),
        .b(_GEN_82)
    );
    wire _node_146;
    wire [8:0] _WTEMP_75;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_305 (
        .y(_WTEMP_75),
        .in(7'h4A)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_306 (
        .y(_node_146),
        .a(_WTEMP_75),
        .b(_arrivedPointer__q)
    );
    wire _node_147;
    BITWISEAND #(.width(1)) bitwiseand_307 (
        .y(_node_147),
        .a(1'h1),
        .b(_node_146)
    );
    wire [7:0] _GEN_84;
    MUX_UNSIGNED #(.width(8)) u_mux_308 (
        .y(_GEN_84),
        .sel(_node_147),
        .a(helloWorld_74),
        .b(_GEN_83)
    );
    wire _node_148;
    wire [8:0] _WTEMP_76;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_309 (
        .y(_WTEMP_76),
        .in(7'h4B)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_310 (
        .y(_node_148),
        .a(_WTEMP_76),
        .b(_arrivedPointer__q)
    );
    wire _node_149;
    BITWISEAND #(.width(1)) bitwiseand_311 (
        .y(_node_149),
        .a(1'h1),
        .b(_node_148)
    );
    wire [7:0] _GEN_85;
    MUX_UNSIGNED #(.width(8)) u_mux_312 (
        .y(_GEN_85),
        .sel(_node_149),
        .a(helloWorld_75),
        .b(_GEN_84)
    );
    wire _node_150;
    wire [8:0] _WTEMP_77;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_313 (
        .y(_WTEMP_77),
        .in(7'h4C)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_314 (
        .y(_node_150),
        .a(_WTEMP_77),
        .b(_arrivedPointer__q)
    );
    wire _node_151;
    BITWISEAND #(.width(1)) bitwiseand_315 (
        .y(_node_151),
        .a(1'h1),
        .b(_node_150)
    );
    wire [7:0] _GEN_86;
    MUX_UNSIGNED #(.width(8)) u_mux_316 (
        .y(_GEN_86),
        .sel(_node_151),
        .a(helloWorld_76),
        .b(_GEN_85)
    );
    wire _node_152;
    wire [8:0] _WTEMP_78;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_317 (
        .y(_WTEMP_78),
        .in(7'h4D)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_318 (
        .y(_node_152),
        .a(_WTEMP_78),
        .b(_arrivedPointer__q)
    );
    wire _node_153;
    BITWISEAND #(.width(1)) bitwiseand_319 (
        .y(_node_153),
        .a(1'h1),
        .b(_node_152)
    );
    wire [7:0] _GEN_87;
    MUX_UNSIGNED #(.width(8)) u_mux_320 (
        .y(_GEN_87),
        .sel(_node_153),
        .a(helloWorld_77),
        .b(_GEN_86)
    );
    wire _node_154;
    wire [8:0] _WTEMP_79;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_321 (
        .y(_WTEMP_79),
        .in(7'h4E)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_322 (
        .y(_node_154),
        .a(_WTEMP_79),
        .b(_arrivedPointer__q)
    );
    wire _node_155;
    BITWISEAND #(.width(1)) bitwiseand_323 (
        .y(_node_155),
        .a(1'h1),
        .b(_node_154)
    );
    wire [7:0] _GEN_88;
    MUX_UNSIGNED #(.width(8)) u_mux_324 (
        .y(_GEN_88),
        .sel(_node_155),
        .a(helloWorld_78),
        .b(_GEN_87)
    );
    wire _node_156;
    wire [8:0] _WTEMP_80;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_325 (
        .y(_WTEMP_80),
        .in(7'h4F)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_326 (
        .y(_node_156),
        .a(_WTEMP_80),
        .b(_arrivedPointer__q)
    );
    wire _node_157;
    BITWISEAND #(.width(1)) bitwiseand_327 (
        .y(_node_157),
        .a(1'h1),
        .b(_node_156)
    );
    wire [7:0] _GEN_89;
    MUX_UNSIGNED #(.width(8)) u_mux_328 (
        .y(_GEN_89),
        .sel(_node_157),
        .a(helloWorld_79),
        .b(_GEN_88)
    );
    wire _node_158;
    wire [8:0] _WTEMP_81;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_329 (
        .y(_WTEMP_81),
        .in(7'h50)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_330 (
        .y(_node_158),
        .a(_WTEMP_81),
        .b(_arrivedPointer__q)
    );
    wire _node_159;
    BITWISEAND #(.width(1)) bitwiseand_331 (
        .y(_node_159),
        .a(1'h1),
        .b(_node_158)
    );
    wire [7:0] _GEN_90;
    MUX_UNSIGNED #(.width(8)) u_mux_332 (
        .y(_GEN_90),
        .sel(_node_159),
        .a(helloWorld_80),
        .b(_GEN_89)
    );
    wire _node_160;
    wire [8:0] _WTEMP_82;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_333 (
        .y(_WTEMP_82),
        .in(7'h51)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_334 (
        .y(_node_160),
        .a(_WTEMP_82),
        .b(_arrivedPointer__q)
    );
    wire _node_161;
    BITWISEAND #(.width(1)) bitwiseand_335 (
        .y(_node_161),
        .a(1'h1),
        .b(_node_160)
    );
    wire [7:0] _GEN_91;
    MUX_UNSIGNED #(.width(8)) u_mux_336 (
        .y(_GEN_91),
        .sel(_node_161),
        .a(helloWorld_81),
        .b(_GEN_90)
    );
    wire _node_162;
    wire [8:0] _WTEMP_83;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_337 (
        .y(_WTEMP_83),
        .in(7'h52)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_338 (
        .y(_node_162),
        .a(_WTEMP_83),
        .b(_arrivedPointer__q)
    );
    wire _node_163;
    BITWISEAND #(.width(1)) bitwiseand_339 (
        .y(_node_163),
        .a(1'h1),
        .b(_node_162)
    );
    wire [7:0] _GEN_92;
    MUX_UNSIGNED #(.width(8)) u_mux_340 (
        .y(_GEN_92),
        .sel(_node_163),
        .a(helloWorld_82),
        .b(_GEN_91)
    );
    wire _node_164;
    wire [8:0] _WTEMP_84;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_341 (
        .y(_WTEMP_84),
        .in(7'h53)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_342 (
        .y(_node_164),
        .a(_WTEMP_84),
        .b(_arrivedPointer__q)
    );
    wire _node_165;
    BITWISEAND #(.width(1)) bitwiseand_343 (
        .y(_node_165),
        .a(1'h1),
        .b(_node_164)
    );
    wire [7:0] _GEN_93;
    MUX_UNSIGNED #(.width(8)) u_mux_344 (
        .y(_GEN_93),
        .sel(_node_165),
        .a(helloWorld_83),
        .b(_GEN_92)
    );
    wire _node_166;
    wire [8:0] _WTEMP_85;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_345 (
        .y(_WTEMP_85),
        .in(7'h54)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_346 (
        .y(_node_166),
        .a(_WTEMP_85),
        .b(_arrivedPointer__q)
    );
    wire _node_167;
    BITWISEAND #(.width(1)) bitwiseand_347 (
        .y(_node_167),
        .a(1'h1),
        .b(_node_166)
    );
    wire [7:0] _GEN_94;
    MUX_UNSIGNED #(.width(8)) u_mux_348 (
        .y(_GEN_94),
        .sel(_node_167),
        .a(helloWorld_84),
        .b(_GEN_93)
    );
    wire _node_168;
    wire [8:0] _WTEMP_86;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_349 (
        .y(_WTEMP_86),
        .in(7'h55)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_350 (
        .y(_node_168),
        .a(_WTEMP_86),
        .b(_arrivedPointer__q)
    );
    wire _node_169;
    BITWISEAND #(.width(1)) bitwiseand_351 (
        .y(_node_169),
        .a(1'h1),
        .b(_node_168)
    );
    wire [7:0] _GEN_95;
    MUX_UNSIGNED #(.width(8)) u_mux_352 (
        .y(_GEN_95),
        .sel(_node_169),
        .a(helloWorld_85),
        .b(_GEN_94)
    );
    wire _node_170;
    wire [8:0] _WTEMP_87;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_353 (
        .y(_WTEMP_87),
        .in(7'h56)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_354 (
        .y(_node_170),
        .a(_WTEMP_87),
        .b(_arrivedPointer__q)
    );
    wire _node_171;
    BITWISEAND #(.width(1)) bitwiseand_355 (
        .y(_node_171),
        .a(1'h1),
        .b(_node_170)
    );
    wire [7:0] _GEN_96;
    MUX_UNSIGNED #(.width(8)) u_mux_356 (
        .y(_GEN_96),
        .sel(_node_171),
        .a(helloWorld_86),
        .b(_GEN_95)
    );
    wire _node_172;
    wire [8:0] _WTEMP_88;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_357 (
        .y(_WTEMP_88),
        .in(7'h57)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_358 (
        .y(_node_172),
        .a(_WTEMP_88),
        .b(_arrivedPointer__q)
    );
    wire _node_173;
    BITWISEAND #(.width(1)) bitwiseand_359 (
        .y(_node_173),
        .a(1'h1),
        .b(_node_172)
    );
    wire [7:0] _GEN_97;
    MUX_UNSIGNED #(.width(8)) u_mux_360 (
        .y(_GEN_97),
        .sel(_node_173),
        .a(helloWorld_87),
        .b(_GEN_96)
    );
    wire _node_174;
    wire [8:0] _WTEMP_89;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_361 (
        .y(_WTEMP_89),
        .in(7'h58)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_362 (
        .y(_node_174),
        .a(_WTEMP_89),
        .b(_arrivedPointer__q)
    );
    wire _node_175;
    BITWISEAND #(.width(1)) bitwiseand_363 (
        .y(_node_175),
        .a(1'h1),
        .b(_node_174)
    );
    wire [7:0] _GEN_98;
    MUX_UNSIGNED #(.width(8)) u_mux_364 (
        .y(_GEN_98),
        .sel(_node_175),
        .a(helloWorld_88),
        .b(_GEN_97)
    );
    wire _node_176;
    wire [8:0] _WTEMP_90;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_365 (
        .y(_WTEMP_90),
        .in(7'h59)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_366 (
        .y(_node_176),
        .a(_WTEMP_90),
        .b(_arrivedPointer__q)
    );
    wire _node_177;
    BITWISEAND #(.width(1)) bitwiseand_367 (
        .y(_node_177),
        .a(1'h1),
        .b(_node_176)
    );
    wire [7:0] _GEN_99;
    MUX_UNSIGNED #(.width(8)) u_mux_368 (
        .y(_GEN_99),
        .sel(_node_177),
        .a(helloWorld_89),
        .b(_GEN_98)
    );
    wire _node_178;
    wire [8:0] _WTEMP_91;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_369 (
        .y(_WTEMP_91),
        .in(7'h5A)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_370 (
        .y(_node_178),
        .a(_WTEMP_91),
        .b(_arrivedPointer__q)
    );
    wire _node_179;
    BITWISEAND #(.width(1)) bitwiseand_371 (
        .y(_node_179),
        .a(1'h1),
        .b(_node_178)
    );
    wire [7:0] _GEN_100;
    MUX_UNSIGNED #(.width(8)) u_mux_372 (
        .y(_GEN_100),
        .sel(_node_179),
        .a(helloWorld_90),
        .b(_GEN_99)
    );
    wire _node_180;
    wire [8:0] _WTEMP_92;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_373 (
        .y(_WTEMP_92),
        .in(7'h5B)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_374 (
        .y(_node_180),
        .a(_WTEMP_92),
        .b(_arrivedPointer__q)
    );
    wire _node_181;
    BITWISEAND #(.width(1)) bitwiseand_375 (
        .y(_node_181),
        .a(1'h1),
        .b(_node_180)
    );
    wire [7:0] _GEN_101;
    MUX_UNSIGNED #(.width(8)) u_mux_376 (
        .y(_GEN_101),
        .sel(_node_181),
        .a(helloWorld_91),
        .b(_GEN_100)
    );
    wire _node_182;
    wire [8:0] _WTEMP_93;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_377 (
        .y(_WTEMP_93),
        .in(7'h5C)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_378 (
        .y(_node_182),
        .a(_WTEMP_93),
        .b(_arrivedPointer__q)
    );
    wire _node_183;
    BITWISEAND #(.width(1)) bitwiseand_379 (
        .y(_node_183),
        .a(1'h1),
        .b(_node_182)
    );
    wire [7:0] _GEN_102;
    MUX_UNSIGNED #(.width(8)) u_mux_380 (
        .y(_GEN_102),
        .sel(_node_183),
        .a(helloWorld_92),
        .b(_GEN_101)
    );
    wire _node_184;
    wire [8:0] _WTEMP_94;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_381 (
        .y(_WTEMP_94),
        .in(7'h5D)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_382 (
        .y(_node_184),
        .a(_WTEMP_94),
        .b(_arrivedPointer__q)
    );
    wire _node_185;
    BITWISEAND #(.width(1)) bitwiseand_383 (
        .y(_node_185),
        .a(1'h1),
        .b(_node_184)
    );
    wire [7:0] _GEN_103;
    MUX_UNSIGNED #(.width(8)) u_mux_384 (
        .y(_GEN_103),
        .sel(_node_185),
        .a(helloWorld_93),
        .b(_GEN_102)
    );
    wire _node_186;
    wire [8:0] _WTEMP_95;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_385 (
        .y(_WTEMP_95),
        .in(7'h5E)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_386 (
        .y(_node_186),
        .a(_WTEMP_95),
        .b(_arrivedPointer__q)
    );
    wire _node_187;
    BITWISEAND #(.width(1)) bitwiseand_387 (
        .y(_node_187),
        .a(1'h1),
        .b(_node_186)
    );
    wire [7:0] _GEN_104;
    MUX_UNSIGNED #(.width(8)) u_mux_388 (
        .y(_GEN_104),
        .sel(_node_187),
        .a(helloWorld_94),
        .b(_GEN_103)
    );
    wire _node_188;
    wire [8:0] _WTEMP_96;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_389 (
        .y(_WTEMP_96),
        .in(7'h5F)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_390 (
        .y(_node_188),
        .a(_WTEMP_96),
        .b(_arrivedPointer__q)
    );
    wire _node_189;
    BITWISEAND #(.width(1)) bitwiseand_391 (
        .y(_node_189),
        .a(1'h1),
        .b(_node_188)
    );
    wire [7:0] _GEN_105;
    MUX_UNSIGNED #(.width(8)) u_mux_392 (
        .y(_GEN_105),
        .sel(_node_189),
        .a(helloWorld_95),
        .b(_GEN_104)
    );
    wire _node_190;
    wire [8:0] _WTEMP_97;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_393 (
        .y(_WTEMP_97),
        .in(7'h60)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_394 (
        .y(_node_190),
        .a(_WTEMP_97),
        .b(_arrivedPointer__q)
    );
    wire _node_191;
    BITWISEAND #(.width(1)) bitwiseand_395 (
        .y(_node_191),
        .a(1'h1),
        .b(_node_190)
    );
    wire [7:0] _GEN_106;
    MUX_UNSIGNED #(.width(8)) u_mux_396 (
        .y(_GEN_106),
        .sel(_node_191),
        .a(helloWorld_96),
        .b(_GEN_105)
    );
    wire _node_192;
    wire [8:0] _WTEMP_98;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_397 (
        .y(_WTEMP_98),
        .in(7'h61)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_398 (
        .y(_node_192),
        .a(_WTEMP_98),
        .b(_arrivedPointer__q)
    );
    wire _node_193;
    BITWISEAND #(.width(1)) bitwiseand_399 (
        .y(_node_193),
        .a(1'h1),
        .b(_node_192)
    );
    wire [7:0] _GEN_107;
    MUX_UNSIGNED #(.width(8)) u_mux_400 (
        .y(_GEN_107),
        .sel(_node_193),
        .a(helloWorld_97),
        .b(_GEN_106)
    );
    wire _node_194;
    wire [8:0] _WTEMP_99;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_401 (
        .y(_WTEMP_99),
        .in(7'h62)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_402 (
        .y(_node_194),
        .a(_WTEMP_99),
        .b(_arrivedPointer__q)
    );
    wire _node_195;
    BITWISEAND #(.width(1)) bitwiseand_403 (
        .y(_node_195),
        .a(1'h1),
        .b(_node_194)
    );
    wire [7:0] _GEN_108;
    MUX_UNSIGNED #(.width(8)) u_mux_404 (
        .y(_GEN_108),
        .sel(_node_195),
        .a(helloWorld_98),
        .b(_GEN_107)
    );
    wire _node_196;
    wire [8:0] _WTEMP_100;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_405 (
        .y(_WTEMP_100),
        .in(7'h63)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_406 (
        .y(_node_196),
        .a(_WTEMP_100),
        .b(_arrivedPointer__q)
    );
    wire _node_197;
    BITWISEAND #(.width(1)) bitwiseand_407 (
        .y(_node_197),
        .a(1'h1),
        .b(_node_196)
    );
    wire [7:0] _GEN_109;
    MUX_UNSIGNED #(.width(8)) u_mux_408 (
        .y(_GEN_109),
        .sel(_node_197),
        .a(helloWorld_99),
        .b(_GEN_108)
    );
    wire _node_198;
    wire [8:0] _WTEMP_101;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_409 (
        .y(_WTEMP_101),
        .in(7'h64)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_410 (
        .y(_node_198),
        .a(_WTEMP_101),
        .b(_arrivedPointer__q)
    );
    wire _node_199;
    BITWISEAND #(.width(1)) bitwiseand_411 (
        .y(_node_199),
        .a(1'h1),
        .b(_node_198)
    );
    wire [7:0] _GEN_110;
    MUX_UNSIGNED #(.width(8)) u_mux_412 (
        .y(_GEN_110),
        .sel(_node_199),
        .a(helloWorld_100),
        .b(_GEN_109)
    );
    wire _node_200;
    wire [8:0] _WTEMP_102;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_413 (
        .y(_WTEMP_102),
        .in(7'h65)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_414 (
        .y(_node_200),
        .a(_WTEMP_102),
        .b(_arrivedPointer__q)
    );
    wire _node_201;
    BITWISEAND #(.width(1)) bitwiseand_415 (
        .y(_node_201),
        .a(1'h1),
        .b(_node_200)
    );
    wire [7:0] _GEN_111;
    MUX_UNSIGNED #(.width(8)) u_mux_416 (
        .y(_GEN_111),
        .sel(_node_201),
        .a(helloWorld_101),
        .b(_GEN_110)
    );
    wire _node_202;
    wire [8:0] _WTEMP_103;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_417 (
        .y(_WTEMP_103),
        .in(7'h66)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_418 (
        .y(_node_202),
        .a(_WTEMP_103),
        .b(_arrivedPointer__q)
    );
    wire _node_203;
    BITWISEAND #(.width(1)) bitwiseand_419 (
        .y(_node_203),
        .a(1'h1),
        .b(_node_202)
    );
    wire [7:0] _GEN_112;
    MUX_UNSIGNED #(.width(8)) u_mux_420 (
        .y(_GEN_112),
        .sel(_node_203),
        .a(helloWorld_102),
        .b(_GEN_111)
    );
    wire _node_204;
    wire [8:0] _WTEMP_104;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_421 (
        .y(_WTEMP_104),
        .in(7'h67)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_422 (
        .y(_node_204),
        .a(_WTEMP_104),
        .b(_arrivedPointer__q)
    );
    wire _node_205;
    BITWISEAND #(.width(1)) bitwiseand_423 (
        .y(_node_205),
        .a(1'h1),
        .b(_node_204)
    );
    wire [7:0] _GEN_113;
    MUX_UNSIGNED #(.width(8)) u_mux_424 (
        .y(_GEN_113),
        .sel(_node_205),
        .a(helloWorld_103),
        .b(_GEN_112)
    );
    wire _node_206;
    wire [8:0] _WTEMP_105;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_425 (
        .y(_WTEMP_105),
        .in(7'h68)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_426 (
        .y(_node_206),
        .a(_WTEMP_105),
        .b(_arrivedPointer__q)
    );
    wire _node_207;
    BITWISEAND #(.width(1)) bitwiseand_427 (
        .y(_node_207),
        .a(1'h1),
        .b(_node_206)
    );
    wire [7:0] _GEN_114;
    MUX_UNSIGNED #(.width(8)) u_mux_428 (
        .y(_GEN_114),
        .sel(_node_207),
        .a(helloWorld_104),
        .b(_GEN_113)
    );
    wire _node_208;
    wire [8:0] _WTEMP_106;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_429 (
        .y(_WTEMP_106),
        .in(7'h69)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_430 (
        .y(_node_208),
        .a(_WTEMP_106),
        .b(_arrivedPointer__q)
    );
    wire _node_209;
    BITWISEAND #(.width(1)) bitwiseand_431 (
        .y(_node_209),
        .a(1'h1),
        .b(_node_208)
    );
    wire [7:0] _GEN_115;
    MUX_UNSIGNED #(.width(8)) u_mux_432 (
        .y(_GEN_115),
        .sel(_node_209),
        .a(helloWorld_105),
        .b(_GEN_114)
    );
    wire _node_210;
    wire [8:0] _WTEMP_107;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_433 (
        .y(_WTEMP_107),
        .in(7'h6A)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_434 (
        .y(_node_210),
        .a(_WTEMP_107),
        .b(_arrivedPointer__q)
    );
    wire _node_211;
    BITWISEAND #(.width(1)) bitwiseand_435 (
        .y(_node_211),
        .a(1'h1),
        .b(_node_210)
    );
    wire [7:0] _GEN_116;
    MUX_UNSIGNED #(.width(8)) u_mux_436 (
        .y(_GEN_116),
        .sel(_node_211),
        .a(helloWorld_106),
        .b(_GEN_115)
    );
    wire _node_212;
    wire [8:0] _WTEMP_108;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_437 (
        .y(_WTEMP_108),
        .in(7'h6B)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_438 (
        .y(_node_212),
        .a(_WTEMP_108),
        .b(_arrivedPointer__q)
    );
    wire _node_213;
    BITWISEAND #(.width(1)) bitwiseand_439 (
        .y(_node_213),
        .a(1'h1),
        .b(_node_212)
    );
    wire [7:0] _GEN_117;
    MUX_UNSIGNED #(.width(8)) u_mux_440 (
        .y(_GEN_117),
        .sel(_node_213),
        .a(helloWorld_107),
        .b(_GEN_116)
    );
    wire _node_214;
    wire [8:0] _WTEMP_109;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_441 (
        .y(_WTEMP_109),
        .in(7'h6C)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_442 (
        .y(_node_214),
        .a(_WTEMP_109),
        .b(_arrivedPointer__q)
    );
    wire _node_215;
    BITWISEAND #(.width(1)) bitwiseand_443 (
        .y(_node_215),
        .a(1'h1),
        .b(_node_214)
    );
    wire [7:0] _GEN_118;
    MUX_UNSIGNED #(.width(8)) u_mux_444 (
        .y(_GEN_118),
        .sel(_node_215),
        .a(helloWorld_108),
        .b(_GEN_117)
    );
    wire _node_216;
    wire [8:0] _WTEMP_110;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_445 (
        .y(_WTEMP_110),
        .in(7'h6D)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_446 (
        .y(_node_216),
        .a(_WTEMP_110),
        .b(_arrivedPointer__q)
    );
    wire _node_217;
    BITWISEAND #(.width(1)) bitwiseand_447 (
        .y(_node_217),
        .a(1'h1),
        .b(_node_216)
    );
    wire [7:0] _GEN_119;
    MUX_UNSIGNED #(.width(8)) u_mux_448 (
        .y(_GEN_119),
        .sel(_node_217),
        .a(helloWorld_109),
        .b(_GEN_118)
    );
    wire _node_218;
    wire [8:0] _WTEMP_111;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_449 (
        .y(_WTEMP_111),
        .in(7'h6E)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_450 (
        .y(_node_218),
        .a(_WTEMP_111),
        .b(_arrivedPointer__q)
    );
    wire _node_219;
    BITWISEAND #(.width(1)) bitwiseand_451 (
        .y(_node_219),
        .a(1'h1),
        .b(_node_218)
    );
    wire [7:0] _GEN_120;
    MUX_UNSIGNED #(.width(8)) u_mux_452 (
        .y(_GEN_120),
        .sel(_node_219),
        .a(helloWorld_110),
        .b(_GEN_119)
    );
    wire _node_220;
    wire [8:0] _WTEMP_112;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_453 (
        .y(_WTEMP_112),
        .in(7'h6F)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_454 (
        .y(_node_220),
        .a(_WTEMP_112),
        .b(_arrivedPointer__q)
    );
    wire _node_221;
    BITWISEAND #(.width(1)) bitwiseand_455 (
        .y(_node_221),
        .a(1'h1),
        .b(_node_220)
    );
    wire [7:0] _GEN_121;
    MUX_UNSIGNED #(.width(8)) u_mux_456 (
        .y(_GEN_121),
        .sel(_node_221),
        .a(helloWorld_111),
        .b(_GEN_120)
    );
    wire _node_222;
    wire [8:0] _WTEMP_113;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_457 (
        .y(_WTEMP_113),
        .in(7'h70)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_458 (
        .y(_node_222),
        .a(_WTEMP_113),
        .b(_arrivedPointer__q)
    );
    wire _node_223;
    BITWISEAND #(.width(1)) bitwiseand_459 (
        .y(_node_223),
        .a(1'h1),
        .b(_node_222)
    );
    wire [7:0] _GEN_122;
    MUX_UNSIGNED #(.width(8)) u_mux_460 (
        .y(_GEN_122),
        .sel(_node_223),
        .a(helloWorld_112),
        .b(_GEN_121)
    );
    wire _node_224;
    wire [8:0] _WTEMP_114;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_461 (
        .y(_WTEMP_114),
        .in(7'h71)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_462 (
        .y(_node_224),
        .a(_WTEMP_114),
        .b(_arrivedPointer__q)
    );
    wire _node_225;
    BITWISEAND #(.width(1)) bitwiseand_463 (
        .y(_node_225),
        .a(1'h1),
        .b(_node_224)
    );
    wire [7:0] _GEN_123;
    MUX_UNSIGNED #(.width(8)) u_mux_464 (
        .y(_GEN_123),
        .sel(_node_225),
        .a(helloWorld_113),
        .b(_GEN_122)
    );
    wire _node_226;
    wire [8:0] _WTEMP_115;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_465 (
        .y(_WTEMP_115),
        .in(7'h72)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_466 (
        .y(_node_226),
        .a(_WTEMP_115),
        .b(_arrivedPointer__q)
    );
    wire _node_227;
    BITWISEAND #(.width(1)) bitwiseand_467 (
        .y(_node_227),
        .a(1'h1),
        .b(_node_226)
    );
    wire [7:0] _GEN_124;
    MUX_UNSIGNED #(.width(8)) u_mux_468 (
        .y(_GEN_124),
        .sel(_node_227),
        .a(helloWorld_114),
        .b(_GEN_123)
    );
    wire _node_228;
    wire [8:0] _WTEMP_116;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_469 (
        .y(_WTEMP_116),
        .in(7'h73)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_470 (
        .y(_node_228),
        .a(_WTEMP_116),
        .b(_arrivedPointer__q)
    );
    wire _node_229;
    BITWISEAND #(.width(1)) bitwiseand_471 (
        .y(_node_229),
        .a(1'h1),
        .b(_node_228)
    );
    wire [7:0] _GEN_125;
    MUX_UNSIGNED #(.width(8)) u_mux_472 (
        .y(_GEN_125),
        .sel(_node_229),
        .a(helloWorld_115),
        .b(_GEN_124)
    );
    wire _node_230;
    wire [8:0] _WTEMP_117;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_473 (
        .y(_WTEMP_117),
        .in(7'h74)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_474 (
        .y(_node_230),
        .a(_WTEMP_117),
        .b(_arrivedPointer__q)
    );
    wire _node_231;
    BITWISEAND #(.width(1)) bitwiseand_475 (
        .y(_node_231),
        .a(1'h1),
        .b(_node_230)
    );
    wire [7:0] _GEN_126;
    MUX_UNSIGNED #(.width(8)) u_mux_476 (
        .y(_GEN_126),
        .sel(_node_231),
        .a(helloWorld_116),
        .b(_GEN_125)
    );
    wire _node_232;
    wire [8:0] _WTEMP_118;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_477 (
        .y(_WTEMP_118),
        .in(7'h75)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_478 (
        .y(_node_232),
        .a(_WTEMP_118),
        .b(_arrivedPointer__q)
    );
    wire _node_233;
    BITWISEAND #(.width(1)) bitwiseand_479 (
        .y(_node_233),
        .a(1'h1),
        .b(_node_232)
    );
    wire [7:0] _GEN_127;
    MUX_UNSIGNED #(.width(8)) u_mux_480 (
        .y(_GEN_127),
        .sel(_node_233),
        .a(helloWorld_117),
        .b(_GEN_126)
    );
    wire _node_234;
    wire [8:0] _WTEMP_119;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_481 (
        .y(_WTEMP_119),
        .in(7'h76)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_482 (
        .y(_node_234),
        .a(_WTEMP_119),
        .b(_arrivedPointer__q)
    );
    wire _node_235;
    BITWISEAND #(.width(1)) bitwiseand_483 (
        .y(_node_235),
        .a(1'h1),
        .b(_node_234)
    );
    wire [7:0] _GEN_128;
    MUX_UNSIGNED #(.width(8)) u_mux_484 (
        .y(_GEN_128),
        .sel(_node_235),
        .a(helloWorld_118),
        .b(_GEN_127)
    );
    wire _node_236;
    wire [8:0] _WTEMP_120;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_485 (
        .y(_WTEMP_120),
        .in(7'h77)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_486 (
        .y(_node_236),
        .a(_WTEMP_120),
        .b(_arrivedPointer__q)
    );
    wire _node_237;
    BITWISEAND #(.width(1)) bitwiseand_487 (
        .y(_node_237),
        .a(1'h1),
        .b(_node_236)
    );
    wire [7:0] _GEN_129;
    MUX_UNSIGNED #(.width(8)) u_mux_488 (
        .y(_GEN_129),
        .sel(_node_237),
        .a(helloWorld_119),
        .b(_GEN_128)
    );
    wire _node_238;
    wire [8:0] _WTEMP_121;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_489 (
        .y(_WTEMP_121),
        .in(7'h78)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_490 (
        .y(_node_238),
        .a(_WTEMP_121),
        .b(_arrivedPointer__q)
    );
    wire _node_239;
    BITWISEAND #(.width(1)) bitwiseand_491 (
        .y(_node_239),
        .a(1'h1),
        .b(_node_238)
    );
    wire [7:0] _GEN_130;
    MUX_UNSIGNED #(.width(8)) u_mux_492 (
        .y(_GEN_130),
        .sel(_node_239),
        .a(helloWorld_120),
        .b(_GEN_129)
    );
    wire _node_240;
    wire [8:0] _WTEMP_122;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_493 (
        .y(_WTEMP_122),
        .in(7'h79)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_494 (
        .y(_node_240),
        .a(_WTEMP_122),
        .b(_arrivedPointer__q)
    );
    wire _node_241;
    BITWISEAND #(.width(1)) bitwiseand_495 (
        .y(_node_241),
        .a(1'h1),
        .b(_node_240)
    );
    wire [7:0] _GEN_131;
    MUX_UNSIGNED #(.width(8)) u_mux_496 (
        .y(_GEN_131),
        .sel(_node_241),
        .a(helloWorld_121),
        .b(_GEN_130)
    );
    wire _node_242;
    wire [8:0] _WTEMP_123;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_497 (
        .y(_WTEMP_123),
        .in(7'h7A)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_498 (
        .y(_node_242),
        .a(_WTEMP_123),
        .b(_arrivedPointer__q)
    );
    wire _node_243;
    BITWISEAND #(.width(1)) bitwiseand_499 (
        .y(_node_243),
        .a(1'h1),
        .b(_node_242)
    );
    wire [7:0] _GEN_132;
    MUX_UNSIGNED #(.width(8)) u_mux_500 (
        .y(_GEN_132),
        .sel(_node_243),
        .a(helloWorld_122),
        .b(_GEN_131)
    );
    wire _node_244;
    wire [8:0] _WTEMP_124;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_501 (
        .y(_WTEMP_124),
        .in(7'h7B)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_502 (
        .y(_node_244),
        .a(_WTEMP_124),
        .b(_arrivedPointer__q)
    );
    wire _node_245;
    BITWISEAND #(.width(1)) bitwiseand_503 (
        .y(_node_245),
        .a(1'h1),
        .b(_node_244)
    );
    wire [7:0] _GEN_133;
    MUX_UNSIGNED #(.width(8)) u_mux_504 (
        .y(_GEN_133),
        .sel(_node_245),
        .a(helloWorld_123),
        .b(_GEN_132)
    );
    wire _node_246;
    wire [8:0] _WTEMP_125;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_505 (
        .y(_WTEMP_125),
        .in(7'h7C)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_506 (
        .y(_node_246),
        .a(_WTEMP_125),
        .b(_arrivedPointer__q)
    );
    wire _node_247;
    BITWISEAND #(.width(1)) bitwiseand_507 (
        .y(_node_247),
        .a(1'h1),
        .b(_node_246)
    );
    wire [7:0] _GEN_134;
    MUX_UNSIGNED #(.width(8)) u_mux_508 (
        .y(_GEN_134),
        .sel(_node_247),
        .a(helloWorld_124),
        .b(_GEN_133)
    );
    wire _node_248;
    wire [8:0] _WTEMP_126;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_509 (
        .y(_WTEMP_126),
        .in(7'h7D)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_510 (
        .y(_node_248),
        .a(_WTEMP_126),
        .b(_arrivedPointer__q)
    );
    wire _node_249;
    BITWISEAND #(.width(1)) bitwiseand_511 (
        .y(_node_249),
        .a(1'h1),
        .b(_node_248)
    );
    wire [7:0] _GEN_135;
    MUX_UNSIGNED #(.width(8)) u_mux_512 (
        .y(_GEN_135),
        .sel(_node_249),
        .a(helloWorld_125),
        .b(_GEN_134)
    );
    wire _node_250;
    wire [8:0] _WTEMP_127;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_513 (
        .y(_WTEMP_127),
        .in(7'h7E)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_514 (
        .y(_node_250),
        .a(_WTEMP_127),
        .b(_arrivedPointer__q)
    );
    wire _node_251;
    BITWISEAND #(.width(1)) bitwiseand_515 (
        .y(_node_251),
        .a(1'h1),
        .b(_node_250)
    );
    wire [7:0] _GEN_136;
    MUX_UNSIGNED #(.width(8)) u_mux_516 (
        .y(_GEN_136),
        .sel(_node_251),
        .a(helloWorld_126),
        .b(_GEN_135)
    );
    wire _node_252;
    wire [8:0] _WTEMP_128;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_517 (
        .y(_WTEMP_128),
        .in(7'h7F)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_518 (
        .y(_node_252),
        .a(_WTEMP_128),
        .b(_arrivedPointer__q)
    );
    wire _node_253;
    BITWISEAND #(.width(1)) bitwiseand_519 (
        .y(_node_253),
        .a(1'h1),
        .b(_node_252)
    );
    wire [7:0] _GEN_137;
    MUX_UNSIGNED #(.width(8)) u_mux_520 (
        .y(_GEN_137),
        .sel(_node_253),
        .a(helloWorld_127),
        .b(_GEN_136)
    );
    wire _node_254;
    wire [8:0] _WTEMP_129;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_521 (
        .y(_WTEMP_129),
        .in(8'h80)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_522 (
        .y(_node_254),
        .a(_WTEMP_129),
        .b(_arrivedPointer__q)
    );
    wire _node_255;
    BITWISEAND #(.width(1)) bitwiseand_523 (
        .y(_node_255),
        .a(1'h1),
        .b(_node_254)
    );
    wire [7:0] _GEN_138;
    MUX_UNSIGNED #(.width(8)) u_mux_524 (
        .y(_GEN_138),
        .sel(_node_255),
        .a(helloWorld_128),
        .b(_GEN_137)
    );
    wire _node_256;
    wire [8:0] _WTEMP_130;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_525 (
        .y(_WTEMP_130),
        .in(8'h81)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_526 (
        .y(_node_256),
        .a(_WTEMP_130),
        .b(_arrivedPointer__q)
    );
    wire _node_257;
    BITWISEAND #(.width(1)) bitwiseand_527 (
        .y(_node_257),
        .a(1'h1),
        .b(_node_256)
    );
    wire [7:0] _GEN_139;
    MUX_UNSIGNED #(.width(8)) u_mux_528 (
        .y(_GEN_139),
        .sel(_node_257),
        .a(helloWorld_129),
        .b(_GEN_138)
    );
    wire _node_258;
    wire [8:0] _WTEMP_131;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_529 (
        .y(_WTEMP_131),
        .in(8'h82)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_530 (
        .y(_node_258),
        .a(_WTEMP_131),
        .b(_arrivedPointer__q)
    );
    wire _node_259;
    BITWISEAND #(.width(1)) bitwiseand_531 (
        .y(_node_259),
        .a(1'h1),
        .b(_node_258)
    );
    wire [7:0] _GEN_140;
    MUX_UNSIGNED #(.width(8)) u_mux_532 (
        .y(_GEN_140),
        .sel(_node_259),
        .a(helloWorld_130),
        .b(_GEN_139)
    );
    wire _node_260;
    wire [8:0] _WTEMP_132;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_533 (
        .y(_WTEMP_132),
        .in(8'h83)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_534 (
        .y(_node_260),
        .a(_WTEMP_132),
        .b(_arrivedPointer__q)
    );
    wire _node_261;
    BITWISEAND #(.width(1)) bitwiseand_535 (
        .y(_node_261),
        .a(1'h1),
        .b(_node_260)
    );
    wire [7:0] _GEN_141;
    MUX_UNSIGNED #(.width(8)) u_mux_536 (
        .y(_GEN_141),
        .sel(_node_261),
        .a(helloWorld_131),
        .b(_GEN_140)
    );
    wire _node_262;
    wire [8:0] _WTEMP_133;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_537 (
        .y(_WTEMP_133),
        .in(8'h84)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_538 (
        .y(_node_262),
        .a(_WTEMP_133),
        .b(_arrivedPointer__q)
    );
    wire _node_263;
    BITWISEAND #(.width(1)) bitwiseand_539 (
        .y(_node_263),
        .a(1'h1),
        .b(_node_262)
    );
    wire [7:0] _GEN_142;
    MUX_UNSIGNED #(.width(8)) u_mux_540 (
        .y(_GEN_142),
        .sel(_node_263),
        .a(helloWorld_132),
        .b(_GEN_141)
    );
    wire _node_264;
    wire [8:0] _WTEMP_134;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_541 (
        .y(_WTEMP_134),
        .in(8'h85)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_542 (
        .y(_node_264),
        .a(_WTEMP_134),
        .b(_arrivedPointer__q)
    );
    wire _node_265;
    BITWISEAND #(.width(1)) bitwiseand_543 (
        .y(_node_265),
        .a(1'h1),
        .b(_node_264)
    );
    wire [7:0] _GEN_143;
    MUX_UNSIGNED #(.width(8)) u_mux_544 (
        .y(_GEN_143),
        .sel(_node_265),
        .a(helloWorld_133),
        .b(_GEN_142)
    );
    wire _node_266;
    wire [8:0] _WTEMP_135;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_545 (
        .y(_WTEMP_135),
        .in(8'h86)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_546 (
        .y(_node_266),
        .a(_WTEMP_135),
        .b(_arrivedPointer__q)
    );
    wire _node_267;
    BITWISEAND #(.width(1)) bitwiseand_547 (
        .y(_node_267),
        .a(1'h1),
        .b(_node_266)
    );
    wire [7:0] _GEN_144;
    MUX_UNSIGNED #(.width(8)) u_mux_548 (
        .y(_GEN_144),
        .sel(_node_267),
        .a(helloWorld_134),
        .b(_GEN_143)
    );
    wire _node_268;
    wire [8:0] _WTEMP_136;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_549 (
        .y(_WTEMP_136),
        .in(8'h87)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_550 (
        .y(_node_268),
        .a(_WTEMP_136),
        .b(_arrivedPointer__q)
    );
    wire _node_269;
    BITWISEAND #(.width(1)) bitwiseand_551 (
        .y(_node_269),
        .a(1'h1),
        .b(_node_268)
    );
    wire [7:0] _GEN_145;
    MUX_UNSIGNED #(.width(8)) u_mux_552 (
        .y(_GEN_145),
        .sel(_node_269),
        .a(helloWorld_135),
        .b(_GEN_144)
    );
    wire _node_270;
    wire [8:0] _WTEMP_137;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_553 (
        .y(_WTEMP_137),
        .in(8'h88)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_554 (
        .y(_node_270),
        .a(_WTEMP_137),
        .b(_arrivedPointer__q)
    );
    wire _node_271;
    BITWISEAND #(.width(1)) bitwiseand_555 (
        .y(_node_271),
        .a(1'h1),
        .b(_node_270)
    );
    wire [7:0] _GEN_146;
    MUX_UNSIGNED #(.width(8)) u_mux_556 (
        .y(_GEN_146),
        .sel(_node_271),
        .a(helloWorld_136),
        .b(_GEN_145)
    );
    wire _node_272;
    wire [8:0] _WTEMP_138;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_557 (
        .y(_WTEMP_138),
        .in(8'h89)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_558 (
        .y(_node_272),
        .a(_WTEMP_138),
        .b(_arrivedPointer__q)
    );
    wire _node_273;
    BITWISEAND #(.width(1)) bitwiseand_559 (
        .y(_node_273),
        .a(1'h1),
        .b(_node_272)
    );
    wire [7:0] _GEN_147;
    MUX_UNSIGNED #(.width(8)) u_mux_560 (
        .y(_GEN_147),
        .sel(_node_273),
        .a(helloWorld_137),
        .b(_GEN_146)
    );
    wire _node_274;
    wire [8:0] _WTEMP_139;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_561 (
        .y(_WTEMP_139),
        .in(8'h8A)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_562 (
        .y(_node_274),
        .a(_WTEMP_139),
        .b(_arrivedPointer__q)
    );
    wire _node_275;
    BITWISEAND #(.width(1)) bitwiseand_563 (
        .y(_node_275),
        .a(1'h1),
        .b(_node_274)
    );
    wire [7:0] _GEN_148;
    MUX_UNSIGNED #(.width(8)) u_mux_564 (
        .y(_GEN_148),
        .sel(_node_275),
        .a(helloWorld_138),
        .b(_GEN_147)
    );
    wire _node_276;
    wire [8:0] _WTEMP_140;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_565 (
        .y(_WTEMP_140),
        .in(8'h8B)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_566 (
        .y(_node_276),
        .a(_WTEMP_140),
        .b(_arrivedPointer__q)
    );
    wire _node_277;
    BITWISEAND #(.width(1)) bitwiseand_567 (
        .y(_node_277),
        .a(1'h1),
        .b(_node_276)
    );
    wire [7:0] _GEN_149;
    MUX_UNSIGNED #(.width(8)) u_mux_568 (
        .y(_GEN_149),
        .sel(_node_277),
        .a(helloWorld_139),
        .b(_GEN_148)
    );
    wire _node_278;
    wire [8:0] _WTEMP_141;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_569 (
        .y(_WTEMP_141),
        .in(8'h8C)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_570 (
        .y(_node_278),
        .a(_WTEMP_141),
        .b(_arrivedPointer__q)
    );
    wire _node_279;
    BITWISEAND #(.width(1)) bitwiseand_571 (
        .y(_node_279),
        .a(1'h1),
        .b(_node_278)
    );
    wire [7:0] _GEN_150;
    MUX_UNSIGNED #(.width(8)) u_mux_572 (
        .y(_GEN_150),
        .sel(_node_279),
        .a(helloWorld_140),
        .b(_GEN_149)
    );
    wire _node_280;
    wire [8:0] _WTEMP_142;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_573 (
        .y(_WTEMP_142),
        .in(8'h8D)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_574 (
        .y(_node_280),
        .a(_WTEMP_142),
        .b(_arrivedPointer__q)
    );
    wire _node_281;
    BITWISEAND #(.width(1)) bitwiseand_575 (
        .y(_node_281),
        .a(1'h1),
        .b(_node_280)
    );
    wire [7:0] _GEN_151;
    MUX_UNSIGNED #(.width(8)) u_mux_576 (
        .y(_GEN_151),
        .sel(_node_281),
        .a(helloWorld_141),
        .b(_GEN_150)
    );
    wire _node_282;
    wire [8:0] _WTEMP_143;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_577 (
        .y(_WTEMP_143),
        .in(8'h8E)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_578 (
        .y(_node_282),
        .a(_WTEMP_143),
        .b(_arrivedPointer__q)
    );
    wire _node_283;
    BITWISEAND #(.width(1)) bitwiseand_579 (
        .y(_node_283),
        .a(1'h1),
        .b(_node_282)
    );
    wire [7:0] _GEN_152;
    MUX_UNSIGNED #(.width(8)) u_mux_580 (
        .y(_GEN_152),
        .sel(_node_283),
        .a(helloWorld_142),
        .b(_GEN_151)
    );
    wire _node_284;
    wire [8:0] _WTEMP_144;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_581 (
        .y(_WTEMP_144),
        .in(8'h8F)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_582 (
        .y(_node_284),
        .a(_WTEMP_144),
        .b(_arrivedPointer__q)
    );
    wire _node_285;
    BITWISEAND #(.width(1)) bitwiseand_583 (
        .y(_node_285),
        .a(1'h1),
        .b(_node_284)
    );
    wire [7:0] _GEN_153;
    MUX_UNSIGNED #(.width(8)) u_mux_584 (
        .y(_GEN_153),
        .sel(_node_285),
        .a(helloWorld_143),
        .b(_GEN_152)
    );
    wire _node_286;
    wire [8:0] _WTEMP_145;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_585 (
        .y(_WTEMP_145),
        .in(8'h90)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_586 (
        .y(_node_286),
        .a(_WTEMP_145),
        .b(_arrivedPointer__q)
    );
    wire _node_287;
    BITWISEAND #(.width(1)) bitwiseand_587 (
        .y(_node_287),
        .a(1'h1),
        .b(_node_286)
    );
    wire [7:0] _GEN_154;
    MUX_UNSIGNED #(.width(8)) u_mux_588 (
        .y(_GEN_154),
        .sel(_node_287),
        .a(helloWorld_144),
        .b(_GEN_153)
    );
    wire _node_288;
    wire [8:0] _WTEMP_146;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_589 (
        .y(_WTEMP_146),
        .in(8'h91)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_590 (
        .y(_node_288),
        .a(_WTEMP_146),
        .b(_arrivedPointer__q)
    );
    wire _node_289;
    BITWISEAND #(.width(1)) bitwiseand_591 (
        .y(_node_289),
        .a(1'h1),
        .b(_node_288)
    );
    wire [7:0] _GEN_155;
    MUX_UNSIGNED #(.width(8)) u_mux_592 (
        .y(_GEN_155),
        .sel(_node_289),
        .a(helloWorld_145),
        .b(_GEN_154)
    );
    wire _node_290;
    wire [8:0] _WTEMP_147;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_593 (
        .y(_WTEMP_147),
        .in(8'h92)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_594 (
        .y(_node_290),
        .a(_WTEMP_147),
        .b(_arrivedPointer__q)
    );
    wire _node_291;
    BITWISEAND #(.width(1)) bitwiseand_595 (
        .y(_node_291),
        .a(1'h1),
        .b(_node_290)
    );
    wire [7:0] _GEN_156;
    MUX_UNSIGNED #(.width(8)) u_mux_596 (
        .y(_GEN_156),
        .sel(_node_291),
        .a(helloWorld_146),
        .b(_GEN_155)
    );
    wire _node_292;
    wire [8:0] _WTEMP_148;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_597 (
        .y(_WTEMP_148),
        .in(8'h93)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_598 (
        .y(_node_292),
        .a(_WTEMP_148),
        .b(_arrivedPointer__q)
    );
    wire _node_293;
    BITWISEAND #(.width(1)) bitwiseand_599 (
        .y(_node_293),
        .a(1'h1),
        .b(_node_292)
    );
    wire [7:0] _GEN_157;
    MUX_UNSIGNED #(.width(8)) u_mux_600 (
        .y(_GEN_157),
        .sel(_node_293),
        .a(helloWorld_147),
        .b(_GEN_156)
    );
    wire _node_294;
    wire [8:0] _WTEMP_149;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_601 (
        .y(_WTEMP_149),
        .in(8'h94)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_602 (
        .y(_node_294),
        .a(_WTEMP_149),
        .b(_arrivedPointer__q)
    );
    wire _node_295;
    BITWISEAND #(.width(1)) bitwiseand_603 (
        .y(_node_295),
        .a(1'h1),
        .b(_node_294)
    );
    wire [7:0] _GEN_158;
    MUX_UNSIGNED #(.width(8)) u_mux_604 (
        .y(_GEN_158),
        .sel(_node_295),
        .a(helloWorld_148),
        .b(_GEN_157)
    );
    wire _node_296;
    wire [8:0] _WTEMP_150;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_605 (
        .y(_WTEMP_150),
        .in(8'h95)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_606 (
        .y(_node_296),
        .a(_WTEMP_150),
        .b(_arrivedPointer__q)
    );
    wire _node_297;
    BITWISEAND #(.width(1)) bitwiseand_607 (
        .y(_node_297),
        .a(1'h1),
        .b(_node_296)
    );
    wire [7:0] _GEN_159;
    MUX_UNSIGNED #(.width(8)) u_mux_608 (
        .y(_GEN_159),
        .sel(_node_297),
        .a(helloWorld_149),
        .b(_GEN_158)
    );
    wire _node_298;
    wire [8:0] _WTEMP_151;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_609 (
        .y(_WTEMP_151),
        .in(8'h96)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_610 (
        .y(_node_298),
        .a(_WTEMP_151),
        .b(_arrivedPointer__q)
    );
    wire _node_299;
    BITWISEAND #(.width(1)) bitwiseand_611 (
        .y(_node_299),
        .a(1'h1),
        .b(_node_298)
    );
    wire [7:0] _GEN_160;
    MUX_UNSIGNED #(.width(8)) u_mux_612 (
        .y(_GEN_160),
        .sel(_node_299),
        .a(helloWorld_150),
        .b(_GEN_159)
    );
    wire _node_300;
    wire [8:0] _WTEMP_152;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_613 (
        .y(_WTEMP_152),
        .in(8'h97)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_614 (
        .y(_node_300),
        .a(_WTEMP_152),
        .b(_arrivedPointer__q)
    );
    wire _node_301;
    BITWISEAND #(.width(1)) bitwiseand_615 (
        .y(_node_301),
        .a(1'h1),
        .b(_node_300)
    );
    wire [7:0] _GEN_161;
    MUX_UNSIGNED #(.width(8)) u_mux_616 (
        .y(_GEN_161),
        .sel(_node_301),
        .a(helloWorld_151),
        .b(_GEN_160)
    );
    wire _node_302;
    wire [8:0] _WTEMP_153;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_617 (
        .y(_WTEMP_153),
        .in(8'h98)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_618 (
        .y(_node_302),
        .a(_WTEMP_153),
        .b(_arrivedPointer__q)
    );
    wire _node_303;
    BITWISEAND #(.width(1)) bitwiseand_619 (
        .y(_node_303),
        .a(1'h1),
        .b(_node_302)
    );
    wire [7:0] _GEN_162;
    MUX_UNSIGNED #(.width(8)) u_mux_620 (
        .y(_GEN_162),
        .sel(_node_303),
        .a(helloWorld_152),
        .b(_GEN_161)
    );
    wire _node_304;
    wire [8:0] _WTEMP_154;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_621 (
        .y(_WTEMP_154),
        .in(8'h99)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_622 (
        .y(_node_304),
        .a(_WTEMP_154),
        .b(_arrivedPointer__q)
    );
    wire _node_305;
    BITWISEAND #(.width(1)) bitwiseand_623 (
        .y(_node_305),
        .a(1'h1),
        .b(_node_304)
    );
    wire [7:0] _GEN_163;
    MUX_UNSIGNED #(.width(8)) u_mux_624 (
        .y(_GEN_163),
        .sel(_node_305),
        .a(helloWorld_153),
        .b(_GEN_162)
    );
    wire _node_306;
    wire [8:0] _WTEMP_155;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_625 (
        .y(_WTEMP_155),
        .in(8'h9A)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_626 (
        .y(_node_306),
        .a(_WTEMP_155),
        .b(_arrivedPointer__q)
    );
    wire _node_307;
    BITWISEAND #(.width(1)) bitwiseand_627 (
        .y(_node_307),
        .a(1'h1),
        .b(_node_306)
    );
    wire [7:0] _GEN_164;
    MUX_UNSIGNED #(.width(8)) u_mux_628 (
        .y(_GEN_164),
        .sel(_node_307),
        .a(helloWorld_154),
        .b(_GEN_163)
    );
    wire _node_308;
    wire [8:0] _WTEMP_156;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_629 (
        .y(_WTEMP_156),
        .in(8'h9B)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_630 (
        .y(_node_308),
        .a(_WTEMP_156),
        .b(_arrivedPointer__q)
    );
    wire _node_309;
    BITWISEAND #(.width(1)) bitwiseand_631 (
        .y(_node_309),
        .a(1'h1),
        .b(_node_308)
    );
    wire [7:0] _GEN_165;
    MUX_UNSIGNED #(.width(8)) u_mux_632 (
        .y(_GEN_165),
        .sel(_node_309),
        .a(helloWorld_155),
        .b(_GEN_164)
    );
    wire _node_310;
    wire [8:0] _WTEMP_157;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_633 (
        .y(_WTEMP_157),
        .in(8'h9C)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_634 (
        .y(_node_310),
        .a(_WTEMP_157),
        .b(_arrivedPointer__q)
    );
    wire _node_311;
    BITWISEAND #(.width(1)) bitwiseand_635 (
        .y(_node_311),
        .a(1'h1),
        .b(_node_310)
    );
    wire [7:0] _GEN_166;
    MUX_UNSIGNED #(.width(8)) u_mux_636 (
        .y(_GEN_166),
        .sel(_node_311),
        .a(helloWorld_156),
        .b(_GEN_165)
    );
    wire _node_312;
    wire [8:0] _WTEMP_158;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_637 (
        .y(_WTEMP_158),
        .in(8'h9D)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_638 (
        .y(_node_312),
        .a(_WTEMP_158),
        .b(_arrivedPointer__q)
    );
    wire _node_313;
    BITWISEAND #(.width(1)) bitwiseand_639 (
        .y(_node_313),
        .a(1'h1),
        .b(_node_312)
    );
    wire [7:0] _GEN_167;
    MUX_UNSIGNED #(.width(8)) u_mux_640 (
        .y(_GEN_167),
        .sel(_node_313),
        .a(helloWorld_157),
        .b(_GEN_166)
    );
    wire _node_314;
    wire [8:0] _WTEMP_159;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_641 (
        .y(_WTEMP_159),
        .in(8'h9E)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_642 (
        .y(_node_314),
        .a(_WTEMP_159),
        .b(_arrivedPointer__q)
    );
    wire _node_315;
    BITWISEAND #(.width(1)) bitwiseand_643 (
        .y(_node_315),
        .a(1'h1),
        .b(_node_314)
    );
    wire [7:0] _GEN_168;
    MUX_UNSIGNED #(.width(8)) u_mux_644 (
        .y(_GEN_168),
        .sel(_node_315),
        .a(helloWorld_158),
        .b(_GEN_167)
    );
    wire _node_316;
    wire [8:0] _WTEMP_160;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_645 (
        .y(_WTEMP_160),
        .in(8'h9F)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_646 (
        .y(_node_316),
        .a(_WTEMP_160),
        .b(_arrivedPointer__q)
    );
    wire _node_317;
    BITWISEAND #(.width(1)) bitwiseand_647 (
        .y(_node_317),
        .a(1'h1),
        .b(_node_316)
    );
    wire [7:0] _GEN_169;
    MUX_UNSIGNED #(.width(8)) u_mux_648 (
        .y(_GEN_169),
        .sel(_node_317),
        .a(helloWorld_159),
        .b(_GEN_168)
    );
    wire _node_318;
    wire [8:0] _WTEMP_161;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_649 (
        .y(_WTEMP_161),
        .in(8'hA0)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_650 (
        .y(_node_318),
        .a(_WTEMP_161),
        .b(_arrivedPointer__q)
    );
    wire _node_319;
    BITWISEAND #(.width(1)) bitwiseand_651 (
        .y(_node_319),
        .a(1'h1),
        .b(_node_318)
    );
    wire [7:0] _GEN_170;
    MUX_UNSIGNED #(.width(8)) u_mux_652 (
        .y(_GEN_170),
        .sel(_node_319),
        .a(helloWorld_160),
        .b(_GEN_169)
    );
    wire _node_320;
    wire [8:0] _WTEMP_162;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_653 (
        .y(_WTEMP_162),
        .in(8'hA1)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_654 (
        .y(_node_320),
        .a(_WTEMP_162),
        .b(_arrivedPointer__q)
    );
    wire _node_321;
    BITWISEAND #(.width(1)) bitwiseand_655 (
        .y(_node_321),
        .a(1'h1),
        .b(_node_320)
    );
    wire [7:0] _GEN_171;
    MUX_UNSIGNED #(.width(8)) u_mux_656 (
        .y(_GEN_171),
        .sel(_node_321),
        .a(helloWorld_161),
        .b(_GEN_170)
    );
    wire _node_322;
    wire [8:0] _WTEMP_163;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_657 (
        .y(_WTEMP_163),
        .in(8'hA2)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_658 (
        .y(_node_322),
        .a(_WTEMP_163),
        .b(_arrivedPointer__q)
    );
    wire _node_323;
    BITWISEAND #(.width(1)) bitwiseand_659 (
        .y(_node_323),
        .a(1'h1),
        .b(_node_322)
    );
    wire [7:0] _GEN_172;
    MUX_UNSIGNED #(.width(8)) u_mux_660 (
        .y(_GEN_172),
        .sel(_node_323),
        .a(helloWorld_162),
        .b(_GEN_171)
    );
    wire _node_324;
    wire [8:0] _WTEMP_164;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_661 (
        .y(_WTEMP_164),
        .in(8'hA3)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_662 (
        .y(_node_324),
        .a(_WTEMP_164),
        .b(_arrivedPointer__q)
    );
    wire _node_325;
    BITWISEAND #(.width(1)) bitwiseand_663 (
        .y(_node_325),
        .a(1'h1),
        .b(_node_324)
    );
    wire [7:0] _GEN_173;
    MUX_UNSIGNED #(.width(8)) u_mux_664 (
        .y(_GEN_173),
        .sel(_node_325),
        .a(helloWorld_163),
        .b(_GEN_172)
    );
    wire _node_326;
    wire [8:0] _WTEMP_165;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_665 (
        .y(_WTEMP_165),
        .in(8'hA4)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_666 (
        .y(_node_326),
        .a(_WTEMP_165),
        .b(_arrivedPointer__q)
    );
    wire _node_327;
    BITWISEAND #(.width(1)) bitwiseand_667 (
        .y(_node_327),
        .a(1'h1),
        .b(_node_326)
    );
    wire [7:0] _GEN_174;
    MUX_UNSIGNED #(.width(8)) u_mux_668 (
        .y(_GEN_174),
        .sel(_node_327),
        .a(helloWorld_164),
        .b(_GEN_173)
    );
    wire _node_328;
    wire [8:0] _WTEMP_166;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_669 (
        .y(_WTEMP_166),
        .in(8'hA5)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_670 (
        .y(_node_328),
        .a(_WTEMP_166),
        .b(_arrivedPointer__q)
    );
    wire _node_329;
    BITWISEAND #(.width(1)) bitwiseand_671 (
        .y(_node_329),
        .a(1'h1),
        .b(_node_328)
    );
    wire [7:0] _GEN_175;
    MUX_UNSIGNED #(.width(8)) u_mux_672 (
        .y(_GEN_175),
        .sel(_node_329),
        .a(helloWorld_165),
        .b(_GEN_174)
    );
    wire _node_330;
    wire [8:0] _WTEMP_167;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_673 (
        .y(_WTEMP_167),
        .in(8'hA6)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_674 (
        .y(_node_330),
        .a(_WTEMP_167),
        .b(_arrivedPointer__q)
    );
    wire _node_331;
    BITWISEAND #(.width(1)) bitwiseand_675 (
        .y(_node_331),
        .a(1'h1),
        .b(_node_330)
    );
    wire [7:0] _GEN_176;
    MUX_UNSIGNED #(.width(8)) u_mux_676 (
        .y(_GEN_176),
        .sel(_node_331),
        .a(helloWorld_166),
        .b(_GEN_175)
    );
    wire _node_332;
    wire [8:0] _WTEMP_168;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_677 (
        .y(_WTEMP_168),
        .in(8'hA7)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_678 (
        .y(_node_332),
        .a(_WTEMP_168),
        .b(_arrivedPointer__q)
    );
    wire _node_333;
    BITWISEAND #(.width(1)) bitwiseand_679 (
        .y(_node_333),
        .a(1'h1),
        .b(_node_332)
    );
    wire [7:0] _GEN_177;
    MUX_UNSIGNED #(.width(8)) u_mux_680 (
        .y(_GEN_177),
        .sel(_node_333),
        .a(helloWorld_167),
        .b(_GEN_176)
    );
    wire _node_334;
    wire [8:0] _WTEMP_169;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_681 (
        .y(_WTEMP_169),
        .in(8'hA8)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_682 (
        .y(_node_334),
        .a(_WTEMP_169),
        .b(_arrivedPointer__q)
    );
    wire _node_335;
    BITWISEAND #(.width(1)) bitwiseand_683 (
        .y(_node_335),
        .a(1'h1),
        .b(_node_334)
    );
    wire [7:0] _GEN_178;
    MUX_UNSIGNED #(.width(8)) u_mux_684 (
        .y(_GEN_178),
        .sel(_node_335),
        .a(helloWorld_168),
        .b(_GEN_177)
    );
    wire _node_336;
    wire [8:0] _WTEMP_170;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_685 (
        .y(_WTEMP_170),
        .in(8'hA9)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_686 (
        .y(_node_336),
        .a(_WTEMP_170),
        .b(_arrivedPointer__q)
    );
    wire _node_337;
    BITWISEAND #(.width(1)) bitwiseand_687 (
        .y(_node_337),
        .a(1'h1),
        .b(_node_336)
    );
    wire [7:0] _GEN_179;
    MUX_UNSIGNED #(.width(8)) u_mux_688 (
        .y(_GEN_179),
        .sel(_node_337),
        .a(helloWorld_169),
        .b(_GEN_178)
    );
    wire _node_338;
    wire [8:0] _WTEMP_171;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_689 (
        .y(_WTEMP_171),
        .in(8'hAA)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_690 (
        .y(_node_338),
        .a(_WTEMP_171),
        .b(_arrivedPointer__q)
    );
    wire _node_339;
    BITWISEAND #(.width(1)) bitwiseand_691 (
        .y(_node_339),
        .a(1'h1),
        .b(_node_338)
    );
    wire [7:0] _GEN_180;
    MUX_UNSIGNED #(.width(8)) u_mux_692 (
        .y(_GEN_180),
        .sel(_node_339),
        .a(helloWorld_170),
        .b(_GEN_179)
    );
    wire _node_340;
    wire [8:0] _WTEMP_172;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_693 (
        .y(_WTEMP_172),
        .in(8'hAB)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_694 (
        .y(_node_340),
        .a(_WTEMP_172),
        .b(_arrivedPointer__q)
    );
    wire _node_341;
    BITWISEAND #(.width(1)) bitwiseand_695 (
        .y(_node_341),
        .a(1'h1),
        .b(_node_340)
    );
    wire [7:0] _GEN_181;
    MUX_UNSIGNED #(.width(8)) u_mux_696 (
        .y(_GEN_181),
        .sel(_node_341),
        .a(helloWorld_171),
        .b(_GEN_180)
    );
    wire _node_342;
    wire [8:0] _WTEMP_173;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_697 (
        .y(_WTEMP_173),
        .in(8'hAC)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_698 (
        .y(_node_342),
        .a(_WTEMP_173),
        .b(_arrivedPointer__q)
    );
    wire _node_343;
    BITWISEAND #(.width(1)) bitwiseand_699 (
        .y(_node_343),
        .a(1'h1),
        .b(_node_342)
    );
    wire [7:0] _GEN_182;
    MUX_UNSIGNED #(.width(8)) u_mux_700 (
        .y(_GEN_182),
        .sel(_node_343),
        .a(helloWorld_172),
        .b(_GEN_181)
    );
    wire _node_344;
    wire [8:0] _WTEMP_174;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_701 (
        .y(_WTEMP_174),
        .in(8'hAD)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_702 (
        .y(_node_344),
        .a(_WTEMP_174),
        .b(_arrivedPointer__q)
    );
    wire _node_345;
    BITWISEAND #(.width(1)) bitwiseand_703 (
        .y(_node_345),
        .a(1'h1),
        .b(_node_344)
    );
    wire [7:0] _GEN_183;
    MUX_UNSIGNED #(.width(8)) u_mux_704 (
        .y(_GEN_183),
        .sel(_node_345),
        .a(helloWorld_173),
        .b(_GEN_182)
    );
    wire _node_346;
    wire [8:0] _WTEMP_175;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_705 (
        .y(_WTEMP_175),
        .in(8'hAE)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_706 (
        .y(_node_346),
        .a(_WTEMP_175),
        .b(_arrivedPointer__q)
    );
    wire _node_347;
    BITWISEAND #(.width(1)) bitwiseand_707 (
        .y(_node_347),
        .a(1'h1),
        .b(_node_346)
    );
    wire [7:0] _GEN_184;
    MUX_UNSIGNED #(.width(8)) u_mux_708 (
        .y(_GEN_184),
        .sel(_node_347),
        .a(helloWorld_174),
        .b(_GEN_183)
    );
    wire _node_348;
    wire [8:0] _WTEMP_176;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_709 (
        .y(_WTEMP_176),
        .in(8'hAF)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_710 (
        .y(_node_348),
        .a(_WTEMP_176),
        .b(_arrivedPointer__q)
    );
    wire _node_349;
    BITWISEAND #(.width(1)) bitwiseand_711 (
        .y(_node_349),
        .a(1'h1),
        .b(_node_348)
    );
    wire [7:0] _GEN_185;
    MUX_UNSIGNED #(.width(8)) u_mux_712 (
        .y(_GEN_185),
        .sel(_node_349),
        .a(helloWorld_175),
        .b(_GEN_184)
    );
    wire _node_350;
    wire [8:0] _WTEMP_177;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_713 (
        .y(_WTEMP_177),
        .in(8'hB0)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_714 (
        .y(_node_350),
        .a(_WTEMP_177),
        .b(_arrivedPointer__q)
    );
    wire _node_351;
    BITWISEAND #(.width(1)) bitwiseand_715 (
        .y(_node_351),
        .a(1'h1),
        .b(_node_350)
    );
    wire [7:0] _GEN_186;
    MUX_UNSIGNED #(.width(8)) u_mux_716 (
        .y(_GEN_186),
        .sel(_node_351),
        .a(helloWorld_176),
        .b(_GEN_185)
    );
    wire _node_352;
    wire [8:0] _WTEMP_178;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_717 (
        .y(_WTEMP_178),
        .in(8'hB1)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_718 (
        .y(_node_352),
        .a(_WTEMP_178),
        .b(_arrivedPointer__q)
    );
    wire _node_353;
    BITWISEAND #(.width(1)) bitwiseand_719 (
        .y(_node_353),
        .a(1'h1),
        .b(_node_352)
    );
    wire [7:0] _GEN_187;
    MUX_UNSIGNED #(.width(8)) u_mux_720 (
        .y(_GEN_187),
        .sel(_node_353),
        .a(helloWorld_177),
        .b(_GEN_186)
    );
    wire _node_354;
    wire [8:0] _WTEMP_179;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_721 (
        .y(_WTEMP_179),
        .in(8'hB2)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_722 (
        .y(_node_354),
        .a(_WTEMP_179),
        .b(_arrivedPointer__q)
    );
    wire _node_355;
    BITWISEAND #(.width(1)) bitwiseand_723 (
        .y(_node_355),
        .a(1'h1),
        .b(_node_354)
    );
    wire [7:0] _GEN_188;
    MUX_UNSIGNED #(.width(8)) u_mux_724 (
        .y(_GEN_188),
        .sel(_node_355),
        .a(helloWorld_178),
        .b(_GEN_187)
    );
    wire _node_356;
    wire [8:0] _WTEMP_180;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_725 (
        .y(_WTEMP_180),
        .in(8'hB3)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_726 (
        .y(_node_356),
        .a(_WTEMP_180),
        .b(_arrivedPointer__q)
    );
    wire _node_357;
    BITWISEAND #(.width(1)) bitwiseand_727 (
        .y(_node_357),
        .a(1'h1),
        .b(_node_356)
    );
    wire [7:0] _GEN_189;
    MUX_UNSIGNED #(.width(8)) u_mux_728 (
        .y(_GEN_189),
        .sel(_node_357),
        .a(helloWorld_179),
        .b(_GEN_188)
    );
    wire _node_358;
    wire [8:0] _WTEMP_181;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_729 (
        .y(_WTEMP_181),
        .in(8'hB4)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_730 (
        .y(_node_358),
        .a(_WTEMP_181),
        .b(_arrivedPointer__q)
    );
    wire _node_359;
    BITWISEAND #(.width(1)) bitwiseand_731 (
        .y(_node_359),
        .a(1'h1),
        .b(_node_358)
    );
    wire [7:0] _GEN_190;
    MUX_UNSIGNED #(.width(8)) u_mux_732 (
        .y(_GEN_190),
        .sel(_node_359),
        .a(helloWorld_180),
        .b(_GEN_189)
    );
    wire _node_360;
    wire [8:0] _WTEMP_182;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_733 (
        .y(_WTEMP_182),
        .in(8'hB5)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_734 (
        .y(_node_360),
        .a(_WTEMP_182),
        .b(_arrivedPointer__q)
    );
    wire _node_361;
    BITWISEAND #(.width(1)) bitwiseand_735 (
        .y(_node_361),
        .a(1'h1),
        .b(_node_360)
    );
    wire [7:0] _GEN_191;
    MUX_UNSIGNED #(.width(8)) u_mux_736 (
        .y(_GEN_191),
        .sel(_node_361),
        .a(helloWorld_181),
        .b(_GEN_190)
    );
    wire _node_362;
    wire [8:0] _WTEMP_183;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_737 (
        .y(_WTEMP_183),
        .in(8'hB6)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_738 (
        .y(_node_362),
        .a(_WTEMP_183),
        .b(_arrivedPointer__q)
    );
    wire _node_363;
    BITWISEAND #(.width(1)) bitwiseand_739 (
        .y(_node_363),
        .a(1'h1),
        .b(_node_362)
    );
    wire [7:0] _GEN_192;
    MUX_UNSIGNED #(.width(8)) u_mux_740 (
        .y(_GEN_192),
        .sel(_node_363),
        .a(helloWorld_182),
        .b(_GEN_191)
    );
    wire _node_364;
    wire [8:0] _WTEMP_184;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_741 (
        .y(_WTEMP_184),
        .in(8'hB7)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_742 (
        .y(_node_364),
        .a(_WTEMP_184),
        .b(_arrivedPointer__q)
    );
    wire _node_365;
    BITWISEAND #(.width(1)) bitwiseand_743 (
        .y(_node_365),
        .a(1'h1),
        .b(_node_364)
    );
    wire [7:0] _GEN_193;
    MUX_UNSIGNED #(.width(8)) u_mux_744 (
        .y(_GEN_193),
        .sel(_node_365),
        .a(helloWorld_183),
        .b(_GEN_192)
    );
    wire _node_366;
    wire [8:0] _WTEMP_185;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_745 (
        .y(_WTEMP_185),
        .in(8'hB8)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_746 (
        .y(_node_366),
        .a(_WTEMP_185),
        .b(_arrivedPointer__q)
    );
    wire _node_367;
    BITWISEAND #(.width(1)) bitwiseand_747 (
        .y(_node_367),
        .a(1'h1),
        .b(_node_366)
    );
    wire [7:0] _GEN_194;
    MUX_UNSIGNED #(.width(8)) u_mux_748 (
        .y(_GEN_194),
        .sel(_node_367),
        .a(helloWorld_184),
        .b(_GEN_193)
    );
    wire _node_368;
    wire [8:0] _WTEMP_186;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_749 (
        .y(_WTEMP_186),
        .in(8'hB9)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_750 (
        .y(_node_368),
        .a(_WTEMP_186),
        .b(_arrivedPointer__q)
    );
    wire _node_369;
    BITWISEAND #(.width(1)) bitwiseand_751 (
        .y(_node_369),
        .a(1'h1),
        .b(_node_368)
    );
    wire [7:0] _GEN_195;
    MUX_UNSIGNED #(.width(8)) u_mux_752 (
        .y(_GEN_195),
        .sel(_node_369),
        .a(helloWorld_185),
        .b(_GEN_194)
    );
    wire _node_370;
    wire [8:0] _WTEMP_187;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_753 (
        .y(_WTEMP_187),
        .in(8'hBA)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_754 (
        .y(_node_370),
        .a(_WTEMP_187),
        .b(_arrivedPointer__q)
    );
    wire _node_371;
    BITWISEAND #(.width(1)) bitwiseand_755 (
        .y(_node_371),
        .a(1'h1),
        .b(_node_370)
    );
    wire [7:0] _GEN_196;
    MUX_UNSIGNED #(.width(8)) u_mux_756 (
        .y(_GEN_196),
        .sel(_node_371),
        .a(helloWorld_186),
        .b(_GEN_195)
    );
    wire _node_372;
    wire [8:0] _WTEMP_188;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_757 (
        .y(_WTEMP_188),
        .in(8'hBB)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_758 (
        .y(_node_372),
        .a(_WTEMP_188),
        .b(_arrivedPointer__q)
    );
    wire _node_373;
    BITWISEAND #(.width(1)) bitwiseand_759 (
        .y(_node_373),
        .a(1'h1),
        .b(_node_372)
    );
    wire [7:0] _GEN_197;
    MUX_UNSIGNED #(.width(8)) u_mux_760 (
        .y(_GEN_197),
        .sel(_node_373),
        .a(helloWorld_187),
        .b(_GEN_196)
    );
    wire _node_374;
    wire [8:0] _WTEMP_189;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_761 (
        .y(_WTEMP_189),
        .in(8'hBC)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_762 (
        .y(_node_374),
        .a(_WTEMP_189),
        .b(_arrivedPointer__q)
    );
    wire _node_375;
    BITWISEAND #(.width(1)) bitwiseand_763 (
        .y(_node_375),
        .a(1'h1),
        .b(_node_374)
    );
    wire [7:0] _GEN_198;
    MUX_UNSIGNED #(.width(8)) u_mux_764 (
        .y(_GEN_198),
        .sel(_node_375),
        .a(helloWorld_188),
        .b(_GEN_197)
    );
    wire _node_376;
    wire [8:0] _WTEMP_190;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_765 (
        .y(_WTEMP_190),
        .in(8'hBD)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_766 (
        .y(_node_376),
        .a(_WTEMP_190),
        .b(_arrivedPointer__q)
    );
    wire _node_377;
    BITWISEAND #(.width(1)) bitwiseand_767 (
        .y(_node_377),
        .a(1'h1),
        .b(_node_376)
    );
    wire [7:0] _GEN_199;
    MUX_UNSIGNED #(.width(8)) u_mux_768 (
        .y(_GEN_199),
        .sel(_node_377),
        .a(helloWorld_189),
        .b(_GEN_198)
    );
    wire _node_378;
    wire [8:0] _WTEMP_191;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_769 (
        .y(_WTEMP_191),
        .in(8'hBE)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_770 (
        .y(_node_378),
        .a(_WTEMP_191),
        .b(_arrivedPointer__q)
    );
    wire _node_379;
    BITWISEAND #(.width(1)) bitwiseand_771 (
        .y(_node_379),
        .a(1'h1),
        .b(_node_378)
    );
    wire [7:0] _GEN_200;
    MUX_UNSIGNED #(.width(8)) u_mux_772 (
        .y(_GEN_200),
        .sel(_node_379),
        .a(helloWorld_190),
        .b(_GEN_199)
    );
    wire _node_380;
    wire [8:0] _WTEMP_192;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_773 (
        .y(_WTEMP_192),
        .in(8'hBF)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_774 (
        .y(_node_380),
        .a(_WTEMP_192),
        .b(_arrivedPointer__q)
    );
    wire _node_381;
    BITWISEAND #(.width(1)) bitwiseand_775 (
        .y(_node_381),
        .a(1'h1),
        .b(_node_380)
    );
    wire [7:0] _GEN_201;
    MUX_UNSIGNED #(.width(8)) u_mux_776 (
        .y(_GEN_201),
        .sel(_node_381),
        .a(helloWorld_191),
        .b(_GEN_200)
    );
    wire _node_382;
    wire [8:0] _WTEMP_193;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_777 (
        .y(_WTEMP_193),
        .in(8'hC0)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_778 (
        .y(_node_382),
        .a(_WTEMP_193),
        .b(_arrivedPointer__q)
    );
    wire _node_383;
    BITWISEAND #(.width(1)) bitwiseand_779 (
        .y(_node_383),
        .a(1'h1),
        .b(_node_382)
    );
    wire [7:0] _GEN_202;
    MUX_UNSIGNED #(.width(8)) u_mux_780 (
        .y(_GEN_202),
        .sel(_node_383),
        .a(helloWorld_192),
        .b(_GEN_201)
    );
    wire _node_384;
    wire [8:0] _WTEMP_194;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_781 (
        .y(_WTEMP_194),
        .in(8'hC1)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_782 (
        .y(_node_384),
        .a(_WTEMP_194),
        .b(_arrivedPointer__q)
    );
    wire _node_385;
    BITWISEAND #(.width(1)) bitwiseand_783 (
        .y(_node_385),
        .a(1'h1),
        .b(_node_384)
    );
    wire [7:0] _GEN_203;
    MUX_UNSIGNED #(.width(8)) u_mux_784 (
        .y(_GEN_203),
        .sel(_node_385),
        .a(helloWorld_193),
        .b(_GEN_202)
    );
    wire _node_386;
    wire [8:0] _WTEMP_195;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_785 (
        .y(_WTEMP_195),
        .in(8'hC2)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_786 (
        .y(_node_386),
        .a(_WTEMP_195),
        .b(_arrivedPointer__q)
    );
    wire _node_387;
    BITWISEAND #(.width(1)) bitwiseand_787 (
        .y(_node_387),
        .a(1'h1),
        .b(_node_386)
    );
    wire [7:0] _GEN_204;
    MUX_UNSIGNED #(.width(8)) u_mux_788 (
        .y(_GEN_204),
        .sel(_node_387),
        .a(helloWorld_194),
        .b(_GEN_203)
    );
    wire _node_388;
    wire [8:0] _WTEMP_196;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_789 (
        .y(_WTEMP_196),
        .in(8'hC3)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_790 (
        .y(_node_388),
        .a(_WTEMP_196),
        .b(_arrivedPointer__q)
    );
    wire _node_389;
    BITWISEAND #(.width(1)) bitwiseand_791 (
        .y(_node_389),
        .a(1'h1),
        .b(_node_388)
    );
    wire [7:0] _GEN_205;
    MUX_UNSIGNED #(.width(8)) u_mux_792 (
        .y(_GEN_205),
        .sel(_node_389),
        .a(helloWorld_195),
        .b(_GEN_204)
    );
    wire _node_390;
    wire [8:0] _WTEMP_197;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_793 (
        .y(_WTEMP_197),
        .in(8'hC4)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_794 (
        .y(_node_390),
        .a(_WTEMP_197),
        .b(_arrivedPointer__q)
    );
    wire _node_391;
    BITWISEAND #(.width(1)) bitwiseand_795 (
        .y(_node_391),
        .a(1'h1),
        .b(_node_390)
    );
    wire [7:0] _GEN_206;
    MUX_UNSIGNED #(.width(8)) u_mux_796 (
        .y(_GEN_206),
        .sel(_node_391),
        .a(helloWorld_196),
        .b(_GEN_205)
    );
    wire _node_392;
    wire [8:0] _WTEMP_198;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_797 (
        .y(_WTEMP_198),
        .in(8'hC5)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_798 (
        .y(_node_392),
        .a(_WTEMP_198),
        .b(_arrivedPointer__q)
    );
    wire _node_393;
    BITWISEAND #(.width(1)) bitwiseand_799 (
        .y(_node_393),
        .a(1'h1),
        .b(_node_392)
    );
    wire [7:0] _GEN_207;
    MUX_UNSIGNED #(.width(8)) u_mux_800 (
        .y(_GEN_207),
        .sel(_node_393),
        .a(helloWorld_197),
        .b(_GEN_206)
    );
    wire _node_394;
    wire [8:0] _WTEMP_199;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_801 (
        .y(_WTEMP_199),
        .in(8'hC6)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_802 (
        .y(_node_394),
        .a(_WTEMP_199),
        .b(_arrivedPointer__q)
    );
    wire _node_395;
    BITWISEAND #(.width(1)) bitwiseand_803 (
        .y(_node_395),
        .a(1'h1),
        .b(_node_394)
    );
    wire [7:0] _GEN_208;
    MUX_UNSIGNED #(.width(8)) u_mux_804 (
        .y(_GEN_208),
        .sel(_node_395),
        .a(helloWorld_198),
        .b(_GEN_207)
    );
    wire _node_396;
    wire [8:0] _WTEMP_200;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_805 (
        .y(_WTEMP_200),
        .in(8'hC7)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_806 (
        .y(_node_396),
        .a(_WTEMP_200),
        .b(_arrivedPointer__q)
    );
    wire _node_397;
    BITWISEAND #(.width(1)) bitwiseand_807 (
        .y(_node_397),
        .a(1'h1),
        .b(_node_396)
    );
    wire [7:0] _GEN_209;
    MUX_UNSIGNED #(.width(8)) u_mux_808 (
        .y(_GEN_209),
        .sel(_node_397),
        .a(helloWorld_199),
        .b(_GEN_208)
    );
    wire _node_398;
    wire [8:0] _WTEMP_201;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_809 (
        .y(_WTEMP_201),
        .in(8'hC8)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_810 (
        .y(_node_398),
        .a(_WTEMP_201),
        .b(_arrivedPointer__q)
    );
    wire _node_399;
    BITWISEAND #(.width(1)) bitwiseand_811 (
        .y(_node_399),
        .a(1'h1),
        .b(_node_398)
    );
    wire [7:0] _GEN_210;
    MUX_UNSIGNED #(.width(8)) u_mux_812 (
        .y(_GEN_210),
        .sel(_node_399),
        .a(helloWorld_200),
        .b(_GEN_209)
    );
    wire _node_400;
    wire [8:0] _WTEMP_202;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_813 (
        .y(_WTEMP_202),
        .in(8'hC9)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_814 (
        .y(_node_400),
        .a(_WTEMP_202),
        .b(_arrivedPointer__q)
    );
    wire _node_401;
    BITWISEAND #(.width(1)) bitwiseand_815 (
        .y(_node_401),
        .a(1'h1),
        .b(_node_400)
    );
    wire [7:0] _GEN_211;
    MUX_UNSIGNED #(.width(8)) u_mux_816 (
        .y(_GEN_211),
        .sel(_node_401),
        .a(helloWorld_201),
        .b(_GEN_210)
    );
    wire _node_402;
    wire [8:0] _WTEMP_203;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_817 (
        .y(_WTEMP_203),
        .in(8'hCA)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_818 (
        .y(_node_402),
        .a(_WTEMP_203),
        .b(_arrivedPointer__q)
    );
    wire _node_403;
    BITWISEAND #(.width(1)) bitwiseand_819 (
        .y(_node_403),
        .a(1'h1),
        .b(_node_402)
    );
    wire [7:0] _GEN_212;
    MUX_UNSIGNED #(.width(8)) u_mux_820 (
        .y(_GEN_212),
        .sel(_node_403),
        .a(helloWorld_202),
        .b(_GEN_211)
    );
    wire _node_404;
    wire [8:0] _WTEMP_204;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_821 (
        .y(_WTEMP_204),
        .in(8'hCB)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_822 (
        .y(_node_404),
        .a(_WTEMP_204),
        .b(_arrivedPointer__q)
    );
    wire _node_405;
    BITWISEAND #(.width(1)) bitwiseand_823 (
        .y(_node_405),
        .a(1'h1),
        .b(_node_404)
    );
    wire [7:0] _GEN_213;
    MUX_UNSIGNED #(.width(8)) u_mux_824 (
        .y(_GEN_213),
        .sel(_node_405),
        .a(helloWorld_203),
        .b(_GEN_212)
    );
    wire _node_406;
    wire [8:0] _WTEMP_205;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_825 (
        .y(_WTEMP_205),
        .in(8'hCC)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_826 (
        .y(_node_406),
        .a(_WTEMP_205),
        .b(_arrivedPointer__q)
    );
    wire _node_407;
    BITWISEAND #(.width(1)) bitwiseand_827 (
        .y(_node_407),
        .a(1'h1),
        .b(_node_406)
    );
    wire [7:0] _GEN_214;
    MUX_UNSIGNED #(.width(8)) u_mux_828 (
        .y(_GEN_214),
        .sel(_node_407),
        .a(helloWorld_204),
        .b(_GEN_213)
    );
    wire _node_408;
    wire [8:0] _WTEMP_206;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_829 (
        .y(_WTEMP_206),
        .in(8'hCD)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_830 (
        .y(_node_408),
        .a(_WTEMP_206),
        .b(_arrivedPointer__q)
    );
    wire _node_409;
    BITWISEAND #(.width(1)) bitwiseand_831 (
        .y(_node_409),
        .a(1'h1),
        .b(_node_408)
    );
    wire [7:0] _GEN_215;
    MUX_UNSIGNED #(.width(8)) u_mux_832 (
        .y(_GEN_215),
        .sel(_node_409),
        .a(helloWorld_205),
        .b(_GEN_214)
    );
    wire _node_410;
    wire [8:0] _WTEMP_207;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_833 (
        .y(_WTEMP_207),
        .in(8'hCE)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_834 (
        .y(_node_410),
        .a(_WTEMP_207),
        .b(_arrivedPointer__q)
    );
    wire _node_411;
    BITWISEAND #(.width(1)) bitwiseand_835 (
        .y(_node_411),
        .a(1'h1),
        .b(_node_410)
    );
    wire [7:0] _GEN_216;
    MUX_UNSIGNED #(.width(8)) u_mux_836 (
        .y(_GEN_216),
        .sel(_node_411),
        .a(helloWorld_206),
        .b(_GEN_215)
    );
    wire _node_412;
    wire [8:0] _WTEMP_208;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_837 (
        .y(_WTEMP_208),
        .in(8'hCF)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_838 (
        .y(_node_412),
        .a(_WTEMP_208),
        .b(_arrivedPointer__q)
    );
    wire _node_413;
    BITWISEAND #(.width(1)) bitwiseand_839 (
        .y(_node_413),
        .a(1'h1),
        .b(_node_412)
    );
    wire [7:0] _GEN_217;
    MUX_UNSIGNED #(.width(8)) u_mux_840 (
        .y(_GEN_217),
        .sel(_node_413),
        .a(helloWorld_207),
        .b(_GEN_216)
    );
    wire _node_414;
    wire [8:0] _WTEMP_209;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_841 (
        .y(_WTEMP_209),
        .in(8'hD0)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_842 (
        .y(_node_414),
        .a(_WTEMP_209),
        .b(_arrivedPointer__q)
    );
    wire _node_415;
    BITWISEAND #(.width(1)) bitwiseand_843 (
        .y(_node_415),
        .a(1'h1),
        .b(_node_414)
    );
    wire [7:0] _GEN_218;
    MUX_UNSIGNED #(.width(8)) u_mux_844 (
        .y(_GEN_218),
        .sel(_node_415),
        .a(helloWorld_208),
        .b(_GEN_217)
    );
    wire _node_416;
    wire [8:0] _WTEMP_210;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_845 (
        .y(_WTEMP_210),
        .in(8'hD1)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_846 (
        .y(_node_416),
        .a(_WTEMP_210),
        .b(_arrivedPointer__q)
    );
    wire _node_417;
    BITWISEAND #(.width(1)) bitwiseand_847 (
        .y(_node_417),
        .a(1'h1),
        .b(_node_416)
    );
    wire [7:0] _GEN_219;
    MUX_UNSIGNED #(.width(8)) u_mux_848 (
        .y(_GEN_219),
        .sel(_node_417),
        .a(helloWorld_209),
        .b(_GEN_218)
    );
    wire _node_418;
    wire [8:0] _WTEMP_211;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_849 (
        .y(_WTEMP_211),
        .in(8'hD2)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_850 (
        .y(_node_418),
        .a(_WTEMP_211),
        .b(_arrivedPointer__q)
    );
    wire _node_419;
    BITWISEAND #(.width(1)) bitwiseand_851 (
        .y(_node_419),
        .a(1'h1),
        .b(_node_418)
    );
    wire [7:0] _GEN_220;
    MUX_UNSIGNED #(.width(8)) u_mux_852 (
        .y(_GEN_220),
        .sel(_node_419),
        .a(helloWorld_210),
        .b(_GEN_219)
    );
    wire _node_420;
    wire [8:0] _WTEMP_212;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_853 (
        .y(_WTEMP_212),
        .in(8'hD3)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_854 (
        .y(_node_420),
        .a(_WTEMP_212),
        .b(_arrivedPointer__q)
    );
    wire _node_421;
    BITWISEAND #(.width(1)) bitwiseand_855 (
        .y(_node_421),
        .a(1'h1),
        .b(_node_420)
    );
    wire [7:0] _GEN_221;
    MUX_UNSIGNED #(.width(8)) u_mux_856 (
        .y(_GEN_221),
        .sel(_node_421),
        .a(helloWorld_211),
        .b(_GEN_220)
    );
    wire _node_422;
    wire [8:0] _WTEMP_213;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_857 (
        .y(_WTEMP_213),
        .in(8'hD4)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_858 (
        .y(_node_422),
        .a(_WTEMP_213),
        .b(_arrivedPointer__q)
    );
    wire _node_423;
    BITWISEAND #(.width(1)) bitwiseand_859 (
        .y(_node_423),
        .a(1'h1),
        .b(_node_422)
    );
    wire [7:0] _GEN_222;
    MUX_UNSIGNED #(.width(8)) u_mux_860 (
        .y(_GEN_222),
        .sel(_node_423),
        .a(helloWorld_212),
        .b(_GEN_221)
    );
    wire _node_424;
    wire [8:0] _WTEMP_214;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_861 (
        .y(_WTEMP_214),
        .in(8'hD5)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_862 (
        .y(_node_424),
        .a(_WTEMP_214),
        .b(_arrivedPointer__q)
    );
    wire _node_425;
    BITWISEAND #(.width(1)) bitwiseand_863 (
        .y(_node_425),
        .a(1'h1),
        .b(_node_424)
    );
    wire [7:0] _GEN_223;
    MUX_UNSIGNED #(.width(8)) u_mux_864 (
        .y(_GEN_223),
        .sel(_node_425),
        .a(helloWorld_213),
        .b(_GEN_222)
    );
    wire _node_426;
    wire [8:0] _WTEMP_215;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_865 (
        .y(_WTEMP_215),
        .in(8'hD6)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_866 (
        .y(_node_426),
        .a(_WTEMP_215),
        .b(_arrivedPointer__q)
    );
    wire _node_427;
    BITWISEAND #(.width(1)) bitwiseand_867 (
        .y(_node_427),
        .a(1'h1),
        .b(_node_426)
    );
    wire [7:0] _GEN_224;
    MUX_UNSIGNED #(.width(8)) u_mux_868 (
        .y(_GEN_224),
        .sel(_node_427),
        .a(helloWorld_214),
        .b(_GEN_223)
    );
    wire _node_428;
    wire [8:0] _WTEMP_216;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_869 (
        .y(_WTEMP_216),
        .in(8'hD7)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_870 (
        .y(_node_428),
        .a(_WTEMP_216),
        .b(_arrivedPointer__q)
    );
    wire _node_429;
    BITWISEAND #(.width(1)) bitwiseand_871 (
        .y(_node_429),
        .a(1'h1),
        .b(_node_428)
    );
    wire [7:0] _GEN_225;
    MUX_UNSIGNED #(.width(8)) u_mux_872 (
        .y(_GEN_225),
        .sel(_node_429),
        .a(helloWorld_215),
        .b(_GEN_224)
    );
    wire _node_430;
    wire [8:0] _WTEMP_217;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_873 (
        .y(_WTEMP_217),
        .in(8'hD8)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_874 (
        .y(_node_430),
        .a(_WTEMP_217),
        .b(_arrivedPointer__q)
    );
    wire _node_431;
    BITWISEAND #(.width(1)) bitwiseand_875 (
        .y(_node_431),
        .a(1'h1),
        .b(_node_430)
    );
    wire [7:0] _GEN_226;
    MUX_UNSIGNED #(.width(8)) u_mux_876 (
        .y(_GEN_226),
        .sel(_node_431),
        .a(helloWorld_216),
        .b(_GEN_225)
    );
    wire _node_432;
    wire [8:0] _WTEMP_218;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_877 (
        .y(_WTEMP_218),
        .in(8'hD9)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_878 (
        .y(_node_432),
        .a(_WTEMP_218),
        .b(_arrivedPointer__q)
    );
    wire _node_433;
    BITWISEAND #(.width(1)) bitwiseand_879 (
        .y(_node_433),
        .a(1'h1),
        .b(_node_432)
    );
    wire [7:0] _GEN_227;
    MUX_UNSIGNED #(.width(8)) u_mux_880 (
        .y(_GEN_227),
        .sel(_node_433),
        .a(helloWorld_217),
        .b(_GEN_226)
    );
    wire _node_434;
    wire [8:0] _WTEMP_219;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_881 (
        .y(_WTEMP_219),
        .in(8'hDA)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_882 (
        .y(_node_434),
        .a(_WTEMP_219),
        .b(_arrivedPointer__q)
    );
    wire _node_435;
    BITWISEAND #(.width(1)) bitwiseand_883 (
        .y(_node_435),
        .a(1'h1),
        .b(_node_434)
    );
    wire [7:0] _GEN_228;
    MUX_UNSIGNED #(.width(8)) u_mux_884 (
        .y(_GEN_228),
        .sel(_node_435),
        .a(helloWorld_218),
        .b(_GEN_227)
    );
    wire _node_436;
    wire [8:0] _WTEMP_220;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_885 (
        .y(_WTEMP_220),
        .in(8'hDB)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_886 (
        .y(_node_436),
        .a(_WTEMP_220),
        .b(_arrivedPointer__q)
    );
    wire _node_437;
    BITWISEAND #(.width(1)) bitwiseand_887 (
        .y(_node_437),
        .a(1'h1),
        .b(_node_436)
    );
    wire [7:0] _GEN_229;
    MUX_UNSIGNED #(.width(8)) u_mux_888 (
        .y(_GEN_229),
        .sel(_node_437),
        .a(helloWorld_219),
        .b(_GEN_228)
    );
    wire _node_438;
    wire [8:0] _WTEMP_221;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_889 (
        .y(_WTEMP_221),
        .in(8'hDC)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_890 (
        .y(_node_438),
        .a(_WTEMP_221),
        .b(_arrivedPointer__q)
    );
    wire _node_439;
    BITWISEAND #(.width(1)) bitwiseand_891 (
        .y(_node_439),
        .a(1'h1),
        .b(_node_438)
    );
    wire [7:0] _GEN_230;
    MUX_UNSIGNED #(.width(8)) u_mux_892 (
        .y(_GEN_230),
        .sel(_node_439),
        .a(helloWorld_220),
        .b(_GEN_229)
    );
    wire _node_440;
    wire [8:0] _WTEMP_222;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_893 (
        .y(_WTEMP_222),
        .in(8'hDD)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_894 (
        .y(_node_440),
        .a(_WTEMP_222),
        .b(_arrivedPointer__q)
    );
    wire _node_441;
    BITWISEAND #(.width(1)) bitwiseand_895 (
        .y(_node_441),
        .a(1'h1),
        .b(_node_440)
    );
    wire [7:0] _GEN_231;
    MUX_UNSIGNED #(.width(8)) u_mux_896 (
        .y(_GEN_231),
        .sel(_node_441),
        .a(helloWorld_221),
        .b(_GEN_230)
    );
    wire _node_442;
    wire [8:0] _WTEMP_223;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_897 (
        .y(_WTEMP_223),
        .in(8'hDE)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_898 (
        .y(_node_442),
        .a(_WTEMP_223),
        .b(_arrivedPointer__q)
    );
    wire _node_443;
    BITWISEAND #(.width(1)) bitwiseand_899 (
        .y(_node_443),
        .a(1'h1),
        .b(_node_442)
    );
    wire [7:0] _GEN_232;
    MUX_UNSIGNED #(.width(8)) u_mux_900 (
        .y(_GEN_232),
        .sel(_node_443),
        .a(helloWorld_222),
        .b(_GEN_231)
    );
    wire _node_444;
    wire [8:0] _WTEMP_224;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_901 (
        .y(_WTEMP_224),
        .in(8'hDF)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_902 (
        .y(_node_444),
        .a(_WTEMP_224),
        .b(_arrivedPointer__q)
    );
    wire _node_445;
    BITWISEAND #(.width(1)) bitwiseand_903 (
        .y(_node_445),
        .a(1'h1),
        .b(_node_444)
    );
    wire [7:0] _GEN_233;
    MUX_UNSIGNED #(.width(8)) u_mux_904 (
        .y(_GEN_233),
        .sel(_node_445),
        .a(helloWorld_223),
        .b(_GEN_232)
    );
    wire _node_446;
    wire [8:0] _WTEMP_225;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_905 (
        .y(_WTEMP_225),
        .in(8'hE0)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_906 (
        .y(_node_446),
        .a(_WTEMP_225),
        .b(_arrivedPointer__q)
    );
    wire _node_447;
    BITWISEAND #(.width(1)) bitwiseand_907 (
        .y(_node_447),
        .a(1'h1),
        .b(_node_446)
    );
    wire [7:0] _GEN_234;
    MUX_UNSIGNED #(.width(8)) u_mux_908 (
        .y(_GEN_234),
        .sel(_node_447),
        .a(helloWorld_224),
        .b(_GEN_233)
    );
    wire _node_448;
    wire [8:0] _WTEMP_226;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_909 (
        .y(_WTEMP_226),
        .in(8'hE1)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_910 (
        .y(_node_448),
        .a(_WTEMP_226),
        .b(_arrivedPointer__q)
    );
    wire _node_449;
    BITWISEAND #(.width(1)) bitwiseand_911 (
        .y(_node_449),
        .a(1'h1),
        .b(_node_448)
    );
    wire [7:0] _GEN_235;
    MUX_UNSIGNED #(.width(8)) u_mux_912 (
        .y(_GEN_235),
        .sel(_node_449),
        .a(helloWorld_225),
        .b(_GEN_234)
    );
    wire _node_450;
    wire [8:0] _WTEMP_227;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_913 (
        .y(_WTEMP_227),
        .in(8'hE2)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_914 (
        .y(_node_450),
        .a(_WTEMP_227),
        .b(_arrivedPointer__q)
    );
    wire _node_451;
    BITWISEAND #(.width(1)) bitwiseand_915 (
        .y(_node_451),
        .a(1'h1),
        .b(_node_450)
    );
    wire [7:0] _GEN_236;
    MUX_UNSIGNED #(.width(8)) u_mux_916 (
        .y(_GEN_236),
        .sel(_node_451),
        .a(helloWorld_226),
        .b(_GEN_235)
    );
    wire _node_452;
    wire [8:0] _WTEMP_228;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_917 (
        .y(_WTEMP_228),
        .in(8'hE3)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_918 (
        .y(_node_452),
        .a(_WTEMP_228),
        .b(_arrivedPointer__q)
    );
    wire _node_453;
    BITWISEAND #(.width(1)) bitwiseand_919 (
        .y(_node_453),
        .a(1'h1),
        .b(_node_452)
    );
    wire [7:0] _GEN_237;
    MUX_UNSIGNED #(.width(8)) u_mux_920 (
        .y(_GEN_237),
        .sel(_node_453),
        .a(helloWorld_227),
        .b(_GEN_236)
    );
    wire _node_454;
    wire [8:0] _WTEMP_229;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_921 (
        .y(_WTEMP_229),
        .in(8'hE4)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_922 (
        .y(_node_454),
        .a(_WTEMP_229),
        .b(_arrivedPointer__q)
    );
    wire _node_455;
    BITWISEAND #(.width(1)) bitwiseand_923 (
        .y(_node_455),
        .a(1'h1),
        .b(_node_454)
    );
    wire [7:0] _GEN_238;
    MUX_UNSIGNED #(.width(8)) u_mux_924 (
        .y(_GEN_238),
        .sel(_node_455),
        .a(helloWorld_228),
        .b(_GEN_237)
    );
    wire _node_456;
    wire [8:0] _WTEMP_230;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_925 (
        .y(_WTEMP_230),
        .in(8'hE5)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_926 (
        .y(_node_456),
        .a(_WTEMP_230),
        .b(_arrivedPointer__q)
    );
    wire _node_457;
    BITWISEAND #(.width(1)) bitwiseand_927 (
        .y(_node_457),
        .a(1'h1),
        .b(_node_456)
    );
    wire [7:0] _GEN_239;
    MUX_UNSIGNED #(.width(8)) u_mux_928 (
        .y(_GEN_239),
        .sel(_node_457),
        .a(helloWorld_229),
        .b(_GEN_238)
    );
    wire _node_458;
    wire [8:0] _WTEMP_231;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_929 (
        .y(_WTEMP_231),
        .in(8'hE6)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_930 (
        .y(_node_458),
        .a(_WTEMP_231),
        .b(_arrivedPointer__q)
    );
    wire _node_459;
    BITWISEAND #(.width(1)) bitwiseand_931 (
        .y(_node_459),
        .a(1'h1),
        .b(_node_458)
    );
    wire [7:0] _GEN_240;
    MUX_UNSIGNED #(.width(8)) u_mux_932 (
        .y(_GEN_240),
        .sel(_node_459),
        .a(helloWorld_230),
        .b(_GEN_239)
    );
    wire _node_460;
    wire [8:0] _WTEMP_232;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_933 (
        .y(_WTEMP_232),
        .in(8'hE7)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_934 (
        .y(_node_460),
        .a(_WTEMP_232),
        .b(_arrivedPointer__q)
    );
    wire _node_461;
    BITWISEAND #(.width(1)) bitwiseand_935 (
        .y(_node_461),
        .a(1'h1),
        .b(_node_460)
    );
    wire [7:0] _GEN_241;
    MUX_UNSIGNED #(.width(8)) u_mux_936 (
        .y(_GEN_241),
        .sel(_node_461),
        .a(helloWorld_231),
        .b(_GEN_240)
    );
    wire _node_462;
    wire [8:0] _WTEMP_233;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_937 (
        .y(_WTEMP_233),
        .in(8'hE8)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_938 (
        .y(_node_462),
        .a(_WTEMP_233),
        .b(_arrivedPointer__q)
    );
    wire _node_463;
    BITWISEAND #(.width(1)) bitwiseand_939 (
        .y(_node_463),
        .a(1'h1),
        .b(_node_462)
    );
    wire [7:0] _GEN_242;
    MUX_UNSIGNED #(.width(8)) u_mux_940 (
        .y(_GEN_242),
        .sel(_node_463),
        .a(helloWorld_232),
        .b(_GEN_241)
    );
    wire _node_464;
    wire [8:0] _WTEMP_234;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_941 (
        .y(_WTEMP_234),
        .in(8'hE9)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_942 (
        .y(_node_464),
        .a(_WTEMP_234),
        .b(_arrivedPointer__q)
    );
    wire _node_465;
    BITWISEAND #(.width(1)) bitwiseand_943 (
        .y(_node_465),
        .a(1'h1),
        .b(_node_464)
    );
    wire [7:0] _GEN_243;
    MUX_UNSIGNED #(.width(8)) u_mux_944 (
        .y(_GEN_243),
        .sel(_node_465),
        .a(helloWorld_233),
        .b(_GEN_242)
    );
    wire _node_466;
    wire [8:0] _WTEMP_235;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_945 (
        .y(_WTEMP_235),
        .in(8'hEA)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_946 (
        .y(_node_466),
        .a(_WTEMP_235),
        .b(_arrivedPointer__q)
    );
    wire _node_467;
    BITWISEAND #(.width(1)) bitwiseand_947 (
        .y(_node_467),
        .a(1'h1),
        .b(_node_466)
    );
    wire [7:0] _GEN_244;
    MUX_UNSIGNED #(.width(8)) u_mux_948 (
        .y(_GEN_244),
        .sel(_node_467),
        .a(helloWorld_234),
        .b(_GEN_243)
    );
    wire _node_468;
    wire [8:0] _WTEMP_236;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_949 (
        .y(_WTEMP_236),
        .in(8'hEB)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_950 (
        .y(_node_468),
        .a(_WTEMP_236),
        .b(_arrivedPointer__q)
    );
    wire _node_469;
    BITWISEAND #(.width(1)) bitwiseand_951 (
        .y(_node_469),
        .a(1'h1),
        .b(_node_468)
    );
    wire [7:0] _GEN_245;
    MUX_UNSIGNED #(.width(8)) u_mux_952 (
        .y(_GEN_245),
        .sel(_node_469),
        .a(helloWorld_235),
        .b(_GEN_244)
    );
    wire _node_470;
    wire [8:0] _WTEMP_237;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_953 (
        .y(_WTEMP_237),
        .in(8'hEC)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_954 (
        .y(_node_470),
        .a(_WTEMP_237),
        .b(_arrivedPointer__q)
    );
    wire _node_471;
    BITWISEAND #(.width(1)) bitwiseand_955 (
        .y(_node_471),
        .a(1'h1),
        .b(_node_470)
    );
    wire [7:0] _GEN_246;
    MUX_UNSIGNED #(.width(8)) u_mux_956 (
        .y(_GEN_246),
        .sel(_node_471),
        .a(helloWorld_236),
        .b(_GEN_245)
    );
    wire _node_472;
    wire [8:0] _WTEMP_238;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_957 (
        .y(_WTEMP_238),
        .in(8'hED)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_958 (
        .y(_node_472),
        .a(_WTEMP_238),
        .b(_arrivedPointer__q)
    );
    wire _node_473;
    BITWISEAND #(.width(1)) bitwiseand_959 (
        .y(_node_473),
        .a(1'h1),
        .b(_node_472)
    );
    wire [7:0] _GEN_247;
    MUX_UNSIGNED #(.width(8)) u_mux_960 (
        .y(_GEN_247),
        .sel(_node_473),
        .a(helloWorld_237),
        .b(_GEN_246)
    );
    wire _node_474;
    wire [8:0] _WTEMP_239;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_961 (
        .y(_WTEMP_239),
        .in(8'hEE)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_962 (
        .y(_node_474),
        .a(_WTEMP_239),
        .b(_arrivedPointer__q)
    );
    wire _node_475;
    BITWISEAND #(.width(1)) bitwiseand_963 (
        .y(_node_475),
        .a(1'h1),
        .b(_node_474)
    );
    wire [7:0] _GEN_248;
    MUX_UNSIGNED #(.width(8)) u_mux_964 (
        .y(_GEN_248),
        .sel(_node_475),
        .a(helloWorld_238),
        .b(_GEN_247)
    );
    wire _node_476;
    wire [8:0] _WTEMP_240;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_965 (
        .y(_WTEMP_240),
        .in(8'hEF)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_966 (
        .y(_node_476),
        .a(_WTEMP_240),
        .b(_arrivedPointer__q)
    );
    wire _node_477;
    BITWISEAND #(.width(1)) bitwiseand_967 (
        .y(_node_477),
        .a(1'h1),
        .b(_node_476)
    );
    wire [7:0] _GEN_249;
    MUX_UNSIGNED #(.width(8)) u_mux_968 (
        .y(_GEN_249),
        .sel(_node_477),
        .a(helloWorld_239),
        .b(_GEN_248)
    );
    wire _node_478;
    wire [8:0] _WTEMP_241;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_969 (
        .y(_WTEMP_241),
        .in(8'hF0)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_970 (
        .y(_node_478),
        .a(_WTEMP_241),
        .b(_arrivedPointer__q)
    );
    wire _node_479;
    BITWISEAND #(.width(1)) bitwiseand_971 (
        .y(_node_479),
        .a(1'h1),
        .b(_node_478)
    );
    wire [7:0] _GEN_250;
    MUX_UNSIGNED #(.width(8)) u_mux_972 (
        .y(_GEN_250),
        .sel(_node_479),
        .a(helloWorld_240),
        .b(_GEN_249)
    );
    wire _node_480;
    wire [8:0] _WTEMP_242;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_973 (
        .y(_WTEMP_242),
        .in(8'hF1)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_974 (
        .y(_node_480),
        .a(_WTEMP_242),
        .b(_arrivedPointer__q)
    );
    wire _node_481;
    BITWISEAND #(.width(1)) bitwiseand_975 (
        .y(_node_481),
        .a(1'h1),
        .b(_node_480)
    );
    wire [7:0] _GEN_251;
    MUX_UNSIGNED #(.width(8)) u_mux_976 (
        .y(_GEN_251),
        .sel(_node_481),
        .a(helloWorld_241),
        .b(_GEN_250)
    );
    wire _node_482;
    wire [8:0] _WTEMP_243;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_977 (
        .y(_WTEMP_243),
        .in(8'hF2)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_978 (
        .y(_node_482),
        .a(_WTEMP_243),
        .b(_arrivedPointer__q)
    );
    wire _node_483;
    BITWISEAND #(.width(1)) bitwiseand_979 (
        .y(_node_483),
        .a(1'h1),
        .b(_node_482)
    );
    wire [7:0] _GEN_252;
    MUX_UNSIGNED #(.width(8)) u_mux_980 (
        .y(_GEN_252),
        .sel(_node_483),
        .a(helloWorld_242),
        .b(_GEN_251)
    );
    wire _node_484;
    wire [8:0] _WTEMP_244;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_981 (
        .y(_WTEMP_244),
        .in(8'hF3)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_982 (
        .y(_node_484),
        .a(_WTEMP_244),
        .b(_arrivedPointer__q)
    );
    wire _node_485;
    BITWISEAND #(.width(1)) bitwiseand_983 (
        .y(_node_485),
        .a(1'h1),
        .b(_node_484)
    );
    wire [7:0] _GEN_253;
    MUX_UNSIGNED #(.width(8)) u_mux_984 (
        .y(_GEN_253),
        .sel(_node_485),
        .a(helloWorld_243),
        .b(_GEN_252)
    );
    wire _node_486;
    wire [8:0] _WTEMP_245;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_985 (
        .y(_WTEMP_245),
        .in(8'hF4)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_986 (
        .y(_node_486),
        .a(_WTEMP_245),
        .b(_arrivedPointer__q)
    );
    wire _node_487;
    BITWISEAND #(.width(1)) bitwiseand_987 (
        .y(_node_487),
        .a(1'h1),
        .b(_node_486)
    );
    wire [7:0] _GEN_254;
    MUX_UNSIGNED #(.width(8)) u_mux_988 (
        .y(_GEN_254),
        .sel(_node_487),
        .a(helloWorld_244),
        .b(_GEN_253)
    );
    wire _node_488;
    wire [8:0] _WTEMP_246;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_989 (
        .y(_WTEMP_246),
        .in(8'hF5)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_990 (
        .y(_node_488),
        .a(_WTEMP_246),
        .b(_arrivedPointer__q)
    );
    wire _node_489;
    BITWISEAND #(.width(1)) bitwiseand_991 (
        .y(_node_489),
        .a(1'h1),
        .b(_node_488)
    );
    wire [7:0] _GEN_255;
    MUX_UNSIGNED #(.width(8)) u_mux_992 (
        .y(_GEN_255),
        .sel(_node_489),
        .a(helloWorld_245),
        .b(_GEN_254)
    );
    wire _node_490;
    wire [8:0] _WTEMP_247;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_993 (
        .y(_WTEMP_247),
        .in(8'hF6)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_994 (
        .y(_node_490),
        .a(_WTEMP_247),
        .b(_arrivedPointer__q)
    );
    wire _node_491;
    BITWISEAND #(.width(1)) bitwiseand_995 (
        .y(_node_491),
        .a(1'h1),
        .b(_node_490)
    );
    wire [7:0] _GEN_256;
    MUX_UNSIGNED #(.width(8)) u_mux_996 (
        .y(_GEN_256),
        .sel(_node_491),
        .a(helloWorld_246),
        .b(_GEN_255)
    );
    wire _node_492;
    wire [8:0] _WTEMP_248;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_997 (
        .y(_WTEMP_248),
        .in(8'hF7)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_998 (
        .y(_node_492),
        .a(_WTEMP_248),
        .b(_arrivedPointer__q)
    );
    wire _node_493;
    BITWISEAND #(.width(1)) bitwiseand_999 (
        .y(_node_493),
        .a(1'h1),
        .b(_node_492)
    );
    wire [7:0] _GEN_257;
    MUX_UNSIGNED #(.width(8)) u_mux_1000 (
        .y(_GEN_257),
        .sel(_node_493),
        .a(helloWorld_247),
        .b(_GEN_256)
    );
    wire _node_494;
    wire [8:0] _WTEMP_249;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_1001 (
        .y(_WTEMP_249),
        .in(8'hF8)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_1002 (
        .y(_node_494),
        .a(_WTEMP_249),
        .b(_arrivedPointer__q)
    );
    wire _node_495;
    BITWISEAND #(.width(1)) bitwiseand_1003 (
        .y(_node_495),
        .a(1'h1),
        .b(_node_494)
    );
    wire [7:0] _GEN_258;
    MUX_UNSIGNED #(.width(8)) u_mux_1004 (
        .y(_GEN_258),
        .sel(_node_495),
        .a(helloWorld_248),
        .b(_GEN_257)
    );
    wire _node_496;
    wire [8:0] _WTEMP_250;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_1005 (
        .y(_WTEMP_250),
        .in(8'hF9)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_1006 (
        .y(_node_496),
        .a(_WTEMP_250),
        .b(_arrivedPointer__q)
    );
    wire _node_497;
    BITWISEAND #(.width(1)) bitwiseand_1007 (
        .y(_node_497),
        .a(1'h1),
        .b(_node_496)
    );
    wire [7:0] _GEN_259;
    MUX_UNSIGNED #(.width(8)) u_mux_1008 (
        .y(_GEN_259),
        .sel(_node_497),
        .a(helloWorld_249),
        .b(_GEN_258)
    );
    wire _node_498;
    wire [8:0] _WTEMP_251;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_1009 (
        .y(_WTEMP_251),
        .in(8'hFA)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_1010 (
        .y(_node_498),
        .a(_WTEMP_251),
        .b(_arrivedPointer__q)
    );
    wire _node_499;
    BITWISEAND #(.width(1)) bitwiseand_1011 (
        .y(_node_499),
        .a(1'h1),
        .b(_node_498)
    );
    wire [7:0] _GEN_260;
    MUX_UNSIGNED #(.width(8)) u_mux_1012 (
        .y(_GEN_260),
        .sel(_node_499),
        .a(helloWorld_250),
        .b(_GEN_259)
    );
    wire _node_500;
    wire [8:0] _WTEMP_252;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_1013 (
        .y(_WTEMP_252),
        .in(8'hFB)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_1014 (
        .y(_node_500),
        .a(_WTEMP_252),
        .b(_arrivedPointer__q)
    );
    wire _node_501;
    BITWISEAND #(.width(1)) bitwiseand_1015 (
        .y(_node_501),
        .a(1'h1),
        .b(_node_500)
    );
    wire [7:0] _GEN_261;
    MUX_UNSIGNED #(.width(8)) u_mux_1016 (
        .y(_GEN_261),
        .sel(_node_501),
        .a(helloWorld_251),
        .b(_GEN_260)
    );
    wire _node_502;
    wire [8:0] _WTEMP_253;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_1017 (
        .y(_WTEMP_253),
        .in(8'hFC)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_1018 (
        .y(_node_502),
        .a(_WTEMP_253),
        .b(_arrivedPointer__q)
    );
    wire _node_503;
    BITWISEAND #(.width(1)) bitwiseand_1019 (
        .y(_node_503),
        .a(1'h1),
        .b(_node_502)
    );
    wire [7:0] _GEN_262;
    MUX_UNSIGNED #(.width(8)) u_mux_1020 (
        .y(_GEN_262),
        .sel(_node_503),
        .a(helloWorld_252),
        .b(_GEN_261)
    );
    wire _node_504;
    wire [8:0] _WTEMP_254;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_1021 (
        .y(_WTEMP_254),
        .in(8'hFD)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_1022 (
        .y(_node_504),
        .a(_WTEMP_254),
        .b(_arrivedPointer__q)
    );
    wire _node_505;
    BITWISEAND #(.width(1)) bitwiseand_1023 (
        .y(_node_505),
        .a(1'h1),
        .b(_node_504)
    );
    wire [7:0] _GEN_263;
    MUX_UNSIGNED #(.width(8)) u_mux_1024 (
        .y(_GEN_263),
        .sel(_node_505),
        .a(helloWorld_253),
        .b(_GEN_262)
    );
    wire _node_506;
    wire [8:0] _WTEMP_255;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_1025 (
        .y(_WTEMP_255),
        .in(8'hFE)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_1026 (
        .y(_node_506),
        .a(_WTEMP_255),
        .b(_arrivedPointer__q)
    );
    wire _node_507;
    BITWISEAND #(.width(1)) bitwiseand_1027 (
        .y(_node_507),
        .a(1'h1),
        .b(_node_506)
    );
    wire [7:0] _GEN_264;
    MUX_UNSIGNED #(.width(8)) u_mux_1028 (
        .y(_GEN_264),
        .sel(_node_507),
        .a(helloWorld_254),
        .b(_GEN_263)
    );
    wire _node_508;
    wire [8:0] _WTEMP_256;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_1029 (
        .y(_WTEMP_256),
        .in(8'hFF)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_1030 (
        .y(_node_508),
        .a(_WTEMP_256),
        .b(_arrivedPointer__q)
    );
    wire _node_509;
    BITWISEAND #(.width(1)) bitwiseand_1031 (
        .y(_node_509),
        .a(1'h1),
        .b(_node_508)
    );
    wire [7:0] _GEN_265;
    MUX_UNSIGNED #(.width(8)) u_mux_1032 (
        .y(_GEN_265),
        .sel(_node_509),
        .a(helloWorld_255),
        .b(_GEN_264)
    );
    wire _node_510;
    EQ_UNSIGNED #(.width(9)) u_eq_1033 (
        .y(_node_510),
        .a(9'h100),
        .b(_arrivedPointer__q)
    );
    wire _node_511;
    BITWISEAND #(.width(1)) bitwiseand_1034 (
        .y(_node_511),
        .a(1'h1),
        .b(_node_510)
    );
    wire [7:0] _GEN_266;
    MUX_UNSIGNED #(.width(8)) u_mux_1035 (
        .y(_GEN_266),
        .sel(_node_511),
        .a(helloWorld_256),
        .b(_GEN_265)
    );
    wire _node_512;
    EQ_UNSIGNED #(.width(9)) u_eq_1036 (
        .y(_node_512),
        .a(9'h101),
        .b(_arrivedPointer__q)
    );
    wire _node_513;
    BITWISEAND #(.width(1)) bitwiseand_1037 (
        .y(_node_513),
        .a(1'h1),
        .b(_node_512)
    );
    wire [7:0] _GEN_267;
    MUX_UNSIGNED #(.width(8)) u_mux_1038 (
        .y(_GEN_267),
        .sel(_node_513),
        .a(helloWorld_257),
        .b(_GEN_266)
    );
    wire _node_514;
    EQ_UNSIGNED #(.width(9)) u_eq_1039 (
        .y(_node_514),
        .a(9'h102),
        .b(_arrivedPointer__q)
    );
    wire _node_515;
    BITWISEAND #(.width(1)) bitwiseand_1040 (
        .y(_node_515),
        .a(1'h1),
        .b(_node_514)
    );
    wire [7:0] _GEN_268;
    MUX_UNSIGNED #(.width(8)) u_mux_1041 (
        .y(_GEN_268),
        .sel(_node_515),
        .a(helloWorld_258),
        .b(_GEN_267)
    );
    wire _node_516;
    EQ_UNSIGNED #(.width(9)) u_eq_1042 (
        .y(_node_516),
        .a(9'h103),
        .b(_arrivedPointer__q)
    );
    wire _node_517;
    BITWISEAND #(.width(1)) bitwiseand_1043 (
        .y(_node_517),
        .a(1'h1),
        .b(_node_516)
    );
    wire [7:0] _GEN_269;
    MUX_UNSIGNED #(.width(8)) u_mux_1044 (
        .y(_GEN_269),
        .sel(_node_517),
        .a(helloWorld_259),
        .b(_GEN_268)
    );
    wire _node_518;
    EQ_UNSIGNED #(.width(9)) u_eq_1045 (
        .y(_node_518),
        .a(9'h104),
        .b(_arrivedPointer__q)
    );
    wire _node_519;
    BITWISEAND #(.width(1)) bitwiseand_1046 (
        .y(_node_519),
        .a(1'h1),
        .b(_node_518)
    );
    wire [7:0] _GEN_270;
    MUX_UNSIGNED #(.width(8)) u_mux_1047 (
        .y(_GEN_270),
        .sel(_node_519),
        .a(helloWorld_260),
        .b(_GEN_269)
    );
    wire _node_520;
    EQ_UNSIGNED #(.width(9)) u_eq_1048 (
        .y(_node_520),
        .a(9'h105),
        .b(_arrivedPointer__q)
    );
    wire _node_521;
    BITWISEAND #(.width(1)) bitwiseand_1049 (
        .y(_node_521),
        .a(1'h1),
        .b(_node_520)
    );
    wire [7:0] _GEN_271;
    MUX_UNSIGNED #(.width(8)) u_mux_1050 (
        .y(_GEN_271),
        .sel(_node_521),
        .a(helloWorld_261),
        .b(_GEN_270)
    );
    wire _node_522;
    EQ_UNSIGNED #(.width(9)) u_eq_1051 (
        .y(_node_522),
        .a(9'h106),
        .b(_arrivedPointer__q)
    );
    wire _node_523;
    BITWISEAND #(.width(1)) bitwiseand_1052 (
        .y(_node_523),
        .a(1'h1),
        .b(_node_522)
    );
    wire [7:0] _GEN_272;
    MUX_UNSIGNED #(.width(8)) u_mux_1053 (
        .y(_GEN_272),
        .sel(_node_523),
        .a(helloWorld_262),
        .b(_GEN_271)
    );
    wire _node_524;
    EQ_UNSIGNED #(.width(9)) u_eq_1054 (
        .y(_node_524),
        .a(9'h107),
        .b(_arrivedPointer__q)
    );
    wire _node_525;
    BITWISEAND #(.width(1)) bitwiseand_1055 (
        .y(_node_525),
        .a(1'h1),
        .b(_node_524)
    );
    wire [7:0] _GEN_273;
    MUX_UNSIGNED #(.width(8)) u_mux_1056 (
        .y(_GEN_273),
        .sel(_node_525),
        .a(helloWorld_263),
        .b(_GEN_272)
    );
    wire _node_526;
    EQ_UNSIGNED #(.width(9)) u_eq_1057 (
        .y(_node_526),
        .a(9'h108),
        .b(_arrivedPointer__q)
    );
    wire _node_527;
    BITWISEAND #(.width(1)) bitwiseand_1058 (
        .y(_node_527),
        .a(1'h1),
        .b(_node_526)
    );
    wire [7:0] _GEN_274;
    MUX_UNSIGNED #(.width(8)) u_mux_1059 (
        .y(_GEN_274),
        .sel(_node_527),
        .a(helloWorld_264),
        .b(_GEN_273)
    );
    wire _node_528;
    EQ_UNSIGNED #(.width(9)) u_eq_1060 (
        .y(_node_528),
        .a(9'h109),
        .b(_arrivedPointer__q)
    );
    wire _node_529;
    BITWISEAND #(.width(1)) bitwiseand_1061 (
        .y(_node_529),
        .a(1'h1),
        .b(_node_528)
    );
    wire [7:0] _GEN_275;
    MUX_UNSIGNED #(.width(8)) u_mux_1062 (
        .y(_GEN_275),
        .sel(_node_529),
        .a(helloWorld_265),
        .b(_GEN_274)
    );
    wire _node_530;
    EQ_UNSIGNED #(.width(9)) u_eq_1063 (
        .y(_node_530),
        .a(9'h10A),
        .b(_arrivedPointer__q)
    );
    wire _node_531;
    BITWISEAND #(.width(1)) bitwiseand_1064 (
        .y(_node_531),
        .a(1'h1),
        .b(_node_530)
    );
    wire [7:0] _GEN_276;
    MUX_UNSIGNED #(.width(8)) u_mux_1065 (
        .y(_GEN_276),
        .sel(_node_531),
        .a(helloWorld_266),
        .b(_GEN_275)
    );
    wire _node_532;
    EQ_UNSIGNED #(.width(9)) u_eq_1066 (
        .y(_node_532),
        .a(9'h10B),
        .b(_arrivedPointer__q)
    );
    wire _node_533;
    BITWISEAND #(.width(1)) bitwiseand_1067 (
        .y(_node_533),
        .a(1'h1),
        .b(_node_532)
    );
    wire [7:0] _GEN_277;
    MUX_UNSIGNED #(.width(8)) u_mux_1068 (
        .y(_GEN_277),
        .sel(_node_533),
        .a(helloWorld_267),
        .b(_GEN_276)
    );
    wire _node_534;
    EQ_UNSIGNED #(.width(9)) u_eq_1069 (
        .y(_node_534),
        .a(9'h10C),
        .b(_arrivedPointer__q)
    );
    wire _node_535;
    BITWISEAND #(.width(1)) bitwiseand_1070 (
        .y(_node_535),
        .a(1'h1),
        .b(_node_534)
    );
    wire [7:0] _GEN_278;
    MUX_UNSIGNED #(.width(8)) u_mux_1071 (
        .y(_GEN_278),
        .sel(_node_535),
        .a(helloWorld_268),
        .b(_GEN_277)
    );
    wire _node_536;
    EQ_UNSIGNED #(.width(9)) u_eq_1072 (
        .y(_node_536),
        .a(9'h10D),
        .b(_arrivedPointer__q)
    );
    wire _node_537;
    BITWISEAND #(.width(1)) bitwiseand_1073 (
        .y(_node_537),
        .a(1'h1),
        .b(_node_536)
    );
    wire [7:0] _GEN_279;
    MUX_UNSIGNED #(.width(8)) u_mux_1074 (
        .y(_GEN_279),
        .sel(_node_537),
        .a(helloWorld_269),
        .b(_GEN_278)
    );
    wire _node_538;
    EQ_UNSIGNED #(.width(9)) u_eq_1075 (
        .y(_node_538),
        .a(9'h10E),
        .b(_arrivedPointer__q)
    );
    wire _node_539;
    BITWISEAND #(.width(1)) bitwiseand_1076 (
        .y(_node_539),
        .a(1'h1),
        .b(_node_538)
    );
    wire [7:0] _GEN_280;
    MUX_UNSIGNED #(.width(8)) u_mux_1077 (
        .y(_GEN_280),
        .sel(_node_539),
        .a(helloWorld_270),
        .b(_GEN_279)
    );
    wire _node_540;
    EQ_UNSIGNED #(.width(9)) u_eq_1078 (
        .y(_node_540),
        .a(9'h10F),
        .b(_arrivedPointer__q)
    );
    wire _node_541;
    BITWISEAND #(.width(1)) bitwiseand_1079 (
        .y(_node_541),
        .a(1'h1),
        .b(_node_540)
    );
    wire [7:0] _GEN_281;
    MUX_UNSIGNED #(.width(8)) u_mux_1080 (
        .y(_GEN_281),
        .sel(_node_541),
        .a(helloWorld_271),
        .b(_GEN_280)
    );
    wire _node_542;
    EQ_UNSIGNED #(.width(9)) u_eq_1081 (
        .y(_node_542),
        .a(9'h110),
        .b(_arrivedPointer__q)
    );
    wire _node_543;
    BITWISEAND #(.width(1)) bitwiseand_1082 (
        .y(_node_543),
        .a(1'h1),
        .b(_node_542)
    );
    wire [7:0] _GEN_282;
    MUX_UNSIGNED #(.width(8)) u_mux_1083 (
        .y(_GEN_282),
        .sel(_node_543),
        .a(helloWorld_272),
        .b(_GEN_281)
    );
    wire _node_544;
    EQ_UNSIGNED #(.width(9)) u_eq_1084 (
        .y(_node_544),
        .a(9'h111),
        .b(_arrivedPointer__q)
    );
    wire _node_545;
    BITWISEAND #(.width(1)) bitwiseand_1085 (
        .y(_node_545),
        .a(1'h1),
        .b(_node_544)
    );
    wire [7:0] _GEN_283;
    MUX_UNSIGNED #(.width(8)) u_mux_1086 (
        .y(_GEN_283),
        .sel(_node_545),
        .a(helloWorld_273),
        .b(_GEN_282)
    );
    wire _node_546;
    EQ_UNSIGNED #(.width(9)) u_eq_1087 (
        .y(_node_546),
        .a(9'h112),
        .b(_arrivedPointer__q)
    );
    wire _node_547;
    BITWISEAND #(.width(1)) bitwiseand_1088 (
        .y(_node_547),
        .a(1'h1),
        .b(_node_546)
    );
    wire [7:0] _GEN_284;
    MUX_UNSIGNED #(.width(8)) u_mux_1089 (
        .y(_GEN_284),
        .sel(_node_547),
        .a(helloWorld_274),
        .b(_GEN_283)
    );
    wire _node_548;
    EQ_UNSIGNED #(.width(9)) u_eq_1090 (
        .y(_node_548),
        .a(9'h113),
        .b(_arrivedPointer__q)
    );
    wire _node_549;
    BITWISEAND #(.width(1)) bitwiseand_1091 (
        .y(_node_549),
        .a(1'h1),
        .b(_node_548)
    );
    wire [7:0] _GEN_285;
    MUX_UNSIGNED #(.width(8)) u_mux_1092 (
        .y(_GEN_285),
        .sel(_node_549),
        .a(helloWorld_275),
        .b(_GEN_284)
    );
    wire _node_550;
    EQ_UNSIGNED #(.width(9)) u_eq_1093 (
        .y(_node_550),
        .a(9'h114),
        .b(_arrivedPointer__q)
    );
    wire _node_551;
    BITWISEAND #(.width(1)) bitwiseand_1094 (
        .y(_node_551),
        .a(1'h1),
        .b(_node_550)
    );
    wire [7:0] _GEN_286;
    MUX_UNSIGNED #(.width(8)) u_mux_1095 (
        .y(_GEN_286),
        .sel(_node_551),
        .a(helloWorld_276),
        .b(_GEN_285)
    );
    wire _node_552;
    EQ_UNSIGNED #(.width(9)) u_eq_1096 (
        .y(_node_552),
        .a(9'h115),
        .b(_arrivedPointer__q)
    );
    wire _node_553;
    BITWISEAND #(.width(1)) bitwiseand_1097 (
        .y(_node_553),
        .a(1'h1),
        .b(_node_552)
    );
    wire [7:0] _GEN_287;
    MUX_UNSIGNED #(.width(8)) u_mux_1098 (
        .y(_GEN_287),
        .sel(_node_553),
        .a(helloWorld_277),
        .b(_GEN_286)
    );
    wire _node_554;
    EQ_UNSIGNED #(.width(9)) u_eq_1099 (
        .y(_node_554),
        .a(9'h116),
        .b(_arrivedPointer__q)
    );
    wire _node_555;
    BITWISEAND #(.width(1)) bitwiseand_1100 (
        .y(_node_555),
        .a(1'h1),
        .b(_node_554)
    );
    wire [7:0] _GEN_288;
    MUX_UNSIGNED #(.width(8)) u_mux_1101 (
        .y(_GEN_288),
        .sel(_node_555),
        .a(helloWorld_278),
        .b(_GEN_287)
    );
    wire _node_556;
    EQ_UNSIGNED #(.width(9)) u_eq_1102 (
        .y(_node_556),
        .a(9'h117),
        .b(_arrivedPointer__q)
    );
    wire _node_557;
    BITWISEAND #(.width(1)) bitwiseand_1103 (
        .y(_node_557),
        .a(1'h1),
        .b(_node_556)
    );
    wire [7:0] _GEN_289;
    MUX_UNSIGNED #(.width(8)) u_mux_1104 (
        .y(_GEN_289),
        .sel(_node_557),
        .a(helloWorld_279),
        .b(_GEN_288)
    );
    wire _node_558;
    EQ_UNSIGNED #(.width(9)) u_eq_1105 (
        .y(_node_558),
        .a(9'h118),
        .b(_arrivedPointer__q)
    );
    wire _node_559;
    BITWISEAND #(.width(1)) bitwiseand_1106 (
        .y(_node_559),
        .a(1'h1),
        .b(_node_558)
    );
    wire [7:0] _GEN_290;
    MUX_UNSIGNED #(.width(8)) u_mux_1107 (
        .y(_GEN_290),
        .sel(_node_559),
        .a(helloWorld_280),
        .b(_GEN_289)
    );
    wire _node_560;
    EQ_UNSIGNED #(.width(9)) u_eq_1108 (
        .y(_node_560),
        .a(9'h119),
        .b(_arrivedPointer__q)
    );
    wire _node_561;
    BITWISEAND #(.width(1)) bitwiseand_1109 (
        .y(_node_561),
        .a(1'h1),
        .b(_node_560)
    );
    wire [7:0] _GEN_291;
    MUX_UNSIGNED #(.width(8)) u_mux_1110 (
        .y(_GEN_291),
        .sel(_node_561),
        .a(helloWorld_281),
        .b(_GEN_290)
    );
    wire _node_562;
    EQ_UNSIGNED #(.width(9)) u_eq_1111 (
        .y(_node_562),
        .a(9'h11A),
        .b(_arrivedPointer__q)
    );
    wire _node_563;
    BITWISEAND #(.width(1)) bitwiseand_1112 (
        .y(_node_563),
        .a(1'h1),
        .b(_node_562)
    );
    wire [7:0] _GEN_292;
    MUX_UNSIGNED #(.width(8)) u_mux_1113 (
        .y(_GEN_292),
        .sel(_node_563),
        .a(helloWorld_282),
        .b(_GEN_291)
    );
    wire _node_564;
    EQ_UNSIGNED #(.width(9)) u_eq_1114 (
        .y(_node_564),
        .a(9'h11B),
        .b(_arrivedPointer__q)
    );
    wire _node_565;
    BITWISEAND #(.width(1)) bitwiseand_1115 (
        .y(_node_565),
        .a(1'h1),
        .b(_node_564)
    );
    wire [7:0] _GEN_293;
    MUX_UNSIGNED #(.width(8)) u_mux_1116 (
        .y(_GEN_293),
        .sel(_node_565),
        .a(helloWorld_283),
        .b(_GEN_292)
    );
    wire _node_566;
    EQ_UNSIGNED #(.width(9)) u_eq_1117 (
        .y(_node_566),
        .a(9'h11C),
        .b(_arrivedPointer__q)
    );
    wire _node_567;
    BITWISEAND #(.width(1)) bitwiseand_1118 (
        .y(_node_567),
        .a(1'h1),
        .b(_node_566)
    );
    wire [7:0] _GEN_294;
    MUX_UNSIGNED #(.width(8)) u_mux_1119 (
        .y(_GEN_294),
        .sel(_node_567),
        .a(helloWorld_284),
        .b(_GEN_293)
    );
    wire _node_568;
    EQ_UNSIGNED #(.width(9)) u_eq_1120 (
        .y(_node_568),
        .a(9'h11D),
        .b(_arrivedPointer__q)
    );
    wire _node_569;
    BITWISEAND #(.width(1)) bitwiseand_1121 (
        .y(_node_569),
        .a(1'h1),
        .b(_node_568)
    );
    wire [7:0] _GEN_295;
    MUX_UNSIGNED #(.width(8)) u_mux_1122 (
        .y(_GEN_295),
        .sel(_node_569),
        .a(helloWorld_285),
        .b(_GEN_294)
    );
    wire _node_570;
    EQ_UNSIGNED #(.width(9)) u_eq_1123 (
        .y(_node_570),
        .a(9'h11E),
        .b(_arrivedPointer__q)
    );
    wire _node_571;
    BITWISEAND #(.width(1)) bitwiseand_1124 (
        .y(_node_571),
        .a(1'h1),
        .b(_node_570)
    );
    wire [7:0] _GEN_296;
    MUX_UNSIGNED #(.width(8)) u_mux_1125 (
        .y(_GEN_296),
        .sel(_node_571),
        .a(helloWorld_286),
        .b(_GEN_295)
    );
    wire _node_572;
    EQ_UNSIGNED #(.width(9)) u_eq_1126 (
        .y(_node_572),
        .a(9'h11F),
        .b(_arrivedPointer__q)
    );
    wire _node_573;
    BITWISEAND #(.width(1)) bitwiseand_1127 (
        .y(_node_573),
        .a(1'h1),
        .b(_node_572)
    );
    wire [7:0] _GEN_297;
    MUX_UNSIGNED #(.width(8)) u_mux_1128 (
        .y(_GEN_297),
        .sel(_node_573),
        .a(helloWorld_287),
        .b(_GEN_296)
    );
    wire _node_574;
    EQ_UNSIGNED #(.width(9)) u_eq_1129 (
        .y(_node_574),
        .a(9'h120),
        .b(_arrivedPointer__q)
    );
    wire _node_575;
    BITWISEAND #(.width(1)) bitwiseand_1130 (
        .y(_node_575),
        .a(1'h1),
        .b(_node_574)
    );
    wire [7:0] _GEN_298;
    MUX_UNSIGNED #(.width(8)) u_mux_1131 (
        .y(_GEN_298),
        .sel(_node_575),
        .a(helloWorld_288),
        .b(_GEN_297)
    );
    wire _node_576;
    EQ_UNSIGNED #(.width(9)) u_eq_1132 (
        .y(_node_576),
        .a(9'h121),
        .b(_arrivedPointer__q)
    );
    wire _node_577;
    BITWISEAND #(.width(1)) bitwiseand_1133 (
        .y(_node_577),
        .a(1'h1),
        .b(_node_576)
    );
    wire [7:0] _GEN_299;
    MUX_UNSIGNED #(.width(8)) u_mux_1134 (
        .y(_GEN_299),
        .sel(_node_577),
        .a(helloWorld_289),
        .b(_GEN_298)
    );
    wire _node_578;
    EQ_UNSIGNED #(.width(9)) u_eq_1135 (
        .y(_node_578),
        .a(9'h122),
        .b(_arrivedPointer__q)
    );
    wire _node_579;
    BITWISEAND #(.width(1)) bitwiseand_1136 (
        .y(_node_579),
        .a(1'h1),
        .b(_node_578)
    );
    wire [7:0] _GEN_300;
    MUX_UNSIGNED #(.width(8)) u_mux_1137 (
        .y(_GEN_300),
        .sel(_node_579),
        .a(helloWorld_290),
        .b(_GEN_299)
    );
    wire _node_580;
    EQ_UNSIGNED #(.width(9)) u_eq_1138 (
        .y(_node_580),
        .a(9'h123),
        .b(_arrivedPointer__q)
    );
    wire _node_581;
    BITWISEAND #(.width(1)) bitwiseand_1139 (
        .y(_node_581),
        .a(1'h1),
        .b(_node_580)
    );
    wire [7:0] _GEN_301;
    MUX_UNSIGNED #(.width(8)) u_mux_1140 (
        .y(_GEN_301),
        .sel(_node_581),
        .a(helloWorld_291),
        .b(_GEN_300)
    );
    wire _node_582;
    EQ_UNSIGNED #(.width(9)) u_eq_1141 (
        .y(_node_582),
        .a(9'h124),
        .b(_arrivedPointer__q)
    );
    wire _node_583;
    BITWISEAND #(.width(1)) bitwiseand_1142 (
        .y(_node_583),
        .a(1'h1),
        .b(_node_582)
    );
    wire [7:0] _GEN_302;
    MUX_UNSIGNED #(.width(8)) u_mux_1143 (
        .y(_GEN_302),
        .sel(_node_583),
        .a(helloWorld_292),
        .b(_GEN_301)
    );
    wire _node_584;
    EQ_UNSIGNED #(.width(9)) u_eq_1144 (
        .y(_node_584),
        .a(9'h125),
        .b(_arrivedPointer__q)
    );
    wire _node_585;
    BITWISEAND #(.width(1)) bitwiseand_1145 (
        .y(_node_585),
        .a(1'h1),
        .b(_node_584)
    );
    wire [7:0] _GEN_303;
    MUX_UNSIGNED #(.width(8)) u_mux_1146 (
        .y(_GEN_303),
        .sel(_node_585),
        .a(helloWorld_293),
        .b(_GEN_302)
    );
    wire _node_586;
    EQ_UNSIGNED #(.width(9)) u_eq_1147 (
        .y(_node_586),
        .a(9'h126),
        .b(_arrivedPointer__q)
    );
    wire _node_587;
    BITWISEAND #(.width(1)) bitwiseand_1148 (
        .y(_node_587),
        .a(1'h1),
        .b(_node_586)
    );
    wire [7:0] _GEN_304;
    MUX_UNSIGNED #(.width(8)) u_mux_1149 (
        .y(_GEN_304),
        .sel(_node_587),
        .a(helloWorld_294),
        .b(_GEN_303)
    );
    wire _node_588;
    EQ_UNSIGNED #(.width(9)) u_eq_1150 (
        .y(_node_588),
        .a(9'h127),
        .b(_arrivedPointer__q)
    );
    wire _node_589;
    BITWISEAND #(.width(1)) bitwiseand_1151 (
        .y(_node_589),
        .a(1'h1),
        .b(_node_588)
    );
    wire [7:0] _GEN_305;
    MUX_UNSIGNED #(.width(8)) u_mux_1152 (
        .y(_GEN_305),
        .sel(_node_589),
        .a(helloWorld_295),
        .b(_GEN_304)
    );
    wire _node_590;
    EQ_UNSIGNED #(.width(9)) u_eq_1153 (
        .y(_node_590),
        .a(9'h128),
        .b(_arrivedPointer__q)
    );
    wire _node_591;
    BITWISEAND #(.width(1)) bitwiseand_1154 (
        .y(_node_591),
        .a(1'h1),
        .b(_node_590)
    );
    wire [7:0] _GEN_306;
    MUX_UNSIGNED #(.width(8)) u_mux_1155 (
        .y(_GEN_306),
        .sel(_node_591),
        .a(helloWorld_296),
        .b(_GEN_305)
    );
    wire _node_592;
    EQ_UNSIGNED #(.width(9)) u_eq_1156 (
        .y(_node_592),
        .a(9'h129),
        .b(_arrivedPointer__q)
    );
    wire _node_593;
    BITWISEAND #(.width(1)) bitwiseand_1157 (
        .y(_node_593),
        .a(1'h1),
        .b(_node_592)
    );
    wire [7:0] _GEN_307;
    MUX_UNSIGNED #(.width(8)) u_mux_1158 (
        .y(_GEN_307),
        .sel(_node_593),
        .a(helloWorld_297),
        .b(_GEN_306)
    );
    wire _node_594;
    EQ_UNSIGNED #(.width(9)) u_eq_1159 (
        .y(_node_594),
        .a(9'h12A),
        .b(_arrivedPointer__q)
    );
    wire _node_595;
    BITWISEAND #(.width(1)) bitwiseand_1160 (
        .y(_node_595),
        .a(1'h1),
        .b(_node_594)
    );
    wire [7:0] _GEN_308;
    MUX_UNSIGNED #(.width(8)) u_mux_1161 (
        .y(_GEN_308),
        .sel(_node_595),
        .a(helloWorld_298),
        .b(_GEN_307)
    );
    wire _node_596;
    EQ_UNSIGNED #(.width(9)) u_eq_1162 (
        .y(_node_596),
        .a(9'h12B),
        .b(_arrivedPointer__q)
    );
    wire _node_597;
    BITWISEAND #(.width(1)) bitwiseand_1163 (
        .y(_node_597),
        .a(1'h1),
        .b(_node_596)
    );
    wire [7:0] _GEN_309;
    MUX_UNSIGNED #(.width(8)) u_mux_1164 (
        .y(_GEN_309),
        .sel(_node_597),
        .a(helloWorld_299),
        .b(_GEN_308)
    );
    wire _node_598;
    EQ_UNSIGNED #(.width(9)) u_eq_1165 (
        .y(_node_598),
        .a(9'h12C),
        .b(_arrivedPointer__q)
    );
    wire _node_599;
    BITWISEAND #(.width(1)) bitwiseand_1166 (
        .y(_node_599),
        .a(1'h1),
        .b(_node_598)
    );
    wire [7:0] _GEN_310;
    MUX_UNSIGNED #(.width(8)) u_mux_1167 (
        .y(_GEN_310),
        .sel(_node_599),
        .a(helloWorld_300),
        .b(_GEN_309)
    );
    wire _node_600;
    EQ_UNSIGNED #(.width(9)) u_eq_1168 (
        .y(_node_600),
        .a(9'h12D),
        .b(_arrivedPointer__q)
    );
    wire _node_601;
    BITWISEAND #(.width(1)) bitwiseand_1169 (
        .y(_node_601),
        .a(1'h1),
        .b(_node_600)
    );
    wire [7:0] _GEN_311;
    MUX_UNSIGNED #(.width(8)) u_mux_1170 (
        .y(_GEN_311),
        .sel(_node_601),
        .a(helloWorld_301),
        .b(_GEN_310)
    );
    wire _node_602;
    EQ_UNSIGNED #(.width(9)) u_eq_1171 (
        .y(_node_602),
        .a(9'h12E),
        .b(_arrivedPointer__q)
    );
    wire _node_603;
    BITWISEAND #(.width(1)) bitwiseand_1172 (
        .y(_node_603),
        .a(1'h1),
        .b(_node_602)
    );
    wire [7:0] _GEN_312;
    MUX_UNSIGNED #(.width(8)) u_mux_1173 (
        .y(_GEN_312),
        .sel(_node_603),
        .a(helloWorld_302),
        .b(_GEN_311)
    );
    wire _node_604;
    EQ_UNSIGNED #(.width(9)) u_eq_1174 (
        .y(_node_604),
        .a(9'h12F),
        .b(_arrivedPointer__q)
    );
    wire _node_605;
    BITWISEAND #(.width(1)) bitwiseand_1175 (
        .y(_node_605),
        .a(1'h1),
        .b(_node_604)
    );
    wire [7:0] _GEN_313;
    MUX_UNSIGNED #(.width(8)) u_mux_1176 (
        .y(_GEN_313),
        .sel(_node_605),
        .a(helloWorld_303),
        .b(_GEN_312)
    );
    wire _node_606;
    EQ_UNSIGNED #(.width(9)) u_eq_1177 (
        .y(_node_606),
        .a(9'h130),
        .b(_arrivedPointer__q)
    );
    wire _node_607;
    BITWISEAND #(.width(1)) bitwiseand_1178 (
        .y(_node_607),
        .a(1'h1),
        .b(_node_606)
    );
    wire [7:0] _GEN_314;
    MUX_UNSIGNED #(.width(8)) u_mux_1179 (
        .y(_GEN_314),
        .sel(_node_607),
        .a(helloWorld_304),
        .b(_GEN_313)
    );
    wire _node_608;
    EQ_UNSIGNED #(.width(9)) u_eq_1180 (
        .y(_node_608),
        .a(9'h131),
        .b(_arrivedPointer__q)
    );
    wire _node_609;
    BITWISEAND #(.width(1)) bitwiseand_1181 (
        .y(_node_609),
        .a(1'h1),
        .b(_node_608)
    );
    wire [7:0] _GEN_315;
    MUX_UNSIGNED #(.width(8)) u_mux_1182 (
        .y(_GEN_315),
        .sel(_node_609),
        .a(helloWorld_305),
        .b(_GEN_314)
    );
    wire _node_610;
    EQ_UNSIGNED #(.width(9)) u_eq_1183 (
        .y(_node_610),
        .a(9'h132),
        .b(_arrivedPointer__q)
    );
    wire _node_611;
    BITWISEAND #(.width(1)) bitwiseand_1184 (
        .y(_node_611),
        .a(1'h1),
        .b(_node_610)
    );
    wire [7:0] _GEN_316;
    MUX_UNSIGNED #(.width(8)) u_mux_1185 (
        .y(_GEN_316),
        .sel(_node_611),
        .a(helloWorld_306),
        .b(_GEN_315)
    );
    wire _node_612;
    EQ_UNSIGNED #(.width(9)) u_eq_1186 (
        .y(_node_612),
        .a(9'h133),
        .b(_arrivedPointer__q)
    );
    wire _node_613;
    BITWISEAND #(.width(1)) bitwiseand_1187 (
        .y(_node_613),
        .a(1'h1),
        .b(_node_612)
    );
    wire [7:0] _GEN_317;
    MUX_UNSIGNED #(.width(8)) u_mux_1188 (
        .y(_GEN_317),
        .sel(_node_613),
        .a(helloWorld_307),
        .b(_GEN_316)
    );
    wire _node_614;
    EQ_UNSIGNED #(.width(9)) u_eq_1189 (
        .y(_node_614),
        .a(9'h134),
        .b(_arrivedPointer__q)
    );
    wire _node_615;
    BITWISEAND #(.width(1)) bitwiseand_1190 (
        .y(_node_615),
        .a(1'h1),
        .b(_node_614)
    );
    wire [7:0] _GEN_318;
    MUX_UNSIGNED #(.width(8)) u_mux_1191 (
        .y(_GEN_318),
        .sel(_node_615),
        .a(helloWorld_308),
        .b(_GEN_317)
    );
    wire _node_616;
    EQ_UNSIGNED #(.width(9)) u_eq_1192 (
        .y(_node_616),
        .a(9'h135),
        .b(_arrivedPointer__q)
    );
    wire _node_617;
    BITWISEAND #(.width(1)) bitwiseand_1193 (
        .y(_node_617),
        .a(1'h1),
        .b(_node_616)
    );
    wire [7:0] _GEN_319;
    MUX_UNSIGNED #(.width(8)) u_mux_1194 (
        .y(_GEN_319),
        .sel(_node_617),
        .a(helloWorld_309),
        .b(_GEN_318)
    );
    wire _node_618;
    EQ_UNSIGNED #(.width(9)) u_eq_1195 (
        .y(_node_618),
        .a(9'h136),
        .b(_arrivedPointer__q)
    );
    wire _node_619;
    BITWISEAND #(.width(1)) bitwiseand_1196 (
        .y(_node_619),
        .a(1'h1),
        .b(_node_618)
    );
    wire [7:0] _GEN_320;
    MUX_UNSIGNED #(.width(8)) u_mux_1197 (
        .y(_GEN_320),
        .sel(_node_619),
        .a(helloWorld_310),
        .b(_GEN_319)
    );
    wire _node_620;
    EQ_UNSIGNED #(.width(9)) u_eq_1198 (
        .y(_node_620),
        .a(9'h137),
        .b(_arrivedPointer__q)
    );
    wire _node_621;
    BITWISEAND #(.width(1)) bitwiseand_1199 (
        .y(_node_621),
        .a(1'h1),
        .b(_node_620)
    );
    wire [7:0] _GEN_321;
    MUX_UNSIGNED #(.width(8)) u_mux_1200 (
        .y(_GEN_321),
        .sel(_node_621),
        .a(helloWorld_311),
        .b(_GEN_320)
    );
    wire _node_622;
    EQ_UNSIGNED #(.width(9)) u_eq_1201 (
        .y(_node_622),
        .a(9'h138),
        .b(_arrivedPointer__q)
    );
    wire _node_623;
    BITWISEAND #(.width(1)) bitwiseand_1202 (
        .y(_node_623),
        .a(1'h1),
        .b(_node_622)
    );
    wire [7:0] _GEN_322;
    MUX_UNSIGNED #(.width(8)) u_mux_1203 (
        .y(_GEN_322),
        .sel(_node_623),
        .a(helloWorld_312),
        .b(_GEN_321)
    );
    wire _node_624;
    EQ_UNSIGNED #(.width(9)) u_eq_1204 (
        .y(_node_624),
        .a(9'h139),
        .b(_arrivedPointer__q)
    );
    wire _node_625;
    BITWISEAND #(.width(1)) bitwiseand_1205 (
        .y(_node_625),
        .a(1'h1),
        .b(_node_624)
    );
    wire [7:0] _GEN_323;
    MUX_UNSIGNED #(.width(8)) u_mux_1206 (
        .y(_GEN_323),
        .sel(_node_625),
        .a(helloWorld_313),
        .b(_GEN_322)
    );
    wire _node_626;
    EQ_UNSIGNED #(.width(9)) u_eq_1207 (
        .y(_node_626),
        .a(9'h13A),
        .b(_arrivedPointer__q)
    );
    wire _node_627;
    BITWISEAND #(.width(1)) bitwiseand_1208 (
        .y(_node_627),
        .a(1'h1),
        .b(_node_626)
    );
    wire [7:0] _GEN_324;
    MUX_UNSIGNED #(.width(8)) u_mux_1209 (
        .y(_GEN_324),
        .sel(_node_627),
        .a(helloWorld_314),
        .b(_GEN_323)
    );
    wire _node_628;
    EQ_UNSIGNED #(.width(9)) u_eq_1210 (
        .y(_node_628),
        .a(9'h13B),
        .b(_arrivedPointer__q)
    );
    wire _node_629;
    BITWISEAND #(.width(1)) bitwiseand_1211 (
        .y(_node_629),
        .a(1'h1),
        .b(_node_628)
    );
    wire [7:0] _GEN_325;
    MUX_UNSIGNED #(.width(8)) u_mux_1212 (
        .y(_GEN_325),
        .sel(_node_629),
        .a(helloWorld_315),
        .b(_GEN_324)
    );
    wire _node_630;
    EQ_UNSIGNED #(.width(9)) u_eq_1213 (
        .y(_node_630),
        .a(9'h13C),
        .b(_arrivedPointer__q)
    );
    wire _node_631;
    BITWISEAND #(.width(1)) bitwiseand_1214 (
        .y(_node_631),
        .a(1'h1),
        .b(_node_630)
    );
    wire [7:0] _GEN_326;
    MUX_UNSIGNED #(.width(8)) u_mux_1215 (
        .y(_GEN_326),
        .sel(_node_631),
        .a(helloWorld_316),
        .b(_GEN_325)
    );
    wire _node_632;
    EQ_UNSIGNED #(.width(9)) u_eq_1216 (
        .y(_node_632),
        .a(9'h13D),
        .b(_arrivedPointer__q)
    );
    wire _node_633;
    BITWISEAND #(.width(1)) bitwiseand_1217 (
        .y(_node_633),
        .a(1'h1),
        .b(_node_632)
    );
    wire [7:0] _GEN_327;
    MUX_UNSIGNED #(.width(8)) u_mux_1218 (
        .y(_GEN_327),
        .sel(_node_633),
        .a(helloWorld_317),
        .b(_GEN_326)
    );
    wire _node_634;
    EQ_UNSIGNED #(.width(9)) u_eq_1219 (
        .y(_node_634),
        .a(9'h13E),
        .b(_arrivedPointer__q)
    );
    wire _node_635;
    BITWISEAND #(.width(1)) bitwiseand_1220 (
        .y(_node_635),
        .a(1'h1),
        .b(_node_634)
    );
    wire [7:0] _GEN_328;
    MUX_UNSIGNED #(.width(8)) u_mux_1221 (
        .y(_GEN_328),
        .sel(_node_635),
        .a(helloWorld_318),
        .b(_GEN_327)
    );
    wire _node_636;
    EQ_UNSIGNED #(.width(9)) u_eq_1222 (
        .y(_node_636),
        .a(9'h13F),
        .b(_arrivedPointer__q)
    );
    wire _node_637;
    BITWISEAND #(.width(1)) bitwiseand_1223 (
        .y(_node_637),
        .a(1'h1),
        .b(_node_636)
    );
    wire [7:0] _GEN_329;
    MUX_UNSIGNED #(.width(8)) u_mux_1224 (
        .y(_GEN_329),
        .sel(_node_637),
        .a(helloWorld_319),
        .b(_GEN_328)
    );
    wire _node_638;
    EQ_UNSIGNED #(.width(9)) u_eq_1225 (
        .y(_node_638),
        .a(9'h140),
        .b(_arrivedPointer__q)
    );
    wire _node_639;
    BITWISEAND #(.width(1)) bitwiseand_1226 (
        .y(_node_639),
        .a(1'h1),
        .b(_node_638)
    );
    wire [7:0] _GEN_330;
    MUX_UNSIGNED #(.width(8)) u_mux_1227 (
        .y(_GEN_330),
        .sel(_node_639),
        .a(helloWorld_320),
        .b(_GEN_329)
    );
    wire _node_640;
    EQ_UNSIGNED #(.width(9)) u_eq_1228 (
        .y(_node_640),
        .a(9'h141),
        .b(_arrivedPointer__q)
    );
    wire _node_641;
    BITWISEAND #(.width(1)) bitwiseand_1229 (
        .y(_node_641),
        .a(1'h1),
        .b(_node_640)
    );
    wire [7:0] _GEN_331;
    MUX_UNSIGNED #(.width(8)) u_mux_1230 (
        .y(_GEN_331),
        .sel(_node_641),
        .a(helloWorld_321),
        .b(_GEN_330)
    );
    wire _node_642;
    EQ_UNSIGNED #(.width(9)) u_eq_1231 (
        .y(_node_642),
        .a(9'h142),
        .b(_arrivedPointer__q)
    );
    wire _node_643;
    BITWISEAND #(.width(1)) bitwiseand_1232 (
        .y(_node_643),
        .a(1'h1),
        .b(_node_642)
    );
    wire [7:0] _GEN_332;
    MUX_UNSIGNED #(.width(8)) u_mux_1233 (
        .y(_GEN_332),
        .sel(_node_643),
        .a(helloWorld_322),
        .b(_GEN_331)
    );
    wire _node_644;
    EQ_UNSIGNED #(.width(9)) u_eq_1234 (
        .y(_node_644),
        .a(9'h143),
        .b(_arrivedPointer__q)
    );
    wire _node_645;
    BITWISEAND #(.width(1)) bitwiseand_1235 (
        .y(_node_645),
        .a(1'h1),
        .b(_node_644)
    );
    wire [7:0] _GEN_333;
    MUX_UNSIGNED #(.width(8)) u_mux_1236 (
        .y(_GEN_333),
        .sel(_node_645),
        .a(helloWorld_323),
        .b(_GEN_332)
    );
    wire _node_646;
    EQ_UNSIGNED #(.width(9)) u_eq_1237 (
        .y(_node_646),
        .a(9'h144),
        .b(_arrivedPointer__q)
    );
    wire _node_647;
    BITWISEAND #(.width(1)) bitwiseand_1238 (
        .y(_node_647),
        .a(1'h1),
        .b(_node_646)
    );
    wire [7:0] _GEN_334;
    MUX_UNSIGNED #(.width(8)) u_mux_1239 (
        .y(_GEN_334),
        .sel(_node_647),
        .a(helloWorld_324),
        .b(_GEN_333)
    );
    wire _node_648;
    EQ_UNSIGNED #(.width(9)) u_eq_1240 (
        .y(_node_648),
        .a(9'h145),
        .b(_arrivedPointer__q)
    );
    wire _node_649;
    BITWISEAND #(.width(1)) bitwiseand_1241 (
        .y(_node_649),
        .a(1'h1),
        .b(_node_648)
    );
    wire [7:0] _GEN_335;
    MUX_UNSIGNED #(.width(8)) u_mux_1242 (
        .y(_GEN_335),
        .sel(_node_649),
        .a(helloWorld_325),
        .b(_GEN_334)
    );
    wire _node_650;
    EQ_UNSIGNED #(.width(9)) u_eq_1243 (
        .y(_node_650),
        .a(9'h146),
        .b(_arrivedPointer__q)
    );
    wire _node_651;
    BITWISEAND #(.width(1)) bitwiseand_1244 (
        .y(_node_651),
        .a(1'h1),
        .b(_node_650)
    );
    wire [7:0] _GEN_336;
    MUX_UNSIGNED #(.width(8)) u_mux_1245 (
        .y(_GEN_336),
        .sel(_node_651),
        .a(helloWorld_326),
        .b(_GEN_335)
    );
    wire _node_652;
    EQ_UNSIGNED #(.width(9)) u_eq_1246 (
        .y(_node_652),
        .a(9'h147),
        .b(_arrivedPointer__q)
    );
    wire _node_653;
    BITWISEAND #(.width(1)) bitwiseand_1247 (
        .y(_node_653),
        .a(1'h1),
        .b(_node_652)
    );
    wire [7:0] _GEN_337;
    MUX_UNSIGNED #(.width(8)) u_mux_1248 (
        .y(_GEN_337),
        .sel(_node_653),
        .a(helloWorld_327),
        .b(_GEN_336)
    );
    wire _node_654;
    EQ_UNSIGNED #(.width(9)) u_eq_1249 (
        .y(_node_654),
        .a(9'h148),
        .b(_arrivedPointer__q)
    );
    wire _node_655;
    BITWISEAND #(.width(1)) bitwiseand_1250 (
        .y(_node_655),
        .a(1'h1),
        .b(_node_654)
    );
    wire [7:0] _GEN_338;
    MUX_UNSIGNED #(.width(8)) u_mux_1251 (
        .y(_GEN_338),
        .sel(_node_655),
        .a(helloWorld_328),
        .b(_GEN_337)
    );
    wire _node_656;
    EQ_UNSIGNED #(.width(9)) u_eq_1252 (
        .y(_node_656),
        .a(9'h149),
        .b(_arrivedPointer__q)
    );
    wire _node_657;
    BITWISEAND #(.width(1)) bitwiseand_1253 (
        .y(_node_657),
        .a(1'h1),
        .b(_node_656)
    );
    wire [7:0] _GEN_339;
    MUX_UNSIGNED #(.width(8)) u_mux_1254 (
        .y(_GEN_339),
        .sel(_node_657),
        .a(helloWorld_329),
        .b(_GEN_338)
    );
    wire _node_658;
    EQ_UNSIGNED #(.width(9)) u_eq_1255 (
        .y(_node_658),
        .a(9'h14A),
        .b(_arrivedPointer__q)
    );
    wire _node_659;
    BITWISEAND #(.width(1)) bitwiseand_1256 (
        .y(_node_659),
        .a(1'h1),
        .b(_node_658)
    );
    wire [7:0] _GEN_340;
    MUX_UNSIGNED #(.width(8)) u_mux_1257 (
        .y(_GEN_340),
        .sel(_node_659),
        .a(helloWorld_330),
        .b(_GEN_339)
    );
    wire _node_660;
    EQ_UNSIGNED #(.width(9)) u_eq_1258 (
        .y(_node_660),
        .a(9'h14B),
        .b(_arrivedPointer__q)
    );
    wire _node_661;
    BITWISEAND #(.width(1)) bitwiseand_1259 (
        .y(_node_661),
        .a(1'h1),
        .b(_node_660)
    );
    wire [7:0] _GEN_341;
    MUX_UNSIGNED #(.width(8)) u_mux_1260 (
        .y(_GEN_341),
        .sel(_node_661),
        .a(helloWorld_331),
        .b(_GEN_340)
    );
    wire _node_662;
    EQ_UNSIGNED #(.width(9)) u_eq_1261 (
        .y(_node_662),
        .a(9'h14C),
        .b(_arrivedPointer__q)
    );
    wire _node_663;
    BITWISEAND #(.width(1)) bitwiseand_1262 (
        .y(_node_663),
        .a(1'h1),
        .b(_node_662)
    );
    wire [7:0] _GEN_342;
    MUX_UNSIGNED #(.width(8)) u_mux_1263 (
        .y(_GEN_342),
        .sel(_node_663),
        .a(helloWorld_332),
        .b(_GEN_341)
    );
    wire _node_664;
    EQ_UNSIGNED #(.width(9)) u_eq_1264 (
        .y(_node_664),
        .a(9'h14D),
        .b(_arrivedPointer__q)
    );
    wire _node_665;
    BITWISEAND #(.width(1)) bitwiseand_1265 (
        .y(_node_665),
        .a(1'h1),
        .b(_node_664)
    );
    wire [7:0] _GEN_343;
    MUX_UNSIGNED #(.width(8)) u_mux_1266 (
        .y(_GEN_343),
        .sel(_node_665),
        .a(helloWorld_333),
        .b(_GEN_342)
    );
    wire _node_666;
    EQ_UNSIGNED #(.width(9)) u_eq_1267 (
        .y(_node_666),
        .a(9'h14E),
        .b(_arrivedPointer__q)
    );
    wire _node_667;
    BITWISEAND #(.width(1)) bitwiseand_1268 (
        .y(_node_667),
        .a(1'h1),
        .b(_node_666)
    );
    wire [7:0] _GEN_344;
    MUX_UNSIGNED #(.width(8)) u_mux_1269 (
        .y(_GEN_344),
        .sel(_node_667),
        .a(helloWorld_334),
        .b(_GEN_343)
    );
    wire _node_668;
    EQ_UNSIGNED #(.width(9)) u_eq_1270 (
        .y(_node_668),
        .a(9'h14F),
        .b(_arrivedPointer__q)
    );
    wire _node_669;
    BITWISEAND #(.width(1)) bitwiseand_1271 (
        .y(_node_669),
        .a(1'h1),
        .b(_node_668)
    );
    wire [7:0] _GEN_345;
    MUX_UNSIGNED #(.width(8)) u_mux_1272 (
        .y(_GEN_345),
        .sel(_node_669),
        .a(helloWorld_335),
        .b(_GEN_344)
    );
    wire _node_670;
    EQ_UNSIGNED #(.width(9)) u_eq_1273 (
        .y(_node_670),
        .a(9'h150),
        .b(_arrivedPointer__q)
    );
    wire _node_671;
    BITWISEAND #(.width(1)) bitwiseand_1274 (
        .y(_node_671),
        .a(1'h1),
        .b(_node_670)
    );
    wire [7:0] _GEN_346;
    MUX_UNSIGNED #(.width(8)) u_mux_1275 (
        .y(_GEN_346),
        .sel(_node_671),
        .a(helloWorld_336),
        .b(_GEN_345)
    );
    wire _node_672;
    EQ_UNSIGNED #(.width(9)) u_eq_1276 (
        .y(_node_672),
        .a(9'h151),
        .b(_arrivedPointer__q)
    );
    wire _node_673;
    BITWISEAND #(.width(1)) bitwiseand_1277 (
        .y(_node_673),
        .a(1'h1),
        .b(_node_672)
    );
    wire [7:0] _GEN_347;
    MUX_UNSIGNED #(.width(8)) u_mux_1278 (
        .y(_GEN_347),
        .sel(_node_673),
        .a(helloWorld_337),
        .b(_GEN_346)
    );
    wire _node_674;
    EQ_UNSIGNED #(.width(9)) u_eq_1279 (
        .y(_node_674),
        .a(9'h152),
        .b(_arrivedPointer__q)
    );
    wire _node_675;
    BITWISEAND #(.width(1)) bitwiseand_1280 (
        .y(_node_675),
        .a(1'h1),
        .b(_node_674)
    );
    wire [7:0] _GEN_348;
    MUX_UNSIGNED #(.width(8)) u_mux_1281 (
        .y(_GEN_348),
        .sel(_node_675),
        .a(helloWorld_338),
        .b(_GEN_347)
    );
    wire _node_676;
    EQ_UNSIGNED #(.width(9)) u_eq_1282 (
        .y(_node_676),
        .a(9'h153),
        .b(_arrivedPointer__q)
    );
    wire _node_677;
    BITWISEAND #(.width(1)) bitwiseand_1283 (
        .y(_node_677),
        .a(1'h1),
        .b(_node_676)
    );
    wire [7:0] _GEN_349;
    MUX_UNSIGNED #(.width(8)) u_mux_1284 (
        .y(_GEN_349),
        .sel(_node_677),
        .a(helloWorld_339),
        .b(_GEN_348)
    );
    wire _node_678;
    EQ_UNSIGNED #(.width(9)) u_eq_1285 (
        .y(_node_678),
        .a(9'h154),
        .b(_arrivedPointer__q)
    );
    wire _node_679;
    BITWISEAND #(.width(1)) bitwiseand_1286 (
        .y(_node_679),
        .a(1'h1),
        .b(_node_678)
    );
    wire [7:0] _GEN_350;
    MUX_UNSIGNED #(.width(8)) u_mux_1287 (
        .y(_GEN_350),
        .sel(_node_679),
        .a(helloWorld_340),
        .b(_GEN_349)
    );
    wire _node_680;
    EQ_UNSIGNED #(.width(9)) u_eq_1288 (
        .y(_node_680),
        .a(9'h155),
        .b(_arrivedPointer__q)
    );
    wire _node_681;
    BITWISEAND #(.width(1)) bitwiseand_1289 (
        .y(_node_681),
        .a(1'h1),
        .b(_node_680)
    );
    wire [7:0] _GEN_351;
    MUX_UNSIGNED #(.width(8)) u_mux_1290 (
        .y(_GEN_351),
        .sel(_node_681),
        .a(helloWorld_341),
        .b(_GEN_350)
    );
    wire _node_682;
    EQ_UNSIGNED #(.width(9)) u_eq_1291 (
        .y(_node_682),
        .a(9'h156),
        .b(_arrivedPointer__q)
    );
    wire _node_683;
    BITWISEAND #(.width(1)) bitwiseand_1292 (
        .y(_node_683),
        .a(1'h1),
        .b(_node_682)
    );
    wire [7:0] _GEN_352;
    MUX_UNSIGNED #(.width(8)) u_mux_1293 (
        .y(_GEN_352),
        .sel(_node_683),
        .a(helloWorld_342),
        .b(_GEN_351)
    );
    wire _node_684;
    EQ_UNSIGNED #(.width(9)) u_eq_1294 (
        .y(_node_684),
        .a(9'h157),
        .b(_arrivedPointer__q)
    );
    wire _node_685;
    BITWISEAND #(.width(1)) bitwiseand_1295 (
        .y(_node_685),
        .a(1'h1),
        .b(_node_684)
    );
    wire [7:0] _GEN_353;
    MUX_UNSIGNED #(.width(8)) u_mux_1296 (
        .y(_GEN_353),
        .sel(_node_685),
        .a(helloWorld_343),
        .b(_GEN_352)
    );
    wire _node_686;
    EQ_UNSIGNED #(.width(9)) u_eq_1297 (
        .y(_node_686),
        .a(9'h158),
        .b(_arrivedPointer__q)
    );
    wire _node_687;
    BITWISEAND #(.width(1)) bitwiseand_1298 (
        .y(_node_687),
        .a(1'h1),
        .b(_node_686)
    );
    wire [7:0] _GEN_354;
    MUX_UNSIGNED #(.width(8)) u_mux_1299 (
        .y(_GEN_354),
        .sel(_node_687),
        .a(helloWorld_344),
        .b(_GEN_353)
    );
    wire _node_688;
    EQ_UNSIGNED #(.width(9)) u_eq_1300 (
        .y(_node_688),
        .a(9'h159),
        .b(_arrivedPointer__q)
    );
    wire _node_689;
    BITWISEAND #(.width(1)) bitwiseand_1301 (
        .y(_node_689),
        .a(1'h1),
        .b(_node_688)
    );
    wire [7:0] _GEN_355;
    MUX_UNSIGNED #(.width(8)) u_mux_1302 (
        .y(_GEN_355),
        .sel(_node_689),
        .a(helloWorld_345),
        .b(_GEN_354)
    );
    wire _node_690;
    EQ_UNSIGNED #(.width(9)) u_eq_1303 (
        .y(_node_690),
        .a(9'h15A),
        .b(_arrivedPointer__q)
    );
    wire _node_691;
    BITWISEAND #(.width(1)) bitwiseand_1304 (
        .y(_node_691),
        .a(1'h1),
        .b(_node_690)
    );
    wire [7:0] _GEN_356;
    MUX_UNSIGNED #(.width(8)) u_mux_1305 (
        .y(_GEN_356),
        .sel(_node_691),
        .a(helloWorld_346),
        .b(_GEN_355)
    );
    wire _node_692;
    EQ_UNSIGNED #(.width(9)) u_eq_1306 (
        .y(_node_692),
        .a(9'h15B),
        .b(_arrivedPointer__q)
    );
    wire _node_693;
    BITWISEAND #(.width(1)) bitwiseand_1307 (
        .y(_node_693),
        .a(1'h1),
        .b(_node_692)
    );
    wire [7:0] _GEN_357;
    MUX_UNSIGNED #(.width(8)) u_mux_1308 (
        .y(_GEN_357),
        .sel(_node_693),
        .a(helloWorld_347),
        .b(_GEN_356)
    );
    wire _node_694;
    EQ_UNSIGNED #(.width(9)) u_eq_1309 (
        .y(_node_694),
        .a(9'h15C),
        .b(_arrivedPointer__q)
    );
    wire _node_695;
    BITWISEAND #(.width(1)) bitwiseand_1310 (
        .y(_node_695),
        .a(1'h1),
        .b(_node_694)
    );
    wire [7:0] _GEN_358;
    MUX_UNSIGNED #(.width(8)) u_mux_1311 (
        .y(_GEN_358),
        .sel(_node_695),
        .a(helloWorld_348),
        .b(_GEN_357)
    );
    wire _node_696;
    EQ_UNSIGNED #(.width(9)) u_eq_1312 (
        .y(_node_696),
        .a(9'h15D),
        .b(_arrivedPointer__q)
    );
    wire _node_697;
    BITWISEAND #(.width(1)) bitwiseand_1313 (
        .y(_node_697),
        .a(1'h1),
        .b(_node_696)
    );
    wire [7:0] _GEN_359;
    MUX_UNSIGNED #(.width(8)) u_mux_1314 (
        .y(_GEN_359),
        .sel(_node_697),
        .a(helloWorld_349),
        .b(_GEN_358)
    );
    wire _node_698;
    EQ_UNSIGNED #(.width(9)) u_eq_1315 (
        .y(_node_698),
        .a(9'h15E),
        .b(_arrivedPointer__q)
    );
    wire _node_699;
    BITWISEAND #(.width(1)) bitwiseand_1316 (
        .y(_node_699),
        .a(1'h1),
        .b(_node_698)
    );
    wire [7:0] _GEN_360;
    MUX_UNSIGNED #(.width(8)) u_mux_1317 (
        .y(_GEN_360),
        .sel(_node_699),
        .a(helloWorld_350),
        .b(_GEN_359)
    );
    wire _node_700;
    EQ_UNSIGNED #(.width(9)) u_eq_1318 (
        .y(_node_700),
        .a(9'h15F),
        .b(_arrivedPointer__q)
    );
    wire _node_701;
    BITWISEAND #(.width(1)) bitwiseand_1319 (
        .y(_node_701),
        .a(1'h1),
        .b(_node_700)
    );
    wire [7:0] _GEN_361;
    MUX_UNSIGNED #(.width(8)) u_mux_1320 (
        .y(_GEN_361),
        .sel(_node_701),
        .a(helloWorld_351),
        .b(_GEN_360)
    );
    wire _node_702;
    EQ_UNSIGNED #(.width(9)) u_eq_1321 (
        .y(_node_702),
        .a(9'h160),
        .b(_arrivedPointer__q)
    );
    wire _node_703;
    BITWISEAND #(.width(1)) bitwiseand_1322 (
        .y(_node_703),
        .a(1'h1),
        .b(_node_702)
    );
    wire [7:0] _GEN_362;
    MUX_UNSIGNED #(.width(8)) u_mux_1323 (
        .y(_GEN_362),
        .sel(_node_703),
        .a(helloWorld_352),
        .b(_GEN_361)
    );
    wire _node_704;
    EQ_UNSIGNED #(.width(9)) u_eq_1324 (
        .y(_node_704),
        .a(9'h161),
        .b(_arrivedPointer__q)
    );
    wire _node_705;
    BITWISEAND #(.width(1)) bitwiseand_1325 (
        .y(_node_705),
        .a(1'h1),
        .b(_node_704)
    );
    wire [7:0] _GEN_363;
    MUX_UNSIGNED #(.width(8)) u_mux_1326 (
        .y(_GEN_363),
        .sel(_node_705),
        .a(helloWorld_353),
        .b(_GEN_362)
    );
    wire _node_706;
    EQ_UNSIGNED #(.width(9)) u_eq_1327 (
        .y(_node_706),
        .a(9'h162),
        .b(_arrivedPointer__q)
    );
    wire _node_707;
    BITWISEAND #(.width(1)) bitwiseand_1328 (
        .y(_node_707),
        .a(1'h1),
        .b(_node_706)
    );
    wire [7:0] _GEN_364;
    MUX_UNSIGNED #(.width(8)) u_mux_1329 (
        .y(_GEN_364),
        .sel(_node_707),
        .a(helloWorld_354),
        .b(_GEN_363)
    );
    wire _node_708;
    EQ_UNSIGNED #(.width(9)) u_eq_1330 (
        .y(_node_708),
        .a(9'h163),
        .b(_arrivedPointer__q)
    );
    wire _node_709;
    BITWISEAND #(.width(1)) bitwiseand_1331 (
        .y(_node_709),
        .a(1'h1),
        .b(_node_708)
    );
    wire [7:0] _GEN_365;
    MUX_UNSIGNED #(.width(8)) u_mux_1332 (
        .y(_GEN_365),
        .sel(_node_709),
        .a(helloWorld_355),
        .b(_GEN_364)
    );
    wire _node_710;
    EQ_UNSIGNED #(.width(9)) u_eq_1333 (
        .y(_node_710),
        .a(9'h164),
        .b(_arrivedPointer__q)
    );
    wire _node_711;
    BITWISEAND #(.width(1)) bitwiseand_1334 (
        .y(_node_711),
        .a(1'h1),
        .b(_node_710)
    );
    wire [7:0] _GEN_366;
    MUX_UNSIGNED #(.width(8)) u_mux_1335 (
        .y(_GEN_366),
        .sel(_node_711),
        .a(helloWorld_356),
        .b(_GEN_365)
    );
    wire _node_712;
    EQ_UNSIGNED #(.width(9)) u_eq_1336 (
        .y(_node_712),
        .a(9'h165),
        .b(_arrivedPointer__q)
    );
    wire _node_713;
    BITWISEAND #(.width(1)) bitwiseand_1337 (
        .y(_node_713),
        .a(1'h1),
        .b(_node_712)
    );
    wire [7:0] _GEN_367;
    MUX_UNSIGNED #(.width(8)) u_mux_1338 (
        .y(_GEN_367),
        .sel(_node_713),
        .a(helloWorld_357),
        .b(_GEN_366)
    );
    wire _node_714;
    EQ_UNSIGNED #(.width(9)) u_eq_1339 (
        .y(_node_714),
        .a(9'h166),
        .b(_arrivedPointer__q)
    );
    wire _node_715;
    BITWISEAND #(.width(1)) bitwiseand_1340 (
        .y(_node_715),
        .a(1'h1),
        .b(_node_714)
    );
    wire [7:0] _GEN_368;
    MUX_UNSIGNED #(.width(8)) u_mux_1341 (
        .y(_GEN_368),
        .sel(_node_715),
        .a(helloWorld_358),
        .b(_GEN_367)
    );
    wire _node_716;
    EQ_UNSIGNED #(.width(9)) u_eq_1342 (
        .y(_node_716),
        .a(9'h167),
        .b(_arrivedPointer__q)
    );
    wire _node_717;
    BITWISEAND #(.width(1)) bitwiseand_1343 (
        .y(_node_717),
        .a(1'h1),
        .b(_node_716)
    );
    wire [7:0] _GEN_369;
    MUX_UNSIGNED #(.width(8)) u_mux_1344 (
        .y(_GEN_369),
        .sel(_node_717),
        .a(helloWorld_359),
        .b(_GEN_368)
    );
    wire _node_718;
    EQ_UNSIGNED #(.width(9)) u_eq_1345 (
        .y(_node_718),
        .a(9'h168),
        .b(_arrivedPointer__q)
    );
    wire _node_719;
    BITWISEAND #(.width(1)) bitwiseand_1346 (
        .y(_node_719),
        .a(1'h1),
        .b(_node_718)
    );
    wire [7:0] _GEN_370;
    MUX_UNSIGNED #(.width(8)) u_mux_1347 (
        .y(_GEN_370),
        .sel(_node_719),
        .a(helloWorld_360),
        .b(_GEN_369)
    );
    wire _node_720;
    EQ_UNSIGNED #(.width(9)) u_eq_1348 (
        .y(_node_720),
        .a(9'h169),
        .b(_arrivedPointer__q)
    );
    wire _node_721;
    BITWISEAND #(.width(1)) bitwiseand_1349 (
        .y(_node_721),
        .a(1'h1),
        .b(_node_720)
    );
    wire [7:0] _GEN_371;
    MUX_UNSIGNED #(.width(8)) u_mux_1350 (
        .y(_GEN_371),
        .sel(_node_721),
        .a(helloWorld_361),
        .b(_GEN_370)
    );
    wire _node_722;
    EQ_UNSIGNED #(.width(9)) u_eq_1351 (
        .y(_node_722),
        .a(9'h16A),
        .b(_arrivedPointer__q)
    );
    wire _node_723;
    BITWISEAND #(.width(1)) bitwiseand_1352 (
        .y(_node_723),
        .a(1'h1),
        .b(_node_722)
    );
    wire [7:0] _GEN_372;
    MUX_UNSIGNED #(.width(8)) u_mux_1353 (
        .y(_GEN_372),
        .sel(_node_723),
        .a(helloWorld_362),
        .b(_GEN_371)
    );
    wire _node_724;
    EQ_UNSIGNED #(.width(9)) u_eq_1354 (
        .y(_node_724),
        .a(9'h16B),
        .b(_arrivedPointer__q)
    );
    wire _node_725;
    BITWISEAND #(.width(1)) bitwiseand_1355 (
        .y(_node_725),
        .a(1'h1),
        .b(_node_724)
    );
    wire [7:0] _GEN_373;
    MUX_UNSIGNED #(.width(8)) u_mux_1356 (
        .y(_GEN_373),
        .sel(_node_725),
        .a(helloWorld_363),
        .b(_GEN_372)
    );
    wire _node_726;
    EQ_UNSIGNED #(.width(9)) u_eq_1357 (
        .y(_node_726),
        .a(9'h16C),
        .b(_arrivedPointer__q)
    );
    wire _node_727;
    BITWISEAND #(.width(1)) bitwiseand_1358 (
        .y(_node_727),
        .a(1'h1),
        .b(_node_726)
    );
    wire [7:0] _GEN_374;
    MUX_UNSIGNED #(.width(8)) u_mux_1359 (
        .y(_GEN_374),
        .sel(_node_727),
        .a(helloWorld_364),
        .b(_GEN_373)
    );
    wire _node_728;
    EQ_UNSIGNED #(.width(9)) u_eq_1360 (
        .y(_node_728),
        .a(9'h16D),
        .b(_arrivedPointer__q)
    );
    wire _node_729;
    BITWISEAND #(.width(1)) bitwiseand_1361 (
        .y(_node_729),
        .a(1'h1),
        .b(_node_728)
    );
    wire [7:0] _GEN_375;
    MUX_UNSIGNED #(.width(8)) u_mux_1362 (
        .y(_GEN_375),
        .sel(_node_729),
        .a(helloWorld_365),
        .b(_GEN_374)
    );
    wire _node_730;
    EQ_UNSIGNED #(.width(9)) u_eq_1363 (
        .y(_node_730),
        .a(9'h16E),
        .b(_arrivedPointer__q)
    );
    wire _node_731;
    BITWISEAND #(.width(1)) bitwiseand_1364 (
        .y(_node_731),
        .a(1'h1),
        .b(_node_730)
    );
    wire [7:0] _GEN_376;
    MUX_UNSIGNED #(.width(8)) u_mux_1365 (
        .y(_GEN_376),
        .sel(_node_731),
        .a(helloWorld_366),
        .b(_GEN_375)
    );
    wire _node_732;
    EQ_UNSIGNED #(.width(9)) u_eq_1366 (
        .y(_node_732),
        .a(9'h16F),
        .b(_arrivedPointer__q)
    );
    wire _node_733;
    BITWISEAND #(.width(1)) bitwiseand_1367 (
        .y(_node_733),
        .a(1'h1),
        .b(_node_732)
    );
    wire [7:0] _GEN_377;
    MUX_UNSIGNED #(.width(8)) u_mux_1368 (
        .y(_GEN_377),
        .sel(_node_733),
        .a(helloWorld_367),
        .b(_GEN_376)
    );
    wire _node_734;
    EQ_UNSIGNED #(.width(9)) u_eq_1369 (
        .y(_node_734),
        .a(9'h170),
        .b(_arrivedPointer__q)
    );
    wire _node_735;
    BITWISEAND #(.width(1)) bitwiseand_1370 (
        .y(_node_735),
        .a(1'h1),
        .b(_node_734)
    );
    wire [7:0] _GEN_378;
    MUX_UNSIGNED #(.width(8)) u_mux_1371 (
        .y(_GEN_378),
        .sel(_node_735),
        .a(helloWorld_368),
        .b(_GEN_377)
    );
    wire _node_736;
    EQ_UNSIGNED #(.width(9)) u_eq_1372 (
        .y(_node_736),
        .a(9'h171),
        .b(_arrivedPointer__q)
    );
    wire _node_737;
    BITWISEAND #(.width(1)) bitwiseand_1373 (
        .y(_node_737),
        .a(1'h1),
        .b(_node_736)
    );
    wire [7:0] _GEN_379;
    MUX_UNSIGNED #(.width(8)) u_mux_1374 (
        .y(_GEN_379),
        .sel(_node_737),
        .a(helloWorld_369),
        .b(_GEN_378)
    );
    wire _node_738;
    EQ_UNSIGNED #(.width(9)) u_eq_1375 (
        .y(_node_738),
        .a(9'h172),
        .b(_arrivedPointer__q)
    );
    wire _node_739;
    BITWISEAND #(.width(1)) bitwiseand_1376 (
        .y(_node_739),
        .a(1'h1),
        .b(_node_738)
    );
    wire [7:0] _GEN_380;
    MUX_UNSIGNED #(.width(8)) u_mux_1377 (
        .y(_GEN_380),
        .sel(_node_739),
        .a(helloWorld_370),
        .b(_GEN_379)
    );
    wire _node_740;
    EQ_UNSIGNED #(.width(9)) u_eq_1378 (
        .y(_node_740),
        .a(9'h173),
        .b(_arrivedPointer__q)
    );
    wire _node_741;
    BITWISEAND #(.width(1)) bitwiseand_1379 (
        .y(_node_741),
        .a(1'h1),
        .b(_node_740)
    );
    wire [7:0] _GEN_381;
    MUX_UNSIGNED #(.width(8)) u_mux_1380 (
        .y(_GEN_381),
        .sel(_node_741),
        .a(helloWorld_371),
        .b(_GEN_380)
    );
    wire _node_742;
    EQ_UNSIGNED #(.width(9)) u_eq_1381 (
        .y(_node_742),
        .a(9'h174),
        .b(_arrivedPointer__q)
    );
    wire _node_743;
    BITWISEAND #(.width(1)) bitwiseand_1382 (
        .y(_node_743),
        .a(1'h1),
        .b(_node_742)
    );
    wire [7:0] _GEN_382;
    MUX_UNSIGNED #(.width(8)) u_mux_1383 (
        .y(_GEN_382),
        .sel(_node_743),
        .a(helloWorld_372),
        .b(_GEN_381)
    );
    wire _node_744;
    EQ_UNSIGNED #(.width(9)) u_eq_1384 (
        .y(_node_744),
        .a(9'h175),
        .b(_arrivedPointer__q)
    );
    wire _node_745;
    BITWISEAND #(.width(1)) bitwiseand_1385 (
        .y(_node_745),
        .a(1'h1),
        .b(_node_744)
    );
    wire [7:0] _GEN_383;
    MUX_UNSIGNED #(.width(8)) u_mux_1386 (
        .y(_GEN_383),
        .sel(_node_745),
        .a(helloWorld_373),
        .b(_GEN_382)
    );
    wire _node_746;
    EQ_UNSIGNED #(.width(9)) u_eq_1387 (
        .y(_node_746),
        .a(9'h176),
        .b(_arrivedPointer__q)
    );
    wire _node_747;
    BITWISEAND #(.width(1)) bitwiseand_1388 (
        .y(_node_747),
        .a(1'h1),
        .b(_node_746)
    );
    wire [7:0] _GEN_384;
    MUX_UNSIGNED #(.width(8)) u_mux_1389 (
        .y(_GEN_384),
        .sel(_node_747),
        .a(helloWorld_374),
        .b(_GEN_383)
    );
    wire _node_748;
    EQ_UNSIGNED #(.width(9)) u_eq_1390 (
        .y(_node_748),
        .a(9'h177),
        .b(_arrivedPointer__q)
    );
    wire _node_749;
    BITWISEAND #(.width(1)) bitwiseand_1391 (
        .y(_node_749),
        .a(1'h1),
        .b(_node_748)
    );
    wire [7:0] _GEN_385;
    MUX_UNSIGNED #(.width(8)) u_mux_1392 (
        .y(_GEN_385),
        .sel(_node_749),
        .a(helloWorld_375),
        .b(_GEN_384)
    );
    wire _node_750;
    EQ_UNSIGNED #(.width(9)) u_eq_1393 (
        .y(_node_750),
        .a(9'h178),
        .b(_arrivedPointer__q)
    );
    wire _node_751;
    BITWISEAND #(.width(1)) bitwiseand_1394 (
        .y(_node_751),
        .a(1'h1),
        .b(_node_750)
    );
    wire [7:0] _GEN_386;
    MUX_UNSIGNED #(.width(8)) u_mux_1395 (
        .y(_GEN_386),
        .sel(_node_751),
        .a(helloWorld_376),
        .b(_GEN_385)
    );
    wire _node_752;
    EQ_UNSIGNED #(.width(9)) u_eq_1396 (
        .y(_node_752),
        .a(9'h179),
        .b(_arrivedPointer__q)
    );
    wire _node_753;
    BITWISEAND #(.width(1)) bitwiseand_1397 (
        .y(_node_753),
        .a(1'h1),
        .b(_node_752)
    );
    wire [7:0] _GEN_387;
    MUX_UNSIGNED #(.width(8)) u_mux_1398 (
        .y(_GEN_387),
        .sel(_node_753),
        .a(helloWorld_377),
        .b(_GEN_386)
    );
    wire _node_754;
    EQ_UNSIGNED #(.width(9)) u_eq_1399 (
        .y(_node_754),
        .a(9'h17A),
        .b(_arrivedPointer__q)
    );
    wire _node_755;
    BITWISEAND #(.width(1)) bitwiseand_1400 (
        .y(_node_755),
        .a(1'h1),
        .b(_node_754)
    );
    wire [7:0] _GEN_388;
    MUX_UNSIGNED #(.width(8)) u_mux_1401 (
        .y(_GEN_388),
        .sel(_node_755),
        .a(helloWorld_378),
        .b(_GEN_387)
    );
    wire _node_756;
    EQ_UNSIGNED #(.width(9)) u_eq_1402 (
        .y(_node_756),
        .a(9'h17B),
        .b(_arrivedPointer__q)
    );
    wire _node_757;
    BITWISEAND #(.width(1)) bitwiseand_1403 (
        .y(_node_757),
        .a(1'h1),
        .b(_node_756)
    );
    wire [7:0] _GEN_389;
    MUX_UNSIGNED #(.width(8)) u_mux_1404 (
        .y(_GEN_389),
        .sel(_node_757),
        .a(helloWorld_379),
        .b(_GEN_388)
    );
    wire _node_758;
    EQ_UNSIGNED #(.width(9)) u_eq_1405 (
        .y(_node_758),
        .a(9'h17C),
        .b(_arrivedPointer__q)
    );
    wire _node_759;
    BITWISEAND #(.width(1)) bitwiseand_1406 (
        .y(_node_759),
        .a(1'h1),
        .b(_node_758)
    );
    wire [7:0] _GEN_390;
    MUX_UNSIGNED #(.width(8)) u_mux_1407 (
        .y(_GEN_390),
        .sel(_node_759),
        .a(helloWorld_380),
        .b(_GEN_389)
    );
    wire _node_760;
    EQ_UNSIGNED #(.width(9)) u_eq_1408 (
        .y(_node_760),
        .a(9'h17D),
        .b(_arrivedPointer__q)
    );
    wire _node_761;
    BITWISEAND #(.width(1)) bitwiseand_1409 (
        .y(_node_761),
        .a(1'h1),
        .b(_node_760)
    );
    wire [7:0] _GEN_391;
    MUX_UNSIGNED #(.width(8)) u_mux_1410 (
        .y(_GEN_391),
        .sel(_node_761),
        .a(helloWorld_381),
        .b(_GEN_390)
    );
    wire _node_762;
    EQ_UNSIGNED #(.width(9)) u_eq_1411 (
        .y(_node_762),
        .a(9'h17E),
        .b(_arrivedPointer__q)
    );
    wire _node_763;
    BITWISEAND #(.width(1)) bitwiseand_1412 (
        .y(_node_763),
        .a(1'h1),
        .b(_node_762)
    );
    wire [7:0] _GEN_392;
    MUX_UNSIGNED #(.width(8)) u_mux_1413 (
        .y(_GEN_392),
        .sel(_node_763),
        .a(helloWorld_382),
        .b(_GEN_391)
    );
    wire _node_764;
    EQ_UNSIGNED #(.width(9)) u_eq_1414 (
        .y(_node_764),
        .a(9'h17F),
        .b(_arrivedPointer__q)
    );
    wire _node_765;
    BITWISEAND #(.width(1)) bitwiseand_1415 (
        .y(_node_765),
        .a(1'h1),
        .b(_node_764)
    );
    wire [7:0] _GEN_393;
    MUX_UNSIGNED #(.width(8)) u_mux_1416 (
        .y(_GEN_393),
        .sel(_node_765),
        .a(helloWorld_383),
        .b(_GEN_392)
    );
    wire _node_766;
    EQ_UNSIGNED #(.width(9)) u_eq_1417 (
        .y(_node_766),
        .a(9'h180),
        .b(_arrivedPointer__q)
    );
    wire _node_767;
    BITWISEAND #(.width(1)) bitwiseand_1418 (
        .y(_node_767),
        .a(1'h1),
        .b(_node_766)
    );
    wire [7:0] _GEN_394;
    MUX_UNSIGNED #(.width(8)) u_mux_1419 (
        .y(_GEN_394),
        .sel(_node_767),
        .a(helloWorld_384),
        .b(_GEN_393)
    );
    wire _node_768;
    EQ_UNSIGNED #(.width(9)) u_eq_1420 (
        .y(_node_768),
        .a(9'h181),
        .b(_arrivedPointer__q)
    );
    wire _node_769;
    BITWISEAND #(.width(1)) bitwiseand_1421 (
        .y(_node_769),
        .a(1'h1),
        .b(_node_768)
    );
    wire [7:0] _GEN_395;
    MUX_UNSIGNED #(.width(8)) u_mux_1422 (
        .y(_GEN_395),
        .sel(_node_769),
        .a(helloWorld_385),
        .b(_GEN_394)
    );
    wire _node_770;
    EQ_UNSIGNED #(.width(9)) u_eq_1423 (
        .y(_node_770),
        .a(9'h182),
        .b(_arrivedPointer__q)
    );
    wire _node_771;
    BITWISEAND #(.width(1)) bitwiseand_1424 (
        .y(_node_771),
        .a(1'h1),
        .b(_node_770)
    );
    wire [7:0] _GEN_396;
    MUX_UNSIGNED #(.width(8)) u_mux_1425 (
        .y(_GEN_396),
        .sel(_node_771),
        .a(helloWorld_386),
        .b(_GEN_395)
    );
    wire _node_772;
    EQ_UNSIGNED #(.width(9)) u_eq_1426 (
        .y(_node_772),
        .a(9'h183),
        .b(_arrivedPointer__q)
    );
    wire _node_773;
    BITWISEAND #(.width(1)) bitwiseand_1427 (
        .y(_node_773),
        .a(1'h1),
        .b(_node_772)
    );
    wire [7:0] _GEN_397;
    MUX_UNSIGNED #(.width(8)) u_mux_1428 (
        .y(_GEN_397),
        .sel(_node_773),
        .a(helloWorld_387),
        .b(_GEN_396)
    );
    assign _GEN_0 = _GEN_397;
    assign __T_807__d = _GEN_5;
    assign __T_809__d = _GEN_6;
    assign __T_811__d = _GEN_7;
    assign __T_813__d = _GEN_8;
    assign __T_815__d = _GEN_9;
    MUX_UNSIGNED #(.width(9)) u_mux_1429 (
        .y(_arrivedPointer__d),
        .sel(reset),
        .a(9'h0),
        .b(_GEN_4)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_1430 (
        .y(_characterArrived__d),
        .sel(reset),
        .a(1'h0),
        .b(_GEN_10)
    );
    assign helloWorld_0 = 8'h57;
    assign helloWorld_1 = 8'h65;
    assign helloWorld_10 = 8'h74;
    assign helloWorld_100 = 8'h20;
    assign helloWorld_101 = 8'h62;
    assign helloWorld_102 = 8'h65;
    assign helloWorld_103 = 8'h63;
    assign helloWorld_104 = 8'h61;
    assign helloWorld_105 = 8'h75;
    assign helloWorld_106 = 8'h73;
    assign helloWorld_107 = 8'h65;
    assign helloWorld_108 = 8'h20;
    assign helloWorld_109 = 8'h74;
    assign helloWorld_11 = 8'h6F;
    assign helloWorld_110 = 8'h68;
    assign helloWorld_111 = 8'h65;
    assign helloWorld_112 = 8'h79;
    assign helloWorld_113 = 8'h20;
    assign helloWorld_114 = 8'h61;
    assign helloWorld_115 = 8'h72;
    assign helloWorld_116 = 8'h65;
    assign helloWorld_117 = 8'h20;
    assign helloWorld_118 = 8'h65;
    assign helloWorld_119 = 8'h61;
    assign helloWorld_12 = 8'h20;
    assign helloWorld_120 = 8'h73;
    assign helloWorld_121 = 8'h79;
    assign helloWorld_122 = 8'h2C;
    assign helloWorld_123 = 8'h20;
    assign helloWorld_124 = 8'h62;
    assign helloWorld_125 = 8'h75;
    assign helloWorld_126 = 8'h74;
    assign helloWorld_127 = 8'h20;
    assign helloWorld_128 = 8'h62;
    assign helloWorld_129 = 8'h65;
    assign helloWorld_13 = 8'h67;
    assign helloWorld_130 = 8'h63;
    assign helloWorld_131 = 8'h61;
    assign helloWorld_132 = 8'h75;
    assign helloWorld_133 = 8'h73;
    assign helloWorld_134 = 8'h65;
    assign helloWorld_135 = 8'h20;
    assign helloWorld_136 = 8'h74;
    assign helloWorld_137 = 8'h68;
    assign helloWorld_138 = 8'h65;
    assign helloWorld_139 = 8'h79;
    assign helloWorld_14 = 8'h6F;
    assign helloWorld_140 = 8'h20;
    assign helloWorld_141 = 8'h61;
    assign helloWorld_142 = 8'h72;
    assign helloWorld_143 = 8'h65;
    assign helloWorld_144 = 8'h20;
    assign helloWorld_145 = 8'h68;
    assign helloWorld_146 = 8'h61;
    assign helloWorld_147 = 8'h72;
    assign helloWorld_148 = 8'h64;
    assign helloWorld_149 = 8'h2C;
    assign helloWorld_15 = 8'h20;
    assign helloWorld_150 = 8'h20;
    assign helloWorld_151 = 8'h62;
    assign helloWorld_152 = 8'h65;
    assign helloWorld_153 = 8'h63;
    assign helloWorld_154 = 8'h61;
    assign helloWorld_155 = 8'h75;
    assign helloWorld_156 = 8'h73;
    assign helloWorld_157 = 8'h65;
    assign helloWorld_158 = 8'h20;
    assign helloWorld_159 = 8'h74;
    assign helloWorld_16 = 8'h74;
    assign helloWorld_160 = 8'h68;
    assign helloWorld_161 = 8'h61;
    assign helloWorld_162 = 8'h74;
    assign helloWorld_163 = 8'h20;
    assign helloWorld_164 = 8'h67;
    assign helloWorld_165 = 8'h6F;
    assign helloWorld_166 = 8'h61;
    assign helloWorld_167 = 8'h6C;
    assign helloWorld_168 = 8'h20;
    assign helloWorld_169 = 8'h77;
    assign helloWorld_17 = 8'h6F;
    assign helloWorld_170 = 8'h69;
    assign helloWorld_171 = 8'h6C;
    assign helloWorld_172 = 8'h6C;
    assign helloWorld_173 = 8'h20;
    assign helloWorld_174 = 8'h73;
    assign helloWorld_175 = 8'h65;
    assign helloWorld_176 = 8'h72;
    assign helloWorld_177 = 8'h76;
    assign helloWorld_178 = 8'h65;
    assign helloWorld_179 = 8'h20;
    assign helloWorld_18 = 8'h20;
    assign helloWorld_180 = 8'h74;
    assign helloWorld_181 = 8'h6F;
    assign helloWorld_182 = 8'h20;
    assign helloWorld_183 = 8'h6F;
    assign helloWorld_184 = 8'h72;
    assign helloWorld_185 = 8'h67;
    assign helloWorld_186 = 8'h61;
    assign helloWorld_187 = 8'h6E;
    assign helloWorld_188 = 8'h69;
    assign helloWorld_189 = 8'h7A;
    assign helloWorld_19 = 8'h74;
    assign helloWorld_190 = 8'h65;
    assign helloWorld_191 = 8'h20;
    assign helloWorld_192 = 8'h61;
    assign helloWorld_193 = 8'h6E;
    assign helloWorld_194 = 8'h64;
    assign helloWorld_195 = 8'h20;
    assign helloWorld_196 = 8'h6D;
    assign helloWorld_197 = 8'h65;
    assign helloWorld_198 = 8'h61;
    assign helloWorld_199 = 8'h73;
    assign helloWorld_2 = 8'h20;
    assign helloWorld_20 = 8'h68;
    assign helloWorld_200 = 8'h75;
    assign helloWorld_201 = 8'h72;
    assign helloWorld_202 = 8'h65;
    assign helloWorld_203 = 8'h20;
    assign helloWorld_204 = 8'h74;
    assign helloWorld_205 = 8'h68;
    assign helloWorld_206 = 8'h65;
    assign helloWorld_207 = 8'h20;
    assign helloWorld_208 = 8'h62;
    assign helloWorld_209 = 8'h65;
    assign helloWorld_21 = 8'h65;
    assign helloWorld_210 = 8'h73;
    assign helloWorld_211 = 8'h74;
    assign helloWorld_212 = 8'h20;
    assign helloWorld_213 = 8'h6F;
    assign helloWorld_214 = 8'h66;
    assign helloWorld_215 = 8'h20;
    assign helloWorld_216 = 8'h6F;
    assign helloWorld_217 = 8'h75;
    assign helloWorld_218 = 8'h72;
    assign helloWorld_219 = 8'h20;
    assign helloWorld_22 = 8'h20;
    assign helloWorld_220 = 8'h65;
    assign helloWorld_221 = 8'h6E;
    assign helloWorld_222 = 8'h65;
    assign helloWorld_223 = 8'h72;
    assign helloWorld_224 = 8'h67;
    assign helloWorld_225 = 8'h69;
    assign helloWorld_226 = 8'h65;
    assign helloWorld_227 = 8'h73;
    assign helloWorld_228 = 8'h20;
    assign helloWorld_229 = 8'h61;
    assign helloWorld_23 = 8'h6D;
    assign helloWorld_230 = 8'h6E;
    assign helloWorld_231 = 8'h64;
    assign helloWorld_232 = 8'h20;
    assign helloWorld_233 = 8'h73;
    assign helloWorld_234 = 8'h6B;
    assign helloWorld_235 = 8'h69;
    assign helloWorld_236 = 8'h6C;
    assign helloWorld_237 = 8'h6C;
    assign helloWorld_238 = 8'h73;
    assign helloWorld_239 = 8'h2C;
    assign helloWorld_24 = 8'h6F;
    assign helloWorld_240 = 8'h20;
    assign helloWorld_241 = 8'h62;
    assign helloWorld_242 = 8'h65;
    assign helloWorld_243 = 8'h63;
    assign helloWorld_244 = 8'h61;
    assign helloWorld_245 = 8'h75;
    assign helloWorld_246 = 8'h73;
    assign helloWorld_247 = 8'h65;
    assign helloWorld_248 = 8'h20;
    assign helloWorld_249 = 8'h74;
    assign helloWorld_25 = 8'h6F;
    assign helloWorld_250 = 8'h68;
    assign helloWorld_251 = 8'h61;
    assign helloWorld_252 = 8'h74;
    assign helloWorld_253 = 8'h20;
    assign helloWorld_254 = 8'h63;
    assign helloWorld_255 = 8'h68;
    assign helloWorld_256 = 8'h61;
    assign helloWorld_257 = 8'h6C;
    assign helloWorld_258 = 8'h6C;
    assign helloWorld_259 = 8'h65;
    assign helloWorld_26 = 8'h6E;
    assign helloWorld_260 = 8'h6E;
    assign helloWorld_261 = 8'h67;
    assign helloWorld_262 = 8'h65;
    assign helloWorld_263 = 8'h20;
    assign helloWorld_264 = 8'h69;
    assign helloWorld_265 = 8'h73;
    assign helloWorld_266 = 8'h20;
    assign helloWorld_267 = 8'h6F;
    assign helloWorld_268 = 8'h6E;
    assign helloWorld_269 = 8'h65;
    assign helloWorld_27 = 8'h2E;
    assign helloWorld_270 = 8'h20;
    assign helloWorld_271 = 8'h74;
    assign helloWorld_272 = 8'h68;
    assign helloWorld_273 = 8'h61;
    assign helloWorld_274 = 8'h74;
    assign helloWorld_275 = 8'h20;
    assign helloWorld_276 = 8'h77;
    assign helloWorld_277 = 8'h65;
    assign helloWorld_278 = 8'h20;
    assign helloWorld_279 = 8'h61;
    assign helloWorld_28 = 8'h20;
    assign helloWorld_280 = 8'h72;
    assign helloWorld_281 = 8'h65;
    assign helloWorld_282 = 8'h20;
    assign helloWorld_283 = 8'h77;
    assign helloWorld_284 = 8'h69;
    assign helloWorld_285 = 8'h6C;
    assign helloWorld_286 = 8'h6C;
    assign helloWorld_287 = 8'h69;
    assign helloWorld_288 = 8'h6E;
    assign helloWorld_289 = 8'h67;
    assign helloWorld_29 = 8'h57;
    assign helloWorld_290 = 8'h20;
    assign helloWorld_291 = 8'h74;
    assign helloWorld_292 = 8'h6F;
    assign helloWorld_293 = 8'h20;
    assign helloWorld_294 = 8'h61;
    assign helloWorld_295 = 8'h63;
    assign helloWorld_296 = 8'h63;
    assign helloWorld_297 = 8'h65;
    assign helloWorld_298 = 8'h70;
    assign helloWorld_299 = 8'h74;
    assign helloWorld_3 = 8'h63;
    assign helloWorld_30 = 8'h65;
    assign helloWorld_300 = 8'h2C;
    assign helloWorld_301 = 8'h20;
    assign helloWorld_302 = 8'h6F;
    assign helloWorld_303 = 8'h6E;
    assign helloWorld_304 = 8'h65;
    assign helloWorld_305 = 8'h20;
    assign helloWorld_306 = 8'h77;
    assign helloWorld_307 = 8'h65;
    assign helloWorld_308 = 8'h20;
    assign helloWorld_309 = 8'h61;
    assign helloWorld_31 = 8'h20;
    assign helloWorld_310 = 8'h72;
    assign helloWorld_311 = 8'h65;
    assign helloWorld_312 = 8'h20;
    assign helloWorld_313 = 8'h75;
    assign helloWorld_314 = 8'h6E;
    assign helloWorld_315 = 8'h77;
    assign helloWorld_316 = 8'h69;
    assign helloWorld_317 = 8'h6C;
    assign helloWorld_318 = 8'h6C;
    assign helloWorld_319 = 8'h69;
    assign helloWorld_32 = 8'h63;
    assign helloWorld_320 = 8'h6E;
    assign helloWorld_321 = 8'h67;
    assign helloWorld_322 = 8'h20;
    assign helloWorld_323 = 8'h74;
    assign helloWorld_324 = 8'h6F;
    assign helloWorld_325 = 8'h20;
    assign helloWorld_326 = 8'h70;
    assign helloWorld_327 = 8'h6F;
    assign helloWorld_328 = 8'h73;
    assign helloWorld_329 = 8'h74;
    assign helloWorld_33 = 8'h68;
    assign helloWorld_330 = 8'h70;
    assign helloWorld_331 = 8'h6F;
    assign helloWorld_332 = 8'h6E;
    assign helloWorld_333 = 8'h65;
    assign helloWorld_334 = 8'h2C;
    assign helloWorld_335 = 8'h20;
    assign helloWorld_336 = 8'h61;
    assign helloWorld_337 = 8'h6E;
    assign helloWorld_338 = 8'h64;
    assign helloWorld_339 = 8'h20;
    assign helloWorld_34 = 8'h6F;
    assign helloWorld_340 = 8'h6F;
    assign helloWorld_341 = 8'h6E;
    assign helloWorld_342 = 8'h65;
    assign helloWorld_343 = 8'h20;
    assign helloWorld_344 = 8'h77;
    assign helloWorld_345 = 8'h68;
    assign helloWorld_346 = 8'h69;
    assign helloWorld_347 = 8'h63;
    assign helloWorld_348 = 8'h68;
    assign helloWorld_349 = 8'h20;
    assign helloWorld_35 = 8'h6F;
    assign helloWorld_350 = 8'h77;
    assign helloWorld_351 = 8'h65;
    assign helloWorld_352 = 8'h20;
    assign helloWorld_353 = 8'h69;
    assign helloWorld_354 = 8'h6E;
    assign helloWorld_355 = 8'h74;
    assign helloWorld_356 = 8'h65;
    assign helloWorld_357 = 8'h6E;
    assign helloWorld_358 = 8'h64;
    assign helloWorld_359 = 8'h20;
    assign helloWorld_36 = 8'h73;
    assign helloWorld_360 = 8'h74;
    assign helloWorld_361 = 8'h6F;
    assign helloWorld_362 = 8'h20;
    assign helloWorld_363 = 8'h77;
    assign helloWorld_364 = 8'h69;
    assign helloWorld_365 = 8'h6E;
    assign helloWorld_366 = 8'h2C;
    assign helloWorld_367 = 8'h20;
    assign helloWorld_368 = 8'h61;
    assign helloWorld_369 = 8'h6E;
    assign helloWorld_37 = 8'h65;
    assign helloWorld_370 = 8'h64;
    assign helloWorld_371 = 8'h20;
    assign helloWorld_372 = 8'h74;
    assign helloWorld_373 = 8'h68;
    assign helloWorld_374 = 8'h65;
    assign helloWorld_375 = 8'h20;
    assign helloWorld_376 = 8'h6F;
    assign helloWorld_377 = 8'h74;
    assign helloWorld_378 = 8'h68;
    assign helloWorld_379 = 8'h65;
    assign helloWorld_38 = 8'h20;
    assign helloWorld_380 = 8'h72;
    assign helloWorld_381 = 8'h73;
    assign helloWorld_382 = 8'h2C;
    assign helloWorld_383 = 8'h20;
    assign helloWorld_384 = 8'h74;
    assign helloWorld_385 = 8'h6F;
    assign helloWorld_386 = 8'h6F;
    assign helloWorld_387 = 8'h2E;
    assign helloWorld_39 = 8'h74;
    assign helloWorld_4 = 8'h68;
    assign helloWorld_40 = 8'h6F;
    assign helloWorld_41 = 8'h20;
    assign helloWorld_42 = 8'h67;
    assign helloWorld_43 = 8'h6F;
    assign helloWorld_44 = 8'h20;
    assign helloWorld_45 = 8'h74;
    assign helloWorld_46 = 8'h6F;
    assign helloWorld_47 = 8'h20;
    assign helloWorld_48 = 8'h74;
    assign helloWorld_49 = 8'h68;
    assign helloWorld_5 = 8'h6F;
    assign helloWorld_50 = 8'h65;
    assign helloWorld_51 = 8'h20;
    assign helloWorld_52 = 8'h6D;
    assign helloWorld_53 = 8'h6F;
    assign helloWorld_54 = 8'h6F;
    assign helloWorld_55 = 8'h6E;
    assign helloWorld_56 = 8'h20;
    assign helloWorld_57 = 8'h69;
    assign helloWorld_58 = 8'h6E;
    assign helloWorld_59 = 8'h20;
    assign helloWorld_6 = 8'h6F;
    assign helloWorld_60 = 8'h74;
    assign helloWorld_61 = 8'h68;
    assign helloWorld_62 = 8'h69;
    assign helloWorld_63 = 8'h73;
    assign helloWorld_64 = 8'h20;
    assign helloWorld_65 = 8'h64;
    assign helloWorld_66 = 8'h65;
    assign helloWorld_67 = 8'h63;
    assign helloWorld_68 = 8'h61;
    assign helloWorld_69 = 8'h64;
    assign helloWorld_7 = 8'h73;
    assign helloWorld_70 = 8'h65;
    assign helloWorld_71 = 8'h20;
    assign helloWorld_72 = 8'h61;
    assign helloWorld_73 = 8'h6E;
    assign helloWorld_74 = 8'h64;
    assign helloWorld_75 = 8'h20;
    assign helloWorld_76 = 8'h64;
    assign helloWorld_77 = 8'h6F;
    assign helloWorld_78 = 8'h20;
    assign helloWorld_79 = 8'h74;
    assign helloWorld_8 = 8'h65;
    assign helloWorld_80 = 8'h68;
    assign helloWorld_81 = 8'h65;
    assign helloWorld_82 = 8'h20;
    assign helloWorld_83 = 8'h6F;
    assign helloWorld_84 = 8'h74;
    assign helloWorld_85 = 8'h68;
    assign helloWorld_86 = 8'h65;
    assign helloWorld_87 = 8'h72;
    assign helloWorld_88 = 8'h20;
    assign helloWorld_89 = 8'h74;
    assign helloWorld_9 = 8'h20;
    assign helloWorld_90 = 8'h68;
    assign helloWorld_91 = 8'h69;
    assign helloWorld_92 = 8'h6E;
    assign helloWorld_93 = 8'h67;
    assign helloWorld_94 = 8'h73;
    assign helloWorld_95 = 8'h2C;
    assign helloWorld_96 = 8'h20;
    assign helloWorld_97 = 8'h6E;
    assign helloWorld_98 = 8'h6F;
    assign helloWorld_99 = 8'h74;
    assign io_character = _GEN_0;
    PAD_UNSIGNED #(.width(1), .n(8)) u_pad_1431 (
        .y(io_characterAvailable),
        .in(_characterArrived__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_1432 (
        .y(_lastToggle__d),
        .sel(reset),
        .a(1'h0),
        .b(_GEN_1)
    );
    MUX_UNSIGNED #(.width(9)) u_mux_1433 (
        .y(_pointer__d),
        .sel(reset),
        .a(9'h0),
        .b(_GEN_3)
    );
endmodule //Console
module DFF_POSCLK(q, d, clk);
    parameter width = 4;
    output reg [width-1:0] q;
    input [width-1:0] d;
    input clk;
    always @(posedge clk) begin
        q <= d;
    end
endmodule // DFF_POSCLK
module NEQ_UNSIGNED(y, a, b);
    parameter width = 4;
    output y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a != b;
endmodule // NEQ_UNSIGNED
module EQ_UNSIGNED(y, a, b);
    parameter width = 4;
    output y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a == b;
endmodule // EQ_UNSIGNED
module PAD_UNSIGNED(y, in);
    parameter width = 4;
    parameter n = 4;
    output [(n > width ? n : width)-1:0] y;
    input [width-1:0] in;
    assign y = (n > width) ? {{(n - width){1'b0}}, in} : in;
endmodule // PAD_UNSIGNED
module ADD_UNSIGNED(y, a, b);
    parameter width = 4;
    output [width:0] y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a + b;
endmodule // ADD_UNSIGNED
module TAIL(y, in);
    parameter width = 4;
    parameter n = 2;
    output [width-n-1:0] y;
    input [width-1:0] in;
    assign y = in[width-n-1:0];
endmodule // TAIL
module MUX_UNSIGNED(y, sel, a, b);
    parameter width = 4;
    output [width-1:0] y;
    input sel;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = sel ? a : b;
endmodule // MUX_UNSIGNED
module BITWISEAND(y, a, b);
    parameter width = 4;
    output [width-1:0] y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a & b;
endmodule // BITWISEAND
