module AdderExerciser(
    input clock,
    input reset
);
    wire [31:0] _ticker__q;
    wire [31:0] _ticker__d;
    DFF_POSCLK #(.width(32)) ticker (
        .q(_ticker__q),
        .d(_ticker__d),
        .clk(clock)
    );
    wire [31:0] _WTEMP_0;
    MUX_UNSIGNED #(.width(32)) u_mux_1 (
        .y(_ticker__d),
        .sel(reset),
        .a(32'h0),
        .b(_WTEMP_0)
    );
    wire [31:0] _max_ticks_for_state__q;
    wire [31:0] _max_ticks_for_state__d;
    DFF_POSCLK #(.width(32)) max_ticks_for_state (
        .q(_max_ticks_for_state__q),
        .d(_max_ticks_for_state__d),
        .clk(clock)
    );
    wire [31:0] _WTEMP_1;
    MUX_UNSIGNED #(.width(32)) u_mux_2 (
        .y(_max_ticks_for_state__d),
        .sel(reset),
        .a(32'h0),
        .b(_WTEMP_1)
    );
    wire [31:0] _state_number__q;
    wire [31:0] _state_number__d;
    DFF_POSCLK #(.width(32)) state_number (
        .q(_state_number__q),
        .d(_state_number__d),
        .clk(clock)
    );
    wire [31:0] _WTEMP_2;
    MUX_UNSIGNED #(.width(32)) u_mux_3 (
        .y(_state_number__d),
        .sel(reset),
        .a(32'h0),
        .b(_WTEMP_2)
    );
    wire _state_locked__q;
    wire _state_locked__d;
    DFF_POSCLK #(.width(1)) state_locked (
        .q(_state_locked__q),
        .d(_state_locked__d),
        .clk(clock)
    );
    wire _WTEMP_3;
    MUX_UNSIGNED #(.width(1)) u_mux_4 (
        .y(_state_locked__d),
        .sel(reset),
        .a(1'h1),
        .b(_WTEMP_3)
    );
    wire [32:0] _T_11;
    wire [31:0] _WTEMP_4;
    PAD_UNSIGNED #(.width(1), .n(32)) u_pad_5 (
        .y(_WTEMP_4),
        .in(1'h1)
    );
    ADD_UNSIGNED #(.width(32)) u_add_6 (
        .y(_T_11),
        .a(_ticker__q),
        .b(_WTEMP_4)
    );
    wire [31:0] _T_12;
    TAIL #(.width(33), .n(1)) tail_7 (
        .y(_T_12),
        .in(_T_11)
    );
    wire _T_14;
    EQ_UNSIGNED #(.width(1)) u_eq_8 (
        .y(_T_14),
        .a(_state_locked__q),
        .b(1'h0)
    );
    wire [32:0] _T_17;
    wire [31:0] _WTEMP_5;
    PAD_UNSIGNED #(.width(1), .n(32)) u_pad_9 (
        .y(_WTEMP_5),
        .in(1'h1)
    );
    ADD_UNSIGNED #(.width(32)) u_add_10 (
        .y(_T_17),
        .a(_state_number__q),
        .b(_WTEMP_5)
    );
    wire [31:0] _T_18;
    TAIL #(.width(33), .n(1)) tail_11 (
        .y(_T_18),
        .in(_T_17)
    );
    wire _T_19;
    GT_UNSIGNED #(.width(32)) u_gt_12 (
        .y(_T_19),
        .a(_ticker__q),
        .b(_max_ticks_for_state__q)
    );
    wire _T_21;
    EQ_UNSIGNED #(.width(1)) u_eq_13 (
        .y(_T_21),
        .a(_T_14),
        .b(1'h0)
    );
    wire _T_22;
    BITWISEAND #(.width(1)) bitwiseand_14 (
        .y(_T_22),
        .a(_T_21),
        .b(_T_19)
    );
    wire _T_24;
    EQ_UNSIGNED #(.width(1)) u_eq_15 (
        .y(_T_24),
        .a(reset),
        .b(1'h0)
    );
    wire [32:0] _T_27;
    wire [31:0] _WTEMP_6;
    PAD_UNSIGNED #(.width(1), .n(32)) u_pad_16 (
        .y(_WTEMP_6),
        .in(1'h1)
    );
    ADD_UNSIGNED #(.width(32)) u_add_17 (
        .y(_T_27),
        .a(_state_number__q),
        .b(_WTEMP_6)
    );
    wire [31:0] _T_28;
    TAIL #(.width(33), .n(1)) tail_18 (
        .y(_T_28),
        .in(_T_27)
    );
    wire [31:0] _node_0;
    MUX_UNSIGNED #(.width(32)) u_mux_19 (
        .y(_node_0),
        .sel(_T_14),
        .a(_T_18),
        .b(_state_number__q)
    );
    wire _T_30;
    wire [31:0] _WTEMP_7;
    PAD_UNSIGNED #(.width(7), .n(32)) u_pad_20 (
        .y(_WTEMP_7),
        .in(7'h64)
    );
    GT_UNSIGNED #(.width(32)) u_gt_21 (
        .y(_T_30),
        .a(_ticker__q),
        .b(_WTEMP_7)
    );
    wire _T_32;
    EQ_UNSIGNED #(.width(1)) u_eq_22 (
        .y(_T_32),
        .a(reset),
        .b(1'h0)
    );
    wire _T_34;
    EQ_UNSIGNED #(.width(1)) u_eq_23 (
        .y(_T_34),
        .a(reset),
        .b(1'h0)
    );
    wire _c__clock;
    wire _c__reset;
    wire [31:0] _c__io_in0;
    wire [31:0] _c__io_in1;
    wire [31:0] _c__io_out;
    Adder c (
        .clock(_c__clock),
        .reset(_c__reset),
        .io_in0(_c__io_in0),
        .io_in1(_c__io_in1),
        .io_out(_c__io_out)
    );
    wire _T_36;
    EQ_UNSIGNED #(.width(1)) u_eq_26 (
        .y(_T_36),
        .a(reset),
        .b(1'h0)
    );
    wire [4:0] in0_vec_0;
    wire [4:0] in0_vec_1;
    wire [4:0] in0_vec_2;
    wire [4:0] in0_vec_3;
    wire [4:0] in0_vec_4;
    wire [4:0] in0_vec_5;
    wire [4:0] in0_vec_6;
    wire [4:0] in0_vec_7;
    wire [4:0] in0_vec_8;
    wire [4:0] in0_vec_9;
    wire [4:0] in0_vec_10;
    wire [4:0] in0_vec_11;
    wire [4:0] in0_vec_12;
    wire [4:0] in0_vec_13;
    wire [4:0] in0_vec_14;
    wire [4:0] in0_vec_15;
    wire [4:0] in0_vec_16;
    wire [4:0] in0_vec_17;
    wire [4:0] in0_vec_18;
    wire [4:0] in0_vec_19;
    wire [4:0] in1_vec_0;
    wire [4:0] in1_vec_1;
    wire [4:0] in1_vec_2;
    wire [4:0] in1_vec_3;
    wire [4:0] in1_vec_4;
    wire [4:0] in1_vec_5;
    wire [4:0] in1_vec_6;
    wire [4:0] in1_vec_7;
    wire [4:0] in1_vec_8;
    wire [4:0] in1_vec_9;
    wire [4:0] in1_vec_10;
    wire [4:0] in1_vec_11;
    wire [4:0] in1_vec_12;
    wire [4:0] in1_vec_13;
    wire [4:0] in1_vec_14;
    wire [4:0] in1_vec_15;
    wire [4:0] in1_vec_16;
    wire [4:0] in1_vec_17;
    wire [4:0] in1_vec_18;
    wire [4:0] in1_vec_19;
    wire [5:0] _T_125;
    ADD_UNSIGNED #(.width(5)) u_add_27 (
        .y(_T_125),
        .a(in0_vec_0),
        .b(in1_vec_0)
    );
    wire [4:0] _T_126;
    TAIL #(.width(6), .n(1)) tail_28 (
        .y(_T_126),
        .in(_T_125)
    );
    wire [5:0] _T_127;
    ADD_UNSIGNED #(.width(5)) u_add_29 (
        .y(_T_127),
        .a(in0_vec_1),
        .b(in1_vec_1)
    );
    wire [4:0] _T_128;
    TAIL #(.width(6), .n(1)) tail_30 (
        .y(_T_128),
        .in(_T_127)
    );
    wire [5:0] _T_129;
    ADD_UNSIGNED #(.width(5)) u_add_31 (
        .y(_T_129),
        .a(in0_vec_2),
        .b(in1_vec_2)
    );
    wire [4:0] _T_130;
    TAIL #(.width(6), .n(1)) tail_32 (
        .y(_T_130),
        .in(_T_129)
    );
    wire [5:0] _T_131;
    ADD_UNSIGNED #(.width(5)) u_add_33 (
        .y(_T_131),
        .a(in0_vec_3),
        .b(in1_vec_3)
    );
    wire [4:0] _T_132;
    TAIL #(.width(6), .n(1)) tail_34 (
        .y(_T_132),
        .in(_T_131)
    );
    wire [5:0] _T_133;
    ADD_UNSIGNED #(.width(5)) u_add_35 (
        .y(_T_133),
        .a(in0_vec_4),
        .b(in1_vec_4)
    );
    wire [4:0] _T_134;
    TAIL #(.width(6), .n(1)) tail_36 (
        .y(_T_134),
        .in(_T_133)
    );
    wire [5:0] _T_135;
    ADD_UNSIGNED #(.width(5)) u_add_37 (
        .y(_T_135),
        .a(in0_vec_5),
        .b(in1_vec_5)
    );
    wire [4:0] _T_136;
    TAIL #(.width(6), .n(1)) tail_38 (
        .y(_T_136),
        .in(_T_135)
    );
    wire [5:0] _T_137;
    ADD_UNSIGNED #(.width(5)) u_add_39 (
        .y(_T_137),
        .a(in0_vec_6),
        .b(in1_vec_6)
    );
    wire [4:0] _T_138;
    TAIL #(.width(6), .n(1)) tail_40 (
        .y(_T_138),
        .in(_T_137)
    );
    wire [5:0] _T_139;
    ADD_UNSIGNED #(.width(5)) u_add_41 (
        .y(_T_139),
        .a(in0_vec_7),
        .b(in1_vec_7)
    );
    wire [4:0] _T_140;
    TAIL #(.width(6), .n(1)) tail_42 (
        .y(_T_140),
        .in(_T_139)
    );
    wire [5:0] _T_141;
    ADD_UNSIGNED #(.width(5)) u_add_43 (
        .y(_T_141),
        .a(in0_vec_8),
        .b(in1_vec_8)
    );
    wire [4:0] _T_142;
    TAIL #(.width(6), .n(1)) tail_44 (
        .y(_T_142),
        .in(_T_141)
    );
    wire [5:0] _T_143;
    ADD_UNSIGNED #(.width(5)) u_add_45 (
        .y(_T_143),
        .a(in0_vec_9),
        .b(in1_vec_9)
    );
    wire [4:0] _T_144;
    TAIL #(.width(6), .n(1)) tail_46 (
        .y(_T_144),
        .in(_T_143)
    );
    wire [5:0] _T_145;
    ADD_UNSIGNED #(.width(5)) u_add_47 (
        .y(_T_145),
        .a(in0_vec_10),
        .b(in1_vec_10)
    );
    wire [4:0] _T_146;
    TAIL #(.width(6), .n(1)) tail_48 (
        .y(_T_146),
        .in(_T_145)
    );
    wire [5:0] _T_147;
    ADD_UNSIGNED #(.width(5)) u_add_49 (
        .y(_T_147),
        .a(in0_vec_11),
        .b(in1_vec_11)
    );
    wire [4:0] _T_148;
    TAIL #(.width(6), .n(1)) tail_50 (
        .y(_T_148),
        .in(_T_147)
    );
    wire [5:0] _T_149;
    ADD_UNSIGNED #(.width(5)) u_add_51 (
        .y(_T_149),
        .a(in0_vec_12),
        .b(in1_vec_12)
    );
    wire [4:0] _T_150;
    TAIL #(.width(6), .n(1)) tail_52 (
        .y(_T_150),
        .in(_T_149)
    );
    wire [5:0] _T_151;
    ADD_UNSIGNED #(.width(5)) u_add_53 (
        .y(_T_151),
        .a(in0_vec_13),
        .b(in1_vec_13)
    );
    wire [4:0] _T_152;
    TAIL #(.width(6), .n(1)) tail_54 (
        .y(_T_152),
        .in(_T_151)
    );
    wire [5:0] _T_153;
    ADD_UNSIGNED #(.width(5)) u_add_55 (
        .y(_T_153),
        .a(in0_vec_14),
        .b(in1_vec_14)
    );
    wire [4:0] _T_154;
    TAIL #(.width(6), .n(1)) tail_56 (
        .y(_T_154),
        .in(_T_153)
    );
    wire [5:0] _T_155;
    ADD_UNSIGNED #(.width(5)) u_add_57 (
        .y(_T_155),
        .a(in0_vec_15),
        .b(in1_vec_15)
    );
    wire [4:0] _T_156;
    TAIL #(.width(6), .n(1)) tail_58 (
        .y(_T_156),
        .in(_T_155)
    );
    wire [5:0] _T_157;
    ADD_UNSIGNED #(.width(5)) u_add_59 (
        .y(_T_157),
        .a(in0_vec_16),
        .b(in1_vec_16)
    );
    wire [4:0] _T_158;
    TAIL #(.width(6), .n(1)) tail_60 (
        .y(_T_158),
        .in(_T_157)
    );
    wire [5:0] _T_159;
    ADD_UNSIGNED #(.width(5)) u_add_61 (
        .y(_T_159),
        .a(in0_vec_17),
        .b(in1_vec_17)
    );
    wire [4:0] _T_160;
    TAIL #(.width(6), .n(1)) tail_62 (
        .y(_T_160),
        .in(_T_159)
    );
    wire [5:0] _T_161;
    ADD_UNSIGNED #(.width(5)) u_add_63 (
        .y(_T_161),
        .a(in0_vec_18),
        .b(in1_vec_18)
    );
    wire [4:0] _T_162;
    TAIL #(.width(6), .n(1)) tail_64 (
        .y(_T_162),
        .in(_T_161)
    );
    wire [5:0] _T_163;
    ADD_UNSIGNED #(.width(5)) u_add_65 (
        .y(_T_163),
        .a(in0_vec_19),
        .b(in1_vec_19)
    );
    wire [4:0] _T_164;
    TAIL #(.width(6), .n(1)) tail_66 (
        .y(_T_164),
        .in(_T_163)
    );
    wire [4:0] expected_out_vec_0;
    wire [4:0] expected_out_vec_1;
    wire [4:0] expected_out_vec_2;
    wire [4:0] expected_out_vec_3;
    wire [4:0] expected_out_vec_4;
    wire [4:0] expected_out_vec_5;
    wire [4:0] expected_out_vec_6;
    wire [4:0] expected_out_vec_7;
    wire [4:0] expected_out_vec_8;
    wire [4:0] expected_out_vec_9;
    wire [4:0] expected_out_vec_10;
    wire [4:0] expected_out_vec_11;
    wire [4:0] expected_out_vec_12;
    wire [4:0] expected_out_vec_13;
    wire [4:0] expected_out_vec_14;
    wire [4:0] expected_out_vec_15;
    wire [4:0] expected_out_vec_16;
    wire [4:0] expected_out_vec_17;
    wire [4:0] expected_out_vec_18;
    wire [4:0] expected_out_vec_19;
    wire [31:0] _test_number__q;
    wire [31:0] _test_number__d;
    DFF_POSCLK #(.width(32)) test_number (
        .q(_test_number__q),
        .d(_test_number__d),
        .clk(clock)
    );
    wire [31:0] _WTEMP_8;
    MUX_UNSIGNED #(.width(32)) u_mux_67 (
        .y(_test_number__d),
        .sel(reset),
        .a(32'h0),
        .b(_WTEMP_8)
    );
    wire _T_192;
    wire [31:0] _WTEMP_9;
    PAD_UNSIGNED #(.width(5), .n(32)) u_pad_68 (
        .y(_WTEMP_9),
        .in(5'h14)
    );
    GT_UNSIGNED #(.width(32)) u_gt_69 (
        .y(_T_192),
        .a(_test_number__q),
        .b(_WTEMP_9)
    );
    wire _T_194;
    wire [31:0] _WTEMP_10;
    PAD_UNSIGNED #(.width(6), .n(32)) u_pad_70 (
        .y(_WTEMP_10),
        .in(6'h21)
    );
    EQ_UNSIGNED #(.width(32)) u_eq_71 (
        .y(_T_194),
        .a(_state_number__q),
        .b(_WTEMP_10)
    );
    wire _T_196;
    EQ_UNSIGNED #(.width(1)) u_eq_72 (
        .y(_T_196),
        .a(_state_locked__q),
        .b(1'h0)
    );
    wire _T_198;
    EQ_UNSIGNED #(.width(1)) u_eq_73 (
        .y(_T_198),
        .a(reset),
        .b(1'h0)
    );
    wire _node_1;
    MUX_UNSIGNED #(.width(1)) u_mux_74 (
        .y(_node_1),
        .sel(_T_22),
        .a(1'h0),
        .b(_state_locked__q)
    );
    wire [31:0] _node_2;
    MUX_UNSIGNED #(.width(32)) u_mux_75 (
        .y(_node_2),
        .sel(_T_22),
        .a(_T_28),
        .b(_node_0)
    );
    wire [31:0] _node_3;
    wire [31:0] _WTEMP_11;
    PAD_UNSIGNED #(.width(1), .n(32)) u_pad_76 (
        .y(_WTEMP_11),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(32)) u_mux_77 (
        .y(_node_3),
        .sel(_T_14),
        .a(_WTEMP_11),
        .b(_T_12)
    );
    wire [4:0] _T_204;
    BITS #(.width(32), .high(4), .low(0)) bits_78 (
        .y(_T_204),
        .in(_test_number__q)
    );
    wire [4:0] _T_206;
    BITS #(.width(32), .high(4), .low(0)) bits_79 (
        .y(_T_206),
        .in(_test_number__q)
    );
    wire [4:0] _T_208;
    BITS #(.width(32), .high(4), .low(0)) bits_80 (
        .y(_T_208),
        .in(_test_number__q)
    );
    wire [4:0] _T_210;
    BITS #(.width(32), .high(4), .low(0)) bits_81 (
        .y(_T_210),
        .in(_test_number__q)
    );
    wire _node_4;
    EQ_UNSIGNED #(.width(5)) u_eq_82 (
        .y(_node_4),
        .a(5'd0),
        .b(_T_208)
    );
    wire [4:0] _node_5;
    assign _node_5 = in0_vec_0;
    wire _node_6;
    EQ_UNSIGNED #(.width(5)) u_eq_83 (
        .y(_node_6),
        .a(5'd1),
        .b(_T_208)
    );
    wire [4:0] _node_7;
    MUX_UNSIGNED #(.width(5)) u_mux_84 (
        .y(_node_7),
        .sel(_node_6),
        .a(in0_vec_1),
        .b(_node_5)
    );
    wire _node_8;
    EQ_UNSIGNED #(.width(5)) u_eq_85 (
        .y(_node_8),
        .a(5'd2),
        .b(_T_208)
    );
    wire [4:0] _node_9;
    MUX_UNSIGNED #(.width(5)) u_mux_86 (
        .y(_node_9),
        .sel(_node_8),
        .a(in0_vec_2),
        .b(_node_7)
    );
    wire _node_10;
    EQ_UNSIGNED #(.width(5)) u_eq_87 (
        .y(_node_10),
        .a(5'd3),
        .b(_T_208)
    );
    wire [4:0] _node_11;
    MUX_UNSIGNED #(.width(5)) u_mux_88 (
        .y(_node_11),
        .sel(_node_10),
        .a(in0_vec_3),
        .b(_node_9)
    );
    wire _node_12;
    EQ_UNSIGNED #(.width(5)) u_eq_89 (
        .y(_node_12),
        .a(5'd4),
        .b(_T_208)
    );
    wire [4:0] _node_13;
    MUX_UNSIGNED #(.width(5)) u_mux_90 (
        .y(_node_13),
        .sel(_node_12),
        .a(in0_vec_4),
        .b(_node_11)
    );
    wire _node_14;
    EQ_UNSIGNED #(.width(5)) u_eq_91 (
        .y(_node_14),
        .a(5'd5),
        .b(_T_208)
    );
    wire [4:0] _node_15;
    MUX_UNSIGNED #(.width(5)) u_mux_92 (
        .y(_node_15),
        .sel(_node_14),
        .a(in0_vec_5),
        .b(_node_13)
    );
    wire _node_16;
    EQ_UNSIGNED #(.width(5)) u_eq_93 (
        .y(_node_16),
        .a(5'd6),
        .b(_T_208)
    );
    wire [4:0] _node_17;
    MUX_UNSIGNED #(.width(5)) u_mux_94 (
        .y(_node_17),
        .sel(_node_16),
        .a(in0_vec_6),
        .b(_node_15)
    );
    wire _node_18;
    EQ_UNSIGNED #(.width(5)) u_eq_95 (
        .y(_node_18),
        .a(5'd7),
        .b(_T_208)
    );
    wire [4:0] _node_19;
    MUX_UNSIGNED #(.width(5)) u_mux_96 (
        .y(_node_19),
        .sel(_node_18),
        .a(in0_vec_7),
        .b(_node_17)
    );
    wire _node_20;
    EQ_UNSIGNED #(.width(5)) u_eq_97 (
        .y(_node_20),
        .a(5'd8),
        .b(_T_208)
    );
    wire [4:0] _node_21;
    MUX_UNSIGNED #(.width(5)) u_mux_98 (
        .y(_node_21),
        .sel(_node_20),
        .a(in0_vec_8),
        .b(_node_19)
    );
    wire _node_22;
    EQ_UNSIGNED #(.width(5)) u_eq_99 (
        .y(_node_22),
        .a(5'd9),
        .b(_T_208)
    );
    wire [4:0] _node_23;
    MUX_UNSIGNED #(.width(5)) u_mux_100 (
        .y(_node_23),
        .sel(_node_22),
        .a(in0_vec_9),
        .b(_node_21)
    );
    wire _node_24;
    EQ_UNSIGNED #(.width(5)) u_eq_101 (
        .y(_node_24),
        .a(5'd10),
        .b(_T_208)
    );
    wire [4:0] _node_25;
    MUX_UNSIGNED #(.width(5)) u_mux_102 (
        .y(_node_25),
        .sel(_node_24),
        .a(in0_vec_10),
        .b(_node_23)
    );
    wire _node_26;
    EQ_UNSIGNED #(.width(5)) u_eq_103 (
        .y(_node_26),
        .a(5'd11),
        .b(_T_208)
    );
    wire [4:0] _node_27;
    MUX_UNSIGNED #(.width(5)) u_mux_104 (
        .y(_node_27),
        .sel(_node_26),
        .a(in0_vec_11),
        .b(_node_25)
    );
    wire _node_28;
    EQ_UNSIGNED #(.width(5)) u_eq_105 (
        .y(_node_28),
        .a(5'd12),
        .b(_T_208)
    );
    wire [4:0] _node_29;
    MUX_UNSIGNED #(.width(5)) u_mux_106 (
        .y(_node_29),
        .sel(_node_28),
        .a(in0_vec_12),
        .b(_node_27)
    );
    wire _node_30;
    EQ_UNSIGNED #(.width(5)) u_eq_107 (
        .y(_node_30),
        .a(5'd13),
        .b(_T_208)
    );
    wire [4:0] _node_31;
    MUX_UNSIGNED #(.width(5)) u_mux_108 (
        .y(_node_31),
        .sel(_node_30),
        .a(in0_vec_13),
        .b(_node_29)
    );
    wire _node_32;
    EQ_UNSIGNED #(.width(5)) u_eq_109 (
        .y(_node_32),
        .a(5'd14),
        .b(_T_208)
    );
    wire [4:0] _node_33;
    MUX_UNSIGNED #(.width(5)) u_mux_110 (
        .y(_node_33),
        .sel(_node_32),
        .a(in0_vec_14),
        .b(_node_31)
    );
    wire _node_34;
    EQ_UNSIGNED #(.width(5)) u_eq_111 (
        .y(_node_34),
        .a(5'd15),
        .b(_T_208)
    );
    wire [4:0] _node_35;
    MUX_UNSIGNED #(.width(5)) u_mux_112 (
        .y(_node_35),
        .sel(_node_34),
        .a(in0_vec_15),
        .b(_node_33)
    );
    wire _node_36;
    EQ_UNSIGNED #(.width(5)) u_eq_113 (
        .y(_node_36),
        .a(5'd16),
        .b(_T_208)
    );
    wire [4:0] _node_37;
    MUX_UNSIGNED #(.width(5)) u_mux_114 (
        .y(_node_37),
        .sel(_node_36),
        .a(in0_vec_16),
        .b(_node_35)
    );
    wire _node_38;
    EQ_UNSIGNED #(.width(5)) u_eq_115 (
        .y(_node_38),
        .a(5'd17),
        .b(_T_208)
    );
    wire [4:0] _node_39;
    MUX_UNSIGNED #(.width(5)) u_mux_116 (
        .y(_node_39),
        .sel(_node_38),
        .a(in0_vec_17),
        .b(_node_37)
    );
    wire _node_40;
    EQ_UNSIGNED #(.width(5)) u_eq_117 (
        .y(_node_40),
        .a(5'd18),
        .b(_T_208)
    );
    wire [4:0] _node_41;
    MUX_UNSIGNED #(.width(5)) u_mux_118 (
        .y(_node_41),
        .sel(_node_40),
        .a(in0_vec_18),
        .b(_node_39)
    );
    wire _node_42;
    EQ_UNSIGNED #(.width(5)) u_eq_119 (
        .y(_node_42),
        .a(5'd19),
        .b(_T_208)
    );
    wire [4:0] _node_43;
    MUX_UNSIGNED #(.width(5)) u_mux_120 (
        .y(_node_43),
        .sel(_node_42),
        .a(in0_vec_19),
        .b(_node_41)
    );
    wire _node_44;
    EQ_UNSIGNED #(.width(5)) u_eq_121 (
        .y(_node_44),
        .a(5'd0),
        .b(_T_210)
    );
    wire [4:0] _node_45;
    assign _node_45 = in1_vec_0;
    wire _node_46;
    EQ_UNSIGNED #(.width(5)) u_eq_122 (
        .y(_node_46),
        .a(5'd1),
        .b(_T_210)
    );
    wire [4:0] _node_47;
    MUX_UNSIGNED #(.width(5)) u_mux_123 (
        .y(_node_47),
        .sel(_node_46),
        .a(in1_vec_1),
        .b(_node_45)
    );
    wire _node_48;
    EQ_UNSIGNED #(.width(5)) u_eq_124 (
        .y(_node_48),
        .a(5'd2),
        .b(_T_210)
    );
    wire [4:0] _node_49;
    MUX_UNSIGNED #(.width(5)) u_mux_125 (
        .y(_node_49),
        .sel(_node_48),
        .a(in1_vec_2),
        .b(_node_47)
    );
    wire _node_50;
    EQ_UNSIGNED #(.width(5)) u_eq_126 (
        .y(_node_50),
        .a(5'd3),
        .b(_T_210)
    );
    wire [4:0] _node_51;
    MUX_UNSIGNED #(.width(5)) u_mux_127 (
        .y(_node_51),
        .sel(_node_50),
        .a(in1_vec_3),
        .b(_node_49)
    );
    wire _node_52;
    EQ_UNSIGNED #(.width(5)) u_eq_128 (
        .y(_node_52),
        .a(5'd4),
        .b(_T_210)
    );
    wire [4:0] _node_53;
    MUX_UNSIGNED #(.width(5)) u_mux_129 (
        .y(_node_53),
        .sel(_node_52),
        .a(in1_vec_4),
        .b(_node_51)
    );
    wire _node_54;
    EQ_UNSIGNED #(.width(5)) u_eq_130 (
        .y(_node_54),
        .a(5'd5),
        .b(_T_210)
    );
    wire [4:0] _node_55;
    MUX_UNSIGNED #(.width(5)) u_mux_131 (
        .y(_node_55),
        .sel(_node_54),
        .a(in1_vec_5),
        .b(_node_53)
    );
    wire _node_56;
    EQ_UNSIGNED #(.width(5)) u_eq_132 (
        .y(_node_56),
        .a(5'd6),
        .b(_T_210)
    );
    wire [4:0] _node_57;
    MUX_UNSIGNED #(.width(5)) u_mux_133 (
        .y(_node_57),
        .sel(_node_56),
        .a(in1_vec_6),
        .b(_node_55)
    );
    wire _node_58;
    EQ_UNSIGNED #(.width(5)) u_eq_134 (
        .y(_node_58),
        .a(5'd7),
        .b(_T_210)
    );
    wire [4:0] _node_59;
    MUX_UNSIGNED #(.width(5)) u_mux_135 (
        .y(_node_59),
        .sel(_node_58),
        .a(in1_vec_7),
        .b(_node_57)
    );
    wire _node_60;
    EQ_UNSIGNED #(.width(5)) u_eq_136 (
        .y(_node_60),
        .a(5'd8),
        .b(_T_210)
    );
    wire [4:0] _node_61;
    MUX_UNSIGNED #(.width(5)) u_mux_137 (
        .y(_node_61),
        .sel(_node_60),
        .a(in1_vec_8),
        .b(_node_59)
    );
    wire _node_62;
    EQ_UNSIGNED #(.width(5)) u_eq_138 (
        .y(_node_62),
        .a(5'd9),
        .b(_T_210)
    );
    wire [4:0] _node_63;
    MUX_UNSIGNED #(.width(5)) u_mux_139 (
        .y(_node_63),
        .sel(_node_62),
        .a(in1_vec_9),
        .b(_node_61)
    );
    wire _node_64;
    EQ_UNSIGNED #(.width(5)) u_eq_140 (
        .y(_node_64),
        .a(5'd10),
        .b(_T_210)
    );
    wire [4:0] _node_65;
    MUX_UNSIGNED #(.width(5)) u_mux_141 (
        .y(_node_65),
        .sel(_node_64),
        .a(in1_vec_10),
        .b(_node_63)
    );
    wire _node_66;
    EQ_UNSIGNED #(.width(5)) u_eq_142 (
        .y(_node_66),
        .a(5'd11),
        .b(_T_210)
    );
    wire [4:0] _node_67;
    MUX_UNSIGNED #(.width(5)) u_mux_143 (
        .y(_node_67),
        .sel(_node_66),
        .a(in1_vec_11),
        .b(_node_65)
    );
    wire _node_68;
    EQ_UNSIGNED #(.width(5)) u_eq_144 (
        .y(_node_68),
        .a(5'd12),
        .b(_T_210)
    );
    wire [4:0] _node_69;
    MUX_UNSIGNED #(.width(5)) u_mux_145 (
        .y(_node_69),
        .sel(_node_68),
        .a(in1_vec_12),
        .b(_node_67)
    );
    wire _node_70;
    EQ_UNSIGNED #(.width(5)) u_eq_146 (
        .y(_node_70),
        .a(5'd13),
        .b(_T_210)
    );
    wire [4:0] _node_71;
    MUX_UNSIGNED #(.width(5)) u_mux_147 (
        .y(_node_71),
        .sel(_node_70),
        .a(in1_vec_13),
        .b(_node_69)
    );
    wire _node_72;
    EQ_UNSIGNED #(.width(5)) u_eq_148 (
        .y(_node_72),
        .a(5'd14),
        .b(_T_210)
    );
    wire [4:0] _node_73;
    MUX_UNSIGNED #(.width(5)) u_mux_149 (
        .y(_node_73),
        .sel(_node_72),
        .a(in1_vec_14),
        .b(_node_71)
    );
    wire _node_74;
    EQ_UNSIGNED #(.width(5)) u_eq_150 (
        .y(_node_74),
        .a(5'd15),
        .b(_T_210)
    );
    wire [4:0] _node_75;
    MUX_UNSIGNED #(.width(5)) u_mux_151 (
        .y(_node_75),
        .sel(_node_74),
        .a(in1_vec_15),
        .b(_node_73)
    );
    wire _node_76;
    EQ_UNSIGNED #(.width(5)) u_eq_152 (
        .y(_node_76),
        .a(5'd16),
        .b(_T_210)
    );
    wire [4:0] _node_77;
    MUX_UNSIGNED #(.width(5)) u_mux_153 (
        .y(_node_77),
        .sel(_node_76),
        .a(in1_vec_16),
        .b(_node_75)
    );
    wire _node_78;
    EQ_UNSIGNED #(.width(5)) u_eq_154 (
        .y(_node_78),
        .a(5'd17),
        .b(_T_210)
    );
    wire [4:0] _node_79;
    MUX_UNSIGNED #(.width(5)) u_mux_155 (
        .y(_node_79),
        .sel(_node_78),
        .a(in1_vec_17),
        .b(_node_77)
    );
    wire _node_80;
    EQ_UNSIGNED #(.width(5)) u_eq_156 (
        .y(_node_80),
        .a(5'd18),
        .b(_T_210)
    );
    wire [4:0] _node_81;
    MUX_UNSIGNED #(.width(5)) u_mux_157 (
        .y(_node_81),
        .sel(_node_80),
        .a(in1_vec_18),
        .b(_node_79)
    );
    wire _node_82;
    EQ_UNSIGNED #(.width(5)) u_eq_158 (
        .y(_node_82),
        .a(5'd19),
        .b(_T_210)
    );
    wire [4:0] _node_83;
    MUX_UNSIGNED #(.width(5)) u_mux_159 (
        .y(_node_83),
        .sel(_node_82),
        .a(in1_vec_19),
        .b(_node_81)
    );
    wire [5:0] _T_211;
    ADD_UNSIGNED #(.width(5)) u_add_160 (
        .y(_T_211),
        .a(_node_43),
        .b(_node_83)
    );
    wire [4:0] _T_212;
    TAIL #(.width(6), .n(1)) tail_161 (
        .y(_T_212),
        .in(_T_211)
    );
    wire [4:0] _T_214;
    BITS #(.width(32), .high(4), .low(0)) bits_162 (
        .y(_T_214),
        .in(_test_number__q)
    );
    wire _T_216;
    EQ_UNSIGNED #(.width(1)) u_eq_163 (
        .y(_T_216),
        .a(reset),
        .b(1'h0)
    );
    wire [4:0] _T_218;
    BITS #(.width(32), .high(4), .low(0)) bits_164 (
        .y(_T_218),
        .in(_test_number__q)
    );
    wire [4:0] _T_220;
    BITS #(.width(32), .high(4), .low(0)) bits_165 (
        .y(_T_220),
        .in(_test_number__q)
    );
    wire [4:0] _T_222;
    BITS #(.width(32), .high(4), .low(0)) bits_166 (
        .y(_T_222),
        .in(_test_number__q)
    );
    wire _node_84;
    EQ_UNSIGNED #(.width(5)) u_eq_167 (
        .y(_node_84),
        .a(5'd0),
        .b(_T_220)
    );
    wire [4:0] _node_85;
    assign _node_85 = in0_vec_0;
    wire _node_86;
    EQ_UNSIGNED #(.width(5)) u_eq_168 (
        .y(_node_86),
        .a(5'd1),
        .b(_T_220)
    );
    wire [4:0] _node_87;
    MUX_UNSIGNED #(.width(5)) u_mux_169 (
        .y(_node_87),
        .sel(_node_86),
        .a(in0_vec_1),
        .b(_node_85)
    );
    wire _node_88;
    EQ_UNSIGNED #(.width(5)) u_eq_170 (
        .y(_node_88),
        .a(5'd2),
        .b(_T_220)
    );
    wire [4:0] _node_89;
    MUX_UNSIGNED #(.width(5)) u_mux_171 (
        .y(_node_89),
        .sel(_node_88),
        .a(in0_vec_2),
        .b(_node_87)
    );
    wire _node_90;
    EQ_UNSIGNED #(.width(5)) u_eq_172 (
        .y(_node_90),
        .a(5'd3),
        .b(_T_220)
    );
    wire [4:0] _node_91;
    MUX_UNSIGNED #(.width(5)) u_mux_173 (
        .y(_node_91),
        .sel(_node_90),
        .a(in0_vec_3),
        .b(_node_89)
    );
    wire _node_92;
    EQ_UNSIGNED #(.width(5)) u_eq_174 (
        .y(_node_92),
        .a(5'd4),
        .b(_T_220)
    );
    wire [4:0] _node_93;
    MUX_UNSIGNED #(.width(5)) u_mux_175 (
        .y(_node_93),
        .sel(_node_92),
        .a(in0_vec_4),
        .b(_node_91)
    );
    wire _node_94;
    EQ_UNSIGNED #(.width(5)) u_eq_176 (
        .y(_node_94),
        .a(5'd5),
        .b(_T_220)
    );
    wire [4:0] _node_95;
    MUX_UNSIGNED #(.width(5)) u_mux_177 (
        .y(_node_95),
        .sel(_node_94),
        .a(in0_vec_5),
        .b(_node_93)
    );
    wire _node_96;
    EQ_UNSIGNED #(.width(5)) u_eq_178 (
        .y(_node_96),
        .a(5'd6),
        .b(_T_220)
    );
    wire [4:0] _node_97;
    MUX_UNSIGNED #(.width(5)) u_mux_179 (
        .y(_node_97),
        .sel(_node_96),
        .a(in0_vec_6),
        .b(_node_95)
    );
    wire _node_98;
    EQ_UNSIGNED #(.width(5)) u_eq_180 (
        .y(_node_98),
        .a(5'd7),
        .b(_T_220)
    );
    wire [4:0] _node_99;
    MUX_UNSIGNED #(.width(5)) u_mux_181 (
        .y(_node_99),
        .sel(_node_98),
        .a(in0_vec_7),
        .b(_node_97)
    );
    wire _node_100;
    EQ_UNSIGNED #(.width(5)) u_eq_182 (
        .y(_node_100),
        .a(5'd8),
        .b(_T_220)
    );
    wire [4:0] _node_101;
    MUX_UNSIGNED #(.width(5)) u_mux_183 (
        .y(_node_101),
        .sel(_node_100),
        .a(in0_vec_8),
        .b(_node_99)
    );
    wire _node_102;
    EQ_UNSIGNED #(.width(5)) u_eq_184 (
        .y(_node_102),
        .a(5'd9),
        .b(_T_220)
    );
    wire [4:0] _node_103;
    MUX_UNSIGNED #(.width(5)) u_mux_185 (
        .y(_node_103),
        .sel(_node_102),
        .a(in0_vec_9),
        .b(_node_101)
    );
    wire _node_104;
    EQ_UNSIGNED #(.width(5)) u_eq_186 (
        .y(_node_104),
        .a(5'd10),
        .b(_T_220)
    );
    wire [4:0] _node_105;
    MUX_UNSIGNED #(.width(5)) u_mux_187 (
        .y(_node_105),
        .sel(_node_104),
        .a(in0_vec_10),
        .b(_node_103)
    );
    wire _node_106;
    EQ_UNSIGNED #(.width(5)) u_eq_188 (
        .y(_node_106),
        .a(5'd11),
        .b(_T_220)
    );
    wire [4:0] _node_107;
    MUX_UNSIGNED #(.width(5)) u_mux_189 (
        .y(_node_107),
        .sel(_node_106),
        .a(in0_vec_11),
        .b(_node_105)
    );
    wire _node_108;
    EQ_UNSIGNED #(.width(5)) u_eq_190 (
        .y(_node_108),
        .a(5'd12),
        .b(_T_220)
    );
    wire [4:0] _node_109;
    MUX_UNSIGNED #(.width(5)) u_mux_191 (
        .y(_node_109),
        .sel(_node_108),
        .a(in0_vec_12),
        .b(_node_107)
    );
    wire _node_110;
    EQ_UNSIGNED #(.width(5)) u_eq_192 (
        .y(_node_110),
        .a(5'd13),
        .b(_T_220)
    );
    wire [4:0] _node_111;
    MUX_UNSIGNED #(.width(5)) u_mux_193 (
        .y(_node_111),
        .sel(_node_110),
        .a(in0_vec_13),
        .b(_node_109)
    );
    wire _node_112;
    EQ_UNSIGNED #(.width(5)) u_eq_194 (
        .y(_node_112),
        .a(5'd14),
        .b(_T_220)
    );
    wire [4:0] _node_113;
    MUX_UNSIGNED #(.width(5)) u_mux_195 (
        .y(_node_113),
        .sel(_node_112),
        .a(in0_vec_14),
        .b(_node_111)
    );
    wire _node_114;
    EQ_UNSIGNED #(.width(5)) u_eq_196 (
        .y(_node_114),
        .a(5'd15),
        .b(_T_220)
    );
    wire [4:0] _node_115;
    MUX_UNSIGNED #(.width(5)) u_mux_197 (
        .y(_node_115),
        .sel(_node_114),
        .a(in0_vec_15),
        .b(_node_113)
    );
    wire _node_116;
    EQ_UNSIGNED #(.width(5)) u_eq_198 (
        .y(_node_116),
        .a(5'd16),
        .b(_T_220)
    );
    wire [4:0] _node_117;
    MUX_UNSIGNED #(.width(5)) u_mux_199 (
        .y(_node_117),
        .sel(_node_116),
        .a(in0_vec_16),
        .b(_node_115)
    );
    wire _node_118;
    EQ_UNSIGNED #(.width(5)) u_eq_200 (
        .y(_node_118),
        .a(5'd17),
        .b(_T_220)
    );
    wire [4:0] _node_119;
    MUX_UNSIGNED #(.width(5)) u_mux_201 (
        .y(_node_119),
        .sel(_node_118),
        .a(in0_vec_17),
        .b(_node_117)
    );
    wire _node_120;
    EQ_UNSIGNED #(.width(5)) u_eq_202 (
        .y(_node_120),
        .a(5'd18),
        .b(_T_220)
    );
    wire [4:0] _node_121;
    MUX_UNSIGNED #(.width(5)) u_mux_203 (
        .y(_node_121),
        .sel(_node_120),
        .a(in0_vec_18),
        .b(_node_119)
    );
    wire _node_122;
    EQ_UNSIGNED #(.width(5)) u_eq_204 (
        .y(_node_122),
        .a(5'd19),
        .b(_T_220)
    );
    wire [4:0] _node_123;
    MUX_UNSIGNED #(.width(5)) u_mux_205 (
        .y(_node_123),
        .sel(_node_122),
        .a(in0_vec_19),
        .b(_node_121)
    );
    wire _node_124;
    EQ_UNSIGNED #(.width(5)) u_eq_206 (
        .y(_node_124),
        .a(5'd0),
        .b(_T_222)
    );
    wire [4:0] _node_125;
    assign _node_125 = in1_vec_0;
    wire _node_126;
    EQ_UNSIGNED #(.width(5)) u_eq_207 (
        .y(_node_126),
        .a(5'd1),
        .b(_T_222)
    );
    wire [4:0] _node_127;
    MUX_UNSIGNED #(.width(5)) u_mux_208 (
        .y(_node_127),
        .sel(_node_126),
        .a(in1_vec_1),
        .b(_node_125)
    );
    wire _node_128;
    EQ_UNSIGNED #(.width(5)) u_eq_209 (
        .y(_node_128),
        .a(5'd2),
        .b(_T_222)
    );
    wire [4:0] _node_129;
    MUX_UNSIGNED #(.width(5)) u_mux_210 (
        .y(_node_129),
        .sel(_node_128),
        .a(in1_vec_2),
        .b(_node_127)
    );
    wire _node_130;
    EQ_UNSIGNED #(.width(5)) u_eq_211 (
        .y(_node_130),
        .a(5'd3),
        .b(_T_222)
    );
    wire [4:0] _node_131;
    MUX_UNSIGNED #(.width(5)) u_mux_212 (
        .y(_node_131),
        .sel(_node_130),
        .a(in1_vec_3),
        .b(_node_129)
    );
    wire _node_132;
    EQ_UNSIGNED #(.width(5)) u_eq_213 (
        .y(_node_132),
        .a(5'd4),
        .b(_T_222)
    );
    wire [4:0] _node_133;
    MUX_UNSIGNED #(.width(5)) u_mux_214 (
        .y(_node_133),
        .sel(_node_132),
        .a(in1_vec_4),
        .b(_node_131)
    );
    wire _node_134;
    EQ_UNSIGNED #(.width(5)) u_eq_215 (
        .y(_node_134),
        .a(5'd5),
        .b(_T_222)
    );
    wire [4:0] _node_135;
    MUX_UNSIGNED #(.width(5)) u_mux_216 (
        .y(_node_135),
        .sel(_node_134),
        .a(in1_vec_5),
        .b(_node_133)
    );
    wire _node_136;
    EQ_UNSIGNED #(.width(5)) u_eq_217 (
        .y(_node_136),
        .a(5'd6),
        .b(_T_222)
    );
    wire [4:0] _node_137;
    MUX_UNSIGNED #(.width(5)) u_mux_218 (
        .y(_node_137),
        .sel(_node_136),
        .a(in1_vec_6),
        .b(_node_135)
    );
    wire _node_138;
    EQ_UNSIGNED #(.width(5)) u_eq_219 (
        .y(_node_138),
        .a(5'd7),
        .b(_T_222)
    );
    wire [4:0] _node_139;
    MUX_UNSIGNED #(.width(5)) u_mux_220 (
        .y(_node_139),
        .sel(_node_138),
        .a(in1_vec_7),
        .b(_node_137)
    );
    wire _node_140;
    EQ_UNSIGNED #(.width(5)) u_eq_221 (
        .y(_node_140),
        .a(5'd8),
        .b(_T_222)
    );
    wire [4:0] _node_141;
    MUX_UNSIGNED #(.width(5)) u_mux_222 (
        .y(_node_141),
        .sel(_node_140),
        .a(in1_vec_8),
        .b(_node_139)
    );
    wire _node_142;
    EQ_UNSIGNED #(.width(5)) u_eq_223 (
        .y(_node_142),
        .a(5'd9),
        .b(_T_222)
    );
    wire [4:0] _node_143;
    MUX_UNSIGNED #(.width(5)) u_mux_224 (
        .y(_node_143),
        .sel(_node_142),
        .a(in1_vec_9),
        .b(_node_141)
    );
    wire _node_144;
    EQ_UNSIGNED #(.width(5)) u_eq_225 (
        .y(_node_144),
        .a(5'd10),
        .b(_T_222)
    );
    wire [4:0] _node_145;
    MUX_UNSIGNED #(.width(5)) u_mux_226 (
        .y(_node_145),
        .sel(_node_144),
        .a(in1_vec_10),
        .b(_node_143)
    );
    wire _node_146;
    EQ_UNSIGNED #(.width(5)) u_eq_227 (
        .y(_node_146),
        .a(5'd11),
        .b(_T_222)
    );
    wire [4:0] _node_147;
    MUX_UNSIGNED #(.width(5)) u_mux_228 (
        .y(_node_147),
        .sel(_node_146),
        .a(in1_vec_11),
        .b(_node_145)
    );
    wire _node_148;
    EQ_UNSIGNED #(.width(5)) u_eq_229 (
        .y(_node_148),
        .a(5'd12),
        .b(_T_222)
    );
    wire [4:0] _node_149;
    MUX_UNSIGNED #(.width(5)) u_mux_230 (
        .y(_node_149),
        .sel(_node_148),
        .a(in1_vec_12),
        .b(_node_147)
    );
    wire _node_150;
    EQ_UNSIGNED #(.width(5)) u_eq_231 (
        .y(_node_150),
        .a(5'd13),
        .b(_T_222)
    );
    wire [4:0] _node_151;
    MUX_UNSIGNED #(.width(5)) u_mux_232 (
        .y(_node_151),
        .sel(_node_150),
        .a(in1_vec_13),
        .b(_node_149)
    );
    wire _node_152;
    EQ_UNSIGNED #(.width(5)) u_eq_233 (
        .y(_node_152),
        .a(5'd14),
        .b(_T_222)
    );
    wire [4:0] _node_153;
    MUX_UNSIGNED #(.width(5)) u_mux_234 (
        .y(_node_153),
        .sel(_node_152),
        .a(in1_vec_14),
        .b(_node_151)
    );
    wire _node_154;
    EQ_UNSIGNED #(.width(5)) u_eq_235 (
        .y(_node_154),
        .a(5'd15),
        .b(_T_222)
    );
    wire [4:0] _node_155;
    MUX_UNSIGNED #(.width(5)) u_mux_236 (
        .y(_node_155),
        .sel(_node_154),
        .a(in1_vec_15),
        .b(_node_153)
    );
    wire _node_156;
    EQ_UNSIGNED #(.width(5)) u_eq_237 (
        .y(_node_156),
        .a(5'd16),
        .b(_T_222)
    );
    wire [4:0] _node_157;
    MUX_UNSIGNED #(.width(5)) u_mux_238 (
        .y(_node_157),
        .sel(_node_156),
        .a(in1_vec_16),
        .b(_node_155)
    );
    wire _node_158;
    EQ_UNSIGNED #(.width(5)) u_eq_239 (
        .y(_node_158),
        .a(5'd17),
        .b(_T_222)
    );
    wire [4:0] _node_159;
    MUX_UNSIGNED #(.width(5)) u_mux_240 (
        .y(_node_159),
        .sel(_node_158),
        .a(in1_vec_17),
        .b(_node_157)
    );
    wire _node_160;
    EQ_UNSIGNED #(.width(5)) u_eq_241 (
        .y(_node_160),
        .a(5'd18),
        .b(_T_222)
    );
    wire [4:0] _node_161;
    MUX_UNSIGNED #(.width(5)) u_mux_242 (
        .y(_node_161),
        .sel(_node_160),
        .a(in1_vec_18),
        .b(_node_159)
    );
    wire _node_162;
    EQ_UNSIGNED #(.width(5)) u_eq_243 (
        .y(_node_162),
        .a(5'd19),
        .b(_T_222)
    );
    wire [4:0] _node_163;
    MUX_UNSIGNED #(.width(5)) u_mux_244 (
        .y(_node_163),
        .sel(_node_162),
        .a(in1_vec_19),
        .b(_node_161)
    );
    wire [5:0] _T_223;
    ADD_UNSIGNED #(.width(5)) u_add_245 (
        .y(_T_223),
        .a(_node_123),
        .b(_node_163)
    );
    wire [4:0] _T_224;
    TAIL #(.width(6), .n(1)) tail_246 (
        .y(_T_224),
        .in(_T_223)
    );
    wire _node_164;
    EQ_UNSIGNED #(.width(5)) u_eq_247 (
        .y(_node_164),
        .a(5'd0),
        .b(_T_218)
    );
    wire [4:0] _node_165;
    assign _node_165 = expected_out_vec_0;
    wire _node_166;
    EQ_UNSIGNED #(.width(5)) u_eq_248 (
        .y(_node_166),
        .a(5'd1),
        .b(_T_218)
    );
    wire [4:0] _node_167;
    MUX_UNSIGNED #(.width(5)) u_mux_249 (
        .y(_node_167),
        .sel(_node_166),
        .a(expected_out_vec_1),
        .b(_node_165)
    );
    wire _node_168;
    EQ_UNSIGNED #(.width(5)) u_eq_250 (
        .y(_node_168),
        .a(5'd2),
        .b(_T_218)
    );
    wire [4:0] _node_169;
    MUX_UNSIGNED #(.width(5)) u_mux_251 (
        .y(_node_169),
        .sel(_node_168),
        .a(expected_out_vec_2),
        .b(_node_167)
    );
    wire _node_170;
    EQ_UNSIGNED #(.width(5)) u_eq_252 (
        .y(_node_170),
        .a(5'd3),
        .b(_T_218)
    );
    wire [4:0] _node_171;
    MUX_UNSIGNED #(.width(5)) u_mux_253 (
        .y(_node_171),
        .sel(_node_170),
        .a(expected_out_vec_3),
        .b(_node_169)
    );
    wire _node_172;
    EQ_UNSIGNED #(.width(5)) u_eq_254 (
        .y(_node_172),
        .a(5'd4),
        .b(_T_218)
    );
    wire [4:0] _node_173;
    MUX_UNSIGNED #(.width(5)) u_mux_255 (
        .y(_node_173),
        .sel(_node_172),
        .a(expected_out_vec_4),
        .b(_node_171)
    );
    wire _node_174;
    EQ_UNSIGNED #(.width(5)) u_eq_256 (
        .y(_node_174),
        .a(5'd5),
        .b(_T_218)
    );
    wire [4:0] _node_175;
    MUX_UNSIGNED #(.width(5)) u_mux_257 (
        .y(_node_175),
        .sel(_node_174),
        .a(expected_out_vec_5),
        .b(_node_173)
    );
    wire _node_176;
    EQ_UNSIGNED #(.width(5)) u_eq_258 (
        .y(_node_176),
        .a(5'd6),
        .b(_T_218)
    );
    wire [4:0] _node_177;
    MUX_UNSIGNED #(.width(5)) u_mux_259 (
        .y(_node_177),
        .sel(_node_176),
        .a(expected_out_vec_6),
        .b(_node_175)
    );
    wire _node_178;
    EQ_UNSIGNED #(.width(5)) u_eq_260 (
        .y(_node_178),
        .a(5'd7),
        .b(_T_218)
    );
    wire [4:0] _node_179;
    MUX_UNSIGNED #(.width(5)) u_mux_261 (
        .y(_node_179),
        .sel(_node_178),
        .a(expected_out_vec_7),
        .b(_node_177)
    );
    wire _node_180;
    EQ_UNSIGNED #(.width(5)) u_eq_262 (
        .y(_node_180),
        .a(5'd8),
        .b(_T_218)
    );
    wire [4:0] _node_181;
    MUX_UNSIGNED #(.width(5)) u_mux_263 (
        .y(_node_181),
        .sel(_node_180),
        .a(expected_out_vec_8),
        .b(_node_179)
    );
    wire _node_182;
    EQ_UNSIGNED #(.width(5)) u_eq_264 (
        .y(_node_182),
        .a(5'd9),
        .b(_T_218)
    );
    wire [4:0] _node_183;
    MUX_UNSIGNED #(.width(5)) u_mux_265 (
        .y(_node_183),
        .sel(_node_182),
        .a(expected_out_vec_9),
        .b(_node_181)
    );
    wire _node_184;
    EQ_UNSIGNED #(.width(5)) u_eq_266 (
        .y(_node_184),
        .a(5'd10),
        .b(_T_218)
    );
    wire [4:0] _node_185;
    MUX_UNSIGNED #(.width(5)) u_mux_267 (
        .y(_node_185),
        .sel(_node_184),
        .a(expected_out_vec_10),
        .b(_node_183)
    );
    wire _node_186;
    EQ_UNSIGNED #(.width(5)) u_eq_268 (
        .y(_node_186),
        .a(5'd11),
        .b(_T_218)
    );
    wire [4:0] _node_187;
    MUX_UNSIGNED #(.width(5)) u_mux_269 (
        .y(_node_187),
        .sel(_node_186),
        .a(expected_out_vec_11),
        .b(_node_185)
    );
    wire _node_188;
    EQ_UNSIGNED #(.width(5)) u_eq_270 (
        .y(_node_188),
        .a(5'd12),
        .b(_T_218)
    );
    wire [4:0] _node_189;
    MUX_UNSIGNED #(.width(5)) u_mux_271 (
        .y(_node_189),
        .sel(_node_188),
        .a(expected_out_vec_12),
        .b(_node_187)
    );
    wire _node_190;
    EQ_UNSIGNED #(.width(5)) u_eq_272 (
        .y(_node_190),
        .a(5'd13),
        .b(_T_218)
    );
    wire [4:0] _node_191;
    MUX_UNSIGNED #(.width(5)) u_mux_273 (
        .y(_node_191),
        .sel(_node_190),
        .a(expected_out_vec_13),
        .b(_node_189)
    );
    wire _node_192;
    EQ_UNSIGNED #(.width(5)) u_eq_274 (
        .y(_node_192),
        .a(5'd14),
        .b(_T_218)
    );
    wire [4:0] _node_193;
    MUX_UNSIGNED #(.width(5)) u_mux_275 (
        .y(_node_193),
        .sel(_node_192),
        .a(expected_out_vec_14),
        .b(_node_191)
    );
    wire _node_194;
    EQ_UNSIGNED #(.width(5)) u_eq_276 (
        .y(_node_194),
        .a(5'd15),
        .b(_T_218)
    );
    wire [4:0] _node_195;
    MUX_UNSIGNED #(.width(5)) u_mux_277 (
        .y(_node_195),
        .sel(_node_194),
        .a(expected_out_vec_15),
        .b(_node_193)
    );
    wire _node_196;
    EQ_UNSIGNED #(.width(5)) u_eq_278 (
        .y(_node_196),
        .a(5'd16),
        .b(_T_218)
    );
    wire [4:0] _node_197;
    MUX_UNSIGNED #(.width(5)) u_mux_279 (
        .y(_node_197),
        .sel(_node_196),
        .a(expected_out_vec_16),
        .b(_node_195)
    );
    wire _node_198;
    EQ_UNSIGNED #(.width(5)) u_eq_280 (
        .y(_node_198),
        .a(5'd17),
        .b(_T_218)
    );
    wire [4:0] _node_199;
    MUX_UNSIGNED #(.width(5)) u_mux_281 (
        .y(_node_199),
        .sel(_node_198),
        .a(expected_out_vec_17),
        .b(_node_197)
    );
    wire _node_200;
    EQ_UNSIGNED #(.width(5)) u_eq_282 (
        .y(_node_200),
        .a(5'd18),
        .b(_T_218)
    );
    wire [4:0] _node_201;
    MUX_UNSIGNED #(.width(5)) u_mux_283 (
        .y(_node_201),
        .sel(_node_200),
        .a(expected_out_vec_18),
        .b(_node_199)
    );
    wire _node_202;
    EQ_UNSIGNED #(.width(5)) u_eq_284 (
        .y(_node_202),
        .a(5'd19),
        .b(_T_218)
    );
    wire [4:0] _node_203;
    MUX_UNSIGNED #(.width(5)) u_mux_285 (
        .y(_node_203),
        .sel(_node_202),
        .a(expected_out_vec_19),
        .b(_node_201)
    );
    wire _T_225;
    EQ_UNSIGNED #(.width(5)) u_eq_286 (
        .y(_T_225),
        .a(_node_203),
        .b(_T_224)
    );
    wire _T_226;
    BITWISEOR #(.width(1)) bitwiseor_287 (
        .y(_T_226),
        .a(_T_225),
        .b(reset)
    );
    wire _T_228;
    EQ_UNSIGNED #(.width(1)) u_eq_288 (
        .y(_T_228),
        .a(_T_226),
        .b(1'h0)
    );
    wire [32:0] _T_230;
    wire [31:0] _WTEMP_12;
    PAD_UNSIGNED #(.width(1), .n(32)) u_pad_289 (
        .y(_WTEMP_12),
        .in(1'h1)
    );
    ADD_UNSIGNED #(.width(32)) u_add_290 (
        .y(_T_230),
        .a(_test_number__q),
        .b(_WTEMP_12)
    );
    wire [31:0] _T_231;
    TAIL #(.width(33), .n(1)) tail_291 (
        .y(_T_231),
        .in(_T_230)
    );
    wire _T_233;
    EQ_UNSIGNED #(.width(1)) u_eq_292 (
        .y(_T_233),
        .a(reset),
        .b(1'h0)
    );
    wire [32:0] _T_236;
    wire [31:0] _WTEMP_13;
    PAD_UNSIGNED #(.width(1), .n(32)) u_pad_293 (
        .y(_WTEMP_13),
        .in(1'h1)
    );
    ADD_UNSIGNED #(.width(32)) u_add_294 (
        .y(_T_236),
        .a(_state_number__q),
        .b(_WTEMP_13)
    );
    wire [31:0] _T_237;
    TAIL #(.width(33), .n(1)) tail_295 (
        .y(_T_237),
        .in(_T_236)
    );
    wire _node_204;
    MUX_UNSIGNED #(.width(1)) u_mux_296 (
        .y(_node_204),
        .sel(_T_196),
        .a(1'h1),
        .b(_node_1)
    );
    wire [31:0] _node_205;
    wire [31:0] _WTEMP_14;
    PAD_UNSIGNED #(.width(6), .n(32)) u_pad_297 (
        .y(_WTEMP_14),
        .in(6'h21)
    );
    MUX_UNSIGNED #(.width(32)) u_mux_298 (
        .y(_node_205),
        .sel(_T_196),
        .a(_WTEMP_14),
        .b(_node_2)
    );
    wire [31:0] _node_206;
    wire [31:0] _WTEMP_15;
    PAD_UNSIGNED #(.width(7), .n(32)) u_pad_299 (
        .y(_WTEMP_15),
        .in(7'h64)
    );
    MUX_UNSIGNED #(.width(32)) u_mux_300 (
        .y(_node_206),
        .sel(_T_196),
        .a(_WTEMP_15),
        .b(_max_ticks_for_state__q)
    );
    wire _node_207;
    MUX_UNSIGNED #(.width(1)) u_mux_301 (
        .y(_node_207),
        .sel(_T_192),
        .a(1'h0),
        .b(_node_204)
    );
    wire _node_208;
    MUX_UNSIGNED #(.width(1)) u_mux_302 (
        .y(_node_208),
        .sel(_T_22),
        .a(1'h0),
        .b(_state_locked__q)
    );
    wire [31:0] _node_209;
    MUX_UNSIGNED #(.width(32)) u_mux_303 (
        .y(_node_209),
        .sel(_T_192),
        .a(_T_237),
        .b(_node_205)
    );
    wire [31:0] _node_210;
    MUX_UNSIGNED #(.width(32)) u_mux_304 (
        .y(_node_210),
        .sel(_T_22),
        .a(_T_28),
        .b(_node_0)
    );
    wire [31:0] _node_211;
    wire [31:0] _WTEMP_16;
    PAD_UNSIGNED #(.width(1), .n(32)) u_pad_305 (
        .y(_WTEMP_16),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(32)) u_mux_306 (
        .y(_node_211),
        .sel(_T_196),
        .a(_WTEMP_16),
        .b(_node_3)
    );
    wire [31:0] _node_212;
    wire [31:0] _WTEMP_17;
    PAD_UNSIGNED #(.width(1), .n(32)) u_pad_307 (
        .y(_WTEMP_17),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(32)) u_mux_308 (
        .y(_node_212),
        .sel(_T_14),
        .a(_WTEMP_17),
        .b(_T_12)
    );
    wire _T_239;
    wire [31:0] _WTEMP_18;
    PAD_UNSIGNED #(.width(6), .n(32)) u_pad_309 (
        .y(_WTEMP_18),
        .in(6'h22)
    );
    GT_UNSIGNED #(.width(32)) u_gt_310 (
        .y(_T_239),
        .a(_state_number__q),
        .b(_WTEMP_18)
    );
    wire _T_241;
    EQ_UNSIGNED #(.width(1)) u_eq_311 (
        .y(_T_241),
        .a(reset),
        .b(1'h0)
    );
    wire _T_243;
    EQ_UNSIGNED #(.width(1)) u_eq_312 (
        .y(_T_243),
        .a(reset),
        .b(1'h0)
    );
    wire _T_245;
    wire [31:0] _WTEMP_19;
    PAD_UNSIGNED #(.width(6), .n(32)) u_pad_313 (
        .y(_WTEMP_19),
        .in(6'h22)
    );
    GT_UNSIGNED #(.width(32)) u_gt_314 (
        .y(_T_245),
        .a(_state_number__q),
        .b(_WTEMP_19)
    );
    wire _T_247;
    EQ_UNSIGNED #(.width(1)) u_eq_315 (
        .y(_T_247),
        .a(reset),
        .b(1'h0)
    );
    wire _T_249;
    EQ_UNSIGNED #(.width(1)) u_eq_316 (
        .y(_T_249),
        .a(reset),
        .b(1'h0)
    );
    assign _c__clock = clock;
    assign _c__reset = reset;
    assign expected_out_vec_0 = _T_126;
    assign expected_out_vec_1 = _T_128;
    assign expected_out_vec_10 = _T_146;
    assign expected_out_vec_11 = _T_148;
    assign expected_out_vec_12 = _T_150;
    assign expected_out_vec_13 = _T_152;
    assign expected_out_vec_14 = _T_154;
    assign expected_out_vec_15 = _T_156;
    assign expected_out_vec_16 = _T_158;
    assign expected_out_vec_17 = _T_160;
    assign expected_out_vec_18 = _T_162;
    assign expected_out_vec_19 = _T_164;
    assign expected_out_vec_2 = _T_130;
    assign expected_out_vec_3 = _T_132;
    assign expected_out_vec_4 = _T_134;
    assign expected_out_vec_5 = _T_136;
    assign expected_out_vec_6 = _T_138;
    assign expected_out_vec_7 = _T_140;
    assign expected_out_vec_8 = _T_142;
    assign expected_out_vec_9 = _T_144;
    PAD_UNSIGNED #(.width(2), .n(5)) u_pad_317 (
        .y(in0_vec_0),
        .in(2'h3)
    );
    PAD_UNSIGNED #(.width(3), .n(5)) u_pad_318 (
        .y(in0_vec_1),
        .in(3'h4)
    );
    PAD_UNSIGNED #(.width(4), .n(5)) u_pad_319 (
        .y(in0_vec_10),
        .in(4'hD)
    );
    PAD_UNSIGNED #(.width(4), .n(5)) u_pad_320 (
        .y(in0_vec_11),
        .in(4'hE)
    );
    PAD_UNSIGNED #(.width(4), .n(5)) u_pad_321 (
        .y(in0_vec_12),
        .in(4'hF)
    );
    assign in0_vec_13 = 5'h10;
    assign in0_vec_14 = 5'h11;
    assign in0_vec_15 = 5'h12;
    assign in0_vec_16 = 5'h13;
    assign in0_vec_17 = 5'h14;
    assign in0_vec_18 = 5'h15;
    assign in0_vec_19 = 5'h16;
    PAD_UNSIGNED #(.width(3), .n(5)) u_pad_322 (
        .y(in0_vec_2),
        .in(3'h5)
    );
    PAD_UNSIGNED #(.width(3), .n(5)) u_pad_323 (
        .y(in0_vec_3),
        .in(3'h6)
    );
    PAD_UNSIGNED #(.width(3), .n(5)) u_pad_324 (
        .y(in0_vec_4),
        .in(3'h7)
    );
    PAD_UNSIGNED #(.width(4), .n(5)) u_pad_325 (
        .y(in0_vec_5),
        .in(4'h8)
    );
    PAD_UNSIGNED #(.width(4), .n(5)) u_pad_326 (
        .y(in0_vec_6),
        .in(4'h9)
    );
    PAD_UNSIGNED #(.width(4), .n(5)) u_pad_327 (
        .y(in0_vec_7),
        .in(4'hA)
    );
    PAD_UNSIGNED #(.width(4), .n(5)) u_pad_328 (
        .y(in0_vec_8),
        .in(4'hB)
    );
    PAD_UNSIGNED #(.width(4), .n(5)) u_pad_329 (
        .y(in0_vec_9),
        .in(4'hC)
    );
    PAD_UNSIGNED #(.width(3), .n(5)) u_pad_330 (
        .y(in1_vec_0),
        .in(3'h7)
    );
    PAD_UNSIGNED #(.width(4), .n(5)) u_pad_331 (
        .y(in1_vec_1),
        .in(4'h8)
    );
    assign in1_vec_10 = 5'h11;
    assign in1_vec_11 = 5'h12;
    assign in1_vec_12 = 5'h13;
    assign in1_vec_13 = 5'h14;
    assign in1_vec_14 = 5'h15;
    assign in1_vec_15 = 5'h16;
    assign in1_vec_16 = 5'h17;
    assign in1_vec_17 = 5'h18;
    assign in1_vec_18 = 5'h19;
    assign in1_vec_19 = 5'h1A;
    PAD_UNSIGNED #(.width(4), .n(5)) u_pad_332 (
        .y(in1_vec_2),
        .in(4'h9)
    );
    PAD_UNSIGNED #(.width(4), .n(5)) u_pad_333 (
        .y(in1_vec_3),
        .in(4'hA)
    );
    PAD_UNSIGNED #(.width(4), .n(5)) u_pad_334 (
        .y(in1_vec_4),
        .in(4'hB)
    );
    PAD_UNSIGNED #(.width(4), .n(5)) u_pad_335 (
        .y(in1_vec_5),
        .in(4'hC)
    );
    PAD_UNSIGNED #(.width(4), .n(5)) u_pad_336 (
        .y(in1_vec_6),
        .in(4'hD)
    );
    PAD_UNSIGNED #(.width(4), .n(5)) u_pad_337 (
        .y(in1_vec_7),
        .in(4'hE)
    );
    PAD_UNSIGNED #(.width(4), .n(5)) u_pad_338 (
        .y(in1_vec_8),
        .in(4'hF)
    );
    assign in1_vec_9 = 5'h10;
    MUX_UNSIGNED #(.width(32)) u_mux_339 (
        .y(_WTEMP_1),
        .sel(_T_194),
        .a(_node_206),
        .b(_max_ticks_for_state__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_340 (
        .y(_WTEMP_3),
        .sel(_T_194),
        .a(_node_207),
        .b(_node_208)
    );
    MUX_UNSIGNED #(.width(32)) u_mux_341 (
        .y(_WTEMP_2),
        .sel(_T_194),
        .a(_node_209),
        .b(_node_210)
    );
    MUX_UNSIGNED #(.width(32)) u_mux_342 (
        .y(_WTEMP_8),
        .sel(_T_194),
        .a(_T_231),
        .b(_test_number__q)
    );
    MUX_UNSIGNED #(.width(32)) u_mux_343 (
        .y(_WTEMP_0),
        .sel(_T_194),
        .a(_node_211),
        .b(_node_212)
    );
endmodule //AdderExerciser
module DFF_POSCLK(q, d, clk);
    parameter width = 4;
    output reg [width-1:0] q;
    input [width-1:0] d;
    input clk;
    always @(posedge clk) begin
        q <= d;
    end
endmodule // DFF_POSCLK
module MUX_UNSIGNED(y, sel, a, b);
    parameter width = 4;
    output [width-1:0] y;
    input sel;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = sel ? a : b;
endmodule // MUX_UNSIGNED
module PAD_UNSIGNED(y, in);
    parameter width = 4;
    parameter n = 4;
    output [(n > width ? n : width)-1:0] y;
    input [width-1:0] in;
    assign y = (n > width) ? {{(n - width){1'b0}}, in} : in;
endmodule // PAD_UNSIGNED
module ADD_UNSIGNED(y, a, b);
    parameter width = 4;
    output [width:0] y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a + b;
endmodule // ADD_UNSIGNED
module TAIL(y, in);
    parameter width = 4;
    parameter n = 2;
    output [width-n-1:0] y;
    input [width-1:0] in;
    assign y = in[width-n-1:0];
endmodule // TAIL
module EQ_UNSIGNED(y, a, b);
    parameter width = 4;
    output y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a == b;
endmodule // EQ_UNSIGNED
module GT_UNSIGNED(y, a, b);
    parameter width = 4;
    output y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a > b;
endmodule // GT_UNSIGNED
module BITWISEAND(y, a, b);
    parameter width = 4;
    output [width-1:0] y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a & b;
endmodule // BITWISEAND
module Adder(
    input clock,
    input reset,
    input [31:0] io_in0,
    input [31:0] io_in1,
    output [31:0] io_out
);
    wire [32:0] _T_5;
    ADD_UNSIGNED #(.width(32)) u_add_24 (
        .y(_T_5),
        .a(io_in0),
        .b(io_in1)
    );
    wire [31:0] _T_6;
    TAIL #(.width(33), .n(1)) tail_25 (
        .y(_T_6),
        .in(_T_5)
    );
    assign io_out = _T_6;
endmodule //Adder
module BITS(y, in);
    parameter width = 4;
    parameter high = 2;
    parameter low = 0;
    output [high-low:0] y;
    input [width-1:0] in;
    assign y = in[high:low];
endmodule // BITS
module BITWISEOR(y, a, b);
    parameter width = 4;
    output [width-1:0] y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a | b;
endmodule // BITWISEOR
