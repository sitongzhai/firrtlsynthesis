module Queue(
  input   clock
);
endmodule
