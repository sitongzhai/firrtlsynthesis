module FixedPointReduce( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  input  [63:0] io_in_0, // @[:@6.4]
  input  [63:0] io_in_1, // @[:@6.4]
  input  [63:0] io_in_2, // @[:@6.4]
  input  [63:0] io_in_3, // @[:@6.4]
  input  [63:0] io_in_4, // @[:@6.4]
  input  [63:0] io_in_5, // @[:@6.4]
  input  [63:0] io_in_6, // @[:@6.4]
  input  [63:0] io_in_7, // @[:@6.4]
  input  [63:0] io_in_8, // @[:@6.4]
  input  [63:0] io_in_9, // @[:@6.4]
  output [63:0] io_sum // @[:@6.4]
);
  wire [63:0] _T_18 = $signed(io_in_0) + $signed(io_in_1); // @[FixedPointSpec.scala 16:28:@13.4]
  wire [63:0] _T_21 = $signed(_T_18) + $signed(io_in_2); // @[FixedPointSpec.scala 16:28:@16.4]
  wire [63:0] _T_24 = $signed(_T_21) + $signed(io_in_3); // @[FixedPointSpec.scala 16:28:@19.4]
  wire [63:0] _T_27 = $signed(_T_24) + $signed(io_in_4); // @[FixedPointSpec.scala 16:28:@22.4]
  wire [63:0] _T_30 = $signed(_T_27) + $signed(io_in_5); // @[FixedPointSpec.scala 16:28:@25.4]
  wire [63:0] _T_33 = $signed(_T_30) + $signed(io_in_6); // @[FixedPointSpec.scala 16:28:@28.4]
  wire [63:0] _T_36 = $signed(_T_33) + $signed(io_in_7); // @[FixedPointSpec.scala 16:28:@31.4]
  wire [63:0] _T_39 = $signed(_T_36) + $signed(io_in_8); // @[FixedPointSpec.scala 16:28:@34.4]
  assign io_sum = $signed(_T_39) + $signed(io_in_9); // @[FixedPointSpec.scala 16:28:@37.4]
endmodule
