module SmallOdds3Tester(
    input clock,
    input reset
);
    wire _device_under_test__clock;
    wire _device_under_test__reset;
    wire _device_under_test__io_in_ready;
    wire _device_under_test__io_in_valid;
    wire [31:0] _device_under_test__io_in_bits;
    wire _device_under_test__io_out_ready;
    wire _device_under_test__io_out_valid;
    wire [31:0] _device_under_test__io_out_bits;
    SmallOdds3 device_under_test (
        .clock(_device_under_test__clock),
        .reset(_device_under_test__reset),
        .io_in_ready(_device_under_test__io_in_ready),
        .io_in_valid(_device_under_test__io_in_valid),
        .io_in_bits(_device_under_test__io_in_bits),
        .io_out_ready(_device_under_test__io_out_ready),
        .io_out_valid(_device_under_test__io_out_valid),
        .io_out_bits(_device_under_test__io_out_bits)
    );
    wire [8:0] __T_4__q;
    wire [8:0] __T_4__d;
    DFF_POSCLK #(.width(9)) _T_4 (
        .q(__T_4__q),
        .d(__T_4__d),
        .clk(clock)
    );
    wire [8:0] _WTEMP_4;
    MUX_UNSIGNED #(.width(9)) u_mux_24 (
        .y(__T_4__d),
        .sel(reset),
        .a(9'h0),
        .b(_WTEMP_4)
    );
    wire __T_7__q;
    wire __T_7__d;
    DFF_POSCLK #(.width(1)) _T_7 (
        .q(__T_7__q),
        .d(__T_7__d),
        .clk(clock)
    );
    wire _WTEMP_5;
    MUX_UNSIGNED #(.width(1)) u_mux_25 (
        .y(__T_7__d),
        .sel(reset),
        .a(1'h0),
        .b(_WTEMP_5)
    );
    wire [6:0] __T_10__q;
    wire [6:0] __T_10__d;
    DFF_POSCLK #(.width(7)) _T_10 (
        .q(__T_10__q),
        .d(__T_10__d),
        .clk(clock)
    );
    wire [6:0] _WTEMP_6;
    MUX_UNSIGNED #(.width(7)) u_mux_26 (
        .y(__T_10__d),
        .sel(reset),
        .a(7'h0),
        .b(_WTEMP_6)
    );
    wire __T_13__q;
    wire __T_13__d;
    DFF_POSCLK #(.width(1)) _T_13 (
        .q(__T_13__q),
        .d(__T_13__d),
        .clk(clock)
    );
    wire _WTEMP_7;
    MUX_UNSIGNED #(.width(1)) u_mux_27 (
        .y(__T_13__d),
        .sel(reset),
        .a(1'h0),
        .b(_WTEMP_7)
    );
    wire _T_14;
    BITWISEAND #(.width(1)) bitwiseand_28 (
        .y(_T_14),
        .a(__T_7__q),
        .b(__T_13__q)
    );
    wire _T_16;
    EQ_UNSIGNED #(.width(1)) u_eq_29 (
        .y(_T_16),
        .a(reset),
        .b(1'h0)
    );
    wire _T_18;
    EQ_UNSIGNED #(.width(1)) u_eq_30 (
        .y(_T_18),
        .a(reset),
        .b(1'h0)
    );
    wire [13:0] __T_21__q;
    wire [13:0] __T_21__d;
    DFF_POSCLK #(.width(14)) _T_21 (
        .q(__T_21__q),
        .d(__T_21__d),
        .clk(clock)
    );
    wire [13:0] _WTEMP_8;
    MUX_UNSIGNED #(.width(14)) u_mux_31 (
        .y(__T_21__d),
        .sel(reset),
        .a(14'h0),
        .b(_WTEMP_8)
    );
    wire [14:0] _T_23;
    wire [13:0] _WTEMP_9;
    PAD_UNSIGNED #(.width(1), .n(14)) u_pad_32 (
        .y(_WTEMP_9),
        .in(1'h1)
    );
    ADD_UNSIGNED #(.width(14)) u_add_33 (
        .y(_T_23),
        .a(__T_21__q),
        .b(_WTEMP_9)
    );
    wire [13:0] _T_24;
    TAIL #(.width(15), .n(1)) tail_34 (
        .y(_T_24),
        .in(_T_23)
    );
    wire _T_26;
    GT_UNSIGNED #(.width(14)) u_gt_35 (
        .y(_T_26),
        .a(__T_21__q),
        .b(14'h2710)
    );
    wire _T_29;
    EQ_UNSIGNED #(.width(1)) u_eq_36 (
        .y(_T_29),
        .a(reset),
        .b(1'h0)
    );
    wire _T_31;
    EQ_UNSIGNED #(.width(1)) u_eq_37 (
        .y(_T_31),
        .a(reset),
        .b(1'h0)
    );
    wire _T_136_0;
    wire _T_136_1;
    wire _T_136_2;
    wire _T_136_3;
    wire _T_136_4;
    wire _T_136_5;
    wire _T_136_6;
    wire _T_136_7;
    wire _T_136_8;
    wire _T_136_9;
    wire _T_136_10;
    wire _T_136_11;
    wire _T_136_12;
    wire _T_136_13;
    wire _T_136_14;
    wire _T_136_15;
    wire _T_136_16;
    wire _T_136_17;
    wire _T_136_18;
    wire _T_136_19;
    wire _T_136_20;
    wire _T_136_21;
    wire _T_136_22;
    wire _T_136_23;
    wire _T_136_24;
    wire _T_136_25;
    wire _T_136_26;
    wire _T_136_27;
    wire _T_136_28;
    wire _T_136_29;
    wire _T_136_30;
    wire _T_136_31;
    wire _T_136_32;
    wire _T_136_33;
    wire _T_136_34;
    wire _T_136_35;
    wire _T_136_36;
    wire _T_136_37;
    wire _T_136_38;
    wire _T_136_39;
    wire _T_136_40;
    wire _T_136_41;
    wire _T_136_42;
    wire _T_136_43;
    wire _T_136_44;
    wire _T_136_45;
    wire _T_136_46;
    wire _T_136_47;
    wire _T_136_48;
    wire _T_136_49;
    wire _T_136_50;
    wire _T_136_51;
    wire _T_136_52;
    wire _T_136_53;
    wire _T_136_54;
    wire _T_136_55;
    wire _T_136_56;
    wire _T_136_57;
    wire _T_136_58;
    wire _T_136_59;
    wire _T_136_60;
    wire _T_136_61;
    wire _T_136_62;
    wire _T_136_63;
    wire _T_136_64;
    wire _T_136_65;
    wire _T_136_66;
    wire _T_136_67;
    wire _T_136_68;
    wire _T_136_69;
    wire _T_136_70;
    wire _T_136_71;
    wire _T_136_72;
    wire _T_136_73;
    wire _T_136_74;
    wire _T_136_75;
    wire _T_136_76;
    wire _T_136_77;
    wire _T_136_78;
    wire _T_136_79;
    wire _T_136_80;
    wire _T_136_81;
    wire _T_136_82;
    wire _T_136_83;
    wire _T_136_84;
    wire _T_136_85;
    wire _T_136_86;
    wire _T_136_87;
    wire _T_136_88;
    wire _T_136_89;
    wire _T_136_90;
    wire _T_136_91;
    wire _T_136_92;
    wire _T_136_93;
    wire _T_136_94;
    wire _T_136_95;
    wire _T_136_96;
    wire _T_136_97;
    wire _T_136_98;
    wire _T_136_99;
    wire _T_136_100;
    wire _T_136_101;
    wire [6:0] _value__q;
    wire [6:0] _value__d;
    DFF_POSCLK #(.width(7)) value (
        .q(_value__q),
        .d(_value__d),
        .clk(clock)
    );
    wire [6:0] _WTEMP_10;
    MUX_UNSIGNED #(.width(7)) u_mux_38 (
        .y(_value__d),
        .sel(reset),
        .a(7'h0),
        .b(_WTEMP_10)
    );
    wire [4:0] _T_347_0;
    wire [4:0] _T_347_1;
    wire [4:0] _T_347_2;
    wire [4:0] _T_347_3;
    wire [4:0] _T_347_4;
    wire [4:0] _T_347_5;
    wire [4:0] _T_347_6;
    wire [4:0] _T_347_7;
    wire [4:0] _T_347_8;
    wire [4:0] _T_347_9;
    wire [4:0] _T_347_10;
    wire [4:0] _T_347_11;
    wire [4:0] _T_347_12;
    wire [4:0] _T_347_13;
    wire [4:0] _T_347_14;
    wire [4:0] _T_347_15;
    wire [4:0] _T_347_16;
    wire [4:0] _T_347_17;
    wire [4:0] _T_347_18;
    wire [4:0] _T_347_19;
    wire [4:0] _T_347_20;
    wire [4:0] _T_347_21;
    wire [4:0] _T_347_22;
    wire [4:0] _T_347_23;
    wire [4:0] _T_347_24;
    wire [4:0] _T_347_25;
    wire [4:0] _T_347_26;
    wire [4:0] _T_347_27;
    wire [4:0] _T_347_28;
    wire [4:0] _T_347_29;
    wire [4:0] _T_347_30;
    wire [4:0] _T_347_31;
    wire [4:0] _T_347_32;
    wire [4:0] _T_347_33;
    wire [4:0] _T_347_34;
    wire [4:0] _T_347_35;
    wire [4:0] _T_347_36;
    wire [4:0] _T_347_37;
    wire [4:0] _T_347_38;
    wire [4:0] _T_347_39;
    wire [4:0] _T_347_40;
    wire [4:0] _T_347_41;
    wire [4:0] _T_347_42;
    wire [4:0] _T_347_43;
    wire [4:0] _T_347_44;
    wire [4:0] _T_347_45;
    wire [4:0] _T_347_46;
    wire [4:0] _T_347_47;
    wire [4:0] _T_347_48;
    wire [4:0] _T_347_49;
    wire [4:0] _T_347_50;
    wire [4:0] _T_347_51;
    wire [4:0] _T_347_52;
    wire [4:0] _T_347_53;
    wire [4:0] _T_347_54;
    wire [4:0] _T_347_55;
    wire [4:0] _T_347_56;
    wire [4:0] _T_347_57;
    wire [4:0] _T_347_58;
    wire [4:0] _T_347_59;
    wire [4:0] _T_347_60;
    wire [4:0] _T_347_61;
    wire [4:0] _T_347_62;
    wire [4:0] _T_347_63;
    wire [4:0] _T_347_64;
    wire [4:0] _T_347_65;
    wire [4:0] _T_347_66;
    wire [4:0] _T_347_67;
    wire [4:0] _T_347_68;
    wire [4:0] _T_347_69;
    wire [4:0] _T_347_70;
    wire [4:0] _T_347_71;
    wire [4:0] _T_347_72;
    wire [4:0] _T_347_73;
    wire [4:0] _T_347_74;
    wire [4:0] _T_347_75;
    wire [4:0] _T_347_76;
    wire [4:0] _T_347_77;
    wire [4:0] _T_347_78;
    wire [4:0] _T_347_79;
    wire [4:0] _T_347_80;
    wire [4:0] _T_347_81;
    wire [4:0] _T_347_82;
    wire [4:0] _T_347_83;
    wire [4:0] _T_347_84;
    wire [4:0] _T_347_85;
    wire [4:0] _T_347_86;
    wire [4:0] _T_347_87;
    wire [4:0] _T_347_88;
    wire [4:0] _T_347_89;
    wire [4:0] _T_347_90;
    wire [4:0] _T_347_91;
    wire [4:0] _T_347_92;
    wire [4:0] _T_347_93;
    wire [4:0] _T_347_94;
    wire [4:0] _T_347_95;
    wire [4:0] _T_347_96;
    wire [4:0] _T_347_97;
    wire [4:0] _T_347_98;
    wire [4:0] _T_347_99;
    wire [4:0] _T_347_100;
    wire [4:0] _T_347_101;
    wire _node_0;
    EQ_UNSIGNED #(.width(7)) u_eq_39 (
        .y(_node_0),
        .a(7'd0),
        .b(_value__q)
    );
    wire [4:0] _node_1;
    assign _node_1 = _T_347_0;
    wire _node_2;
    EQ_UNSIGNED #(.width(7)) u_eq_40 (
        .y(_node_2),
        .a(7'd1),
        .b(_value__q)
    );
    wire [4:0] _node_3;
    MUX_UNSIGNED #(.width(5)) u_mux_41 (
        .y(_node_3),
        .sel(_node_2),
        .a(_T_347_1),
        .b(_node_1)
    );
    wire _node_4;
    EQ_UNSIGNED #(.width(7)) u_eq_42 (
        .y(_node_4),
        .a(7'd2),
        .b(_value__q)
    );
    wire [4:0] _node_5;
    MUX_UNSIGNED #(.width(5)) u_mux_43 (
        .y(_node_5),
        .sel(_node_4),
        .a(_T_347_2),
        .b(_node_3)
    );
    wire _node_6;
    EQ_UNSIGNED #(.width(7)) u_eq_44 (
        .y(_node_6),
        .a(7'd3),
        .b(_value__q)
    );
    wire [4:0] _node_7;
    MUX_UNSIGNED #(.width(5)) u_mux_45 (
        .y(_node_7),
        .sel(_node_6),
        .a(_T_347_3),
        .b(_node_5)
    );
    wire _node_8;
    EQ_UNSIGNED #(.width(7)) u_eq_46 (
        .y(_node_8),
        .a(7'd4),
        .b(_value__q)
    );
    wire [4:0] _node_9;
    MUX_UNSIGNED #(.width(5)) u_mux_47 (
        .y(_node_9),
        .sel(_node_8),
        .a(_T_347_4),
        .b(_node_7)
    );
    wire _node_10;
    EQ_UNSIGNED #(.width(7)) u_eq_48 (
        .y(_node_10),
        .a(7'd5),
        .b(_value__q)
    );
    wire [4:0] _node_11;
    MUX_UNSIGNED #(.width(5)) u_mux_49 (
        .y(_node_11),
        .sel(_node_10),
        .a(_T_347_5),
        .b(_node_9)
    );
    wire _node_12;
    EQ_UNSIGNED #(.width(7)) u_eq_50 (
        .y(_node_12),
        .a(7'd6),
        .b(_value__q)
    );
    wire [4:0] _node_13;
    MUX_UNSIGNED #(.width(5)) u_mux_51 (
        .y(_node_13),
        .sel(_node_12),
        .a(_T_347_6),
        .b(_node_11)
    );
    wire _node_14;
    EQ_UNSIGNED #(.width(7)) u_eq_52 (
        .y(_node_14),
        .a(7'd7),
        .b(_value__q)
    );
    wire [4:0] _node_15;
    MUX_UNSIGNED #(.width(5)) u_mux_53 (
        .y(_node_15),
        .sel(_node_14),
        .a(_T_347_7),
        .b(_node_13)
    );
    wire _node_16;
    EQ_UNSIGNED #(.width(7)) u_eq_54 (
        .y(_node_16),
        .a(7'd8),
        .b(_value__q)
    );
    wire [4:0] _node_17;
    MUX_UNSIGNED #(.width(5)) u_mux_55 (
        .y(_node_17),
        .sel(_node_16),
        .a(_T_347_8),
        .b(_node_15)
    );
    wire _node_18;
    EQ_UNSIGNED #(.width(7)) u_eq_56 (
        .y(_node_18),
        .a(7'd9),
        .b(_value__q)
    );
    wire [4:0] _node_19;
    MUX_UNSIGNED #(.width(5)) u_mux_57 (
        .y(_node_19),
        .sel(_node_18),
        .a(_T_347_9),
        .b(_node_17)
    );
    wire _node_20;
    EQ_UNSIGNED #(.width(7)) u_eq_58 (
        .y(_node_20),
        .a(7'd10),
        .b(_value__q)
    );
    wire [4:0] _node_21;
    MUX_UNSIGNED #(.width(5)) u_mux_59 (
        .y(_node_21),
        .sel(_node_20),
        .a(_T_347_10),
        .b(_node_19)
    );
    wire _node_22;
    EQ_UNSIGNED #(.width(7)) u_eq_60 (
        .y(_node_22),
        .a(7'd11),
        .b(_value__q)
    );
    wire [4:0] _node_23;
    MUX_UNSIGNED #(.width(5)) u_mux_61 (
        .y(_node_23),
        .sel(_node_22),
        .a(_T_347_11),
        .b(_node_21)
    );
    wire _node_24;
    EQ_UNSIGNED #(.width(7)) u_eq_62 (
        .y(_node_24),
        .a(7'd12),
        .b(_value__q)
    );
    wire [4:0] _node_25;
    MUX_UNSIGNED #(.width(5)) u_mux_63 (
        .y(_node_25),
        .sel(_node_24),
        .a(_T_347_12),
        .b(_node_23)
    );
    wire _node_26;
    EQ_UNSIGNED #(.width(7)) u_eq_64 (
        .y(_node_26),
        .a(7'd13),
        .b(_value__q)
    );
    wire [4:0] _node_27;
    MUX_UNSIGNED #(.width(5)) u_mux_65 (
        .y(_node_27),
        .sel(_node_26),
        .a(_T_347_13),
        .b(_node_25)
    );
    wire _node_28;
    EQ_UNSIGNED #(.width(7)) u_eq_66 (
        .y(_node_28),
        .a(7'd14),
        .b(_value__q)
    );
    wire [4:0] _node_29;
    MUX_UNSIGNED #(.width(5)) u_mux_67 (
        .y(_node_29),
        .sel(_node_28),
        .a(_T_347_14),
        .b(_node_27)
    );
    wire _node_30;
    EQ_UNSIGNED #(.width(7)) u_eq_68 (
        .y(_node_30),
        .a(7'd15),
        .b(_value__q)
    );
    wire [4:0] _node_31;
    MUX_UNSIGNED #(.width(5)) u_mux_69 (
        .y(_node_31),
        .sel(_node_30),
        .a(_T_347_15),
        .b(_node_29)
    );
    wire _node_32;
    EQ_UNSIGNED #(.width(7)) u_eq_70 (
        .y(_node_32),
        .a(7'd16),
        .b(_value__q)
    );
    wire [4:0] _node_33;
    MUX_UNSIGNED #(.width(5)) u_mux_71 (
        .y(_node_33),
        .sel(_node_32),
        .a(_T_347_16),
        .b(_node_31)
    );
    wire _node_34;
    EQ_UNSIGNED #(.width(7)) u_eq_72 (
        .y(_node_34),
        .a(7'd17),
        .b(_value__q)
    );
    wire [4:0] _node_35;
    MUX_UNSIGNED #(.width(5)) u_mux_73 (
        .y(_node_35),
        .sel(_node_34),
        .a(_T_347_17),
        .b(_node_33)
    );
    wire _node_36;
    EQ_UNSIGNED #(.width(7)) u_eq_74 (
        .y(_node_36),
        .a(7'd18),
        .b(_value__q)
    );
    wire [4:0] _node_37;
    MUX_UNSIGNED #(.width(5)) u_mux_75 (
        .y(_node_37),
        .sel(_node_36),
        .a(_T_347_18),
        .b(_node_35)
    );
    wire _node_38;
    EQ_UNSIGNED #(.width(7)) u_eq_76 (
        .y(_node_38),
        .a(7'd19),
        .b(_value__q)
    );
    wire [4:0] _node_39;
    MUX_UNSIGNED #(.width(5)) u_mux_77 (
        .y(_node_39),
        .sel(_node_38),
        .a(_T_347_19),
        .b(_node_37)
    );
    wire _node_40;
    EQ_UNSIGNED #(.width(7)) u_eq_78 (
        .y(_node_40),
        .a(7'd20),
        .b(_value__q)
    );
    wire [4:0] _node_41;
    MUX_UNSIGNED #(.width(5)) u_mux_79 (
        .y(_node_41),
        .sel(_node_40),
        .a(_T_347_20),
        .b(_node_39)
    );
    wire _node_42;
    EQ_UNSIGNED #(.width(7)) u_eq_80 (
        .y(_node_42),
        .a(7'd21),
        .b(_value__q)
    );
    wire [4:0] _node_43;
    MUX_UNSIGNED #(.width(5)) u_mux_81 (
        .y(_node_43),
        .sel(_node_42),
        .a(_T_347_21),
        .b(_node_41)
    );
    wire _node_44;
    EQ_UNSIGNED #(.width(7)) u_eq_82 (
        .y(_node_44),
        .a(7'd22),
        .b(_value__q)
    );
    wire [4:0] _node_45;
    MUX_UNSIGNED #(.width(5)) u_mux_83 (
        .y(_node_45),
        .sel(_node_44),
        .a(_T_347_22),
        .b(_node_43)
    );
    wire _node_46;
    EQ_UNSIGNED #(.width(7)) u_eq_84 (
        .y(_node_46),
        .a(7'd23),
        .b(_value__q)
    );
    wire [4:0] _node_47;
    MUX_UNSIGNED #(.width(5)) u_mux_85 (
        .y(_node_47),
        .sel(_node_46),
        .a(_T_347_23),
        .b(_node_45)
    );
    wire _node_48;
    EQ_UNSIGNED #(.width(7)) u_eq_86 (
        .y(_node_48),
        .a(7'd24),
        .b(_value__q)
    );
    wire [4:0] _node_49;
    MUX_UNSIGNED #(.width(5)) u_mux_87 (
        .y(_node_49),
        .sel(_node_48),
        .a(_T_347_24),
        .b(_node_47)
    );
    wire _node_50;
    EQ_UNSIGNED #(.width(7)) u_eq_88 (
        .y(_node_50),
        .a(7'd25),
        .b(_value__q)
    );
    wire [4:0] _node_51;
    MUX_UNSIGNED #(.width(5)) u_mux_89 (
        .y(_node_51),
        .sel(_node_50),
        .a(_T_347_25),
        .b(_node_49)
    );
    wire _node_52;
    EQ_UNSIGNED #(.width(7)) u_eq_90 (
        .y(_node_52),
        .a(7'd26),
        .b(_value__q)
    );
    wire [4:0] _node_53;
    MUX_UNSIGNED #(.width(5)) u_mux_91 (
        .y(_node_53),
        .sel(_node_52),
        .a(_T_347_26),
        .b(_node_51)
    );
    wire _node_54;
    EQ_UNSIGNED #(.width(7)) u_eq_92 (
        .y(_node_54),
        .a(7'd27),
        .b(_value__q)
    );
    wire [4:0] _node_55;
    MUX_UNSIGNED #(.width(5)) u_mux_93 (
        .y(_node_55),
        .sel(_node_54),
        .a(_T_347_27),
        .b(_node_53)
    );
    wire _node_56;
    EQ_UNSIGNED #(.width(7)) u_eq_94 (
        .y(_node_56),
        .a(7'd28),
        .b(_value__q)
    );
    wire [4:0] _node_57;
    MUX_UNSIGNED #(.width(5)) u_mux_95 (
        .y(_node_57),
        .sel(_node_56),
        .a(_T_347_28),
        .b(_node_55)
    );
    wire _node_58;
    EQ_UNSIGNED #(.width(7)) u_eq_96 (
        .y(_node_58),
        .a(7'd29),
        .b(_value__q)
    );
    wire [4:0] _node_59;
    MUX_UNSIGNED #(.width(5)) u_mux_97 (
        .y(_node_59),
        .sel(_node_58),
        .a(_T_347_29),
        .b(_node_57)
    );
    wire _node_60;
    EQ_UNSIGNED #(.width(7)) u_eq_98 (
        .y(_node_60),
        .a(7'd30),
        .b(_value__q)
    );
    wire [4:0] _node_61;
    MUX_UNSIGNED #(.width(5)) u_mux_99 (
        .y(_node_61),
        .sel(_node_60),
        .a(_T_347_30),
        .b(_node_59)
    );
    wire _node_62;
    EQ_UNSIGNED #(.width(7)) u_eq_100 (
        .y(_node_62),
        .a(7'd31),
        .b(_value__q)
    );
    wire [4:0] _node_63;
    MUX_UNSIGNED #(.width(5)) u_mux_101 (
        .y(_node_63),
        .sel(_node_62),
        .a(_T_347_31),
        .b(_node_61)
    );
    wire _node_64;
    EQ_UNSIGNED #(.width(7)) u_eq_102 (
        .y(_node_64),
        .a(7'd32),
        .b(_value__q)
    );
    wire [4:0] _node_65;
    MUX_UNSIGNED #(.width(5)) u_mux_103 (
        .y(_node_65),
        .sel(_node_64),
        .a(_T_347_32),
        .b(_node_63)
    );
    wire _node_66;
    EQ_UNSIGNED #(.width(7)) u_eq_104 (
        .y(_node_66),
        .a(7'd33),
        .b(_value__q)
    );
    wire [4:0] _node_67;
    MUX_UNSIGNED #(.width(5)) u_mux_105 (
        .y(_node_67),
        .sel(_node_66),
        .a(_T_347_33),
        .b(_node_65)
    );
    wire _node_68;
    EQ_UNSIGNED #(.width(7)) u_eq_106 (
        .y(_node_68),
        .a(7'd34),
        .b(_value__q)
    );
    wire [4:0] _node_69;
    MUX_UNSIGNED #(.width(5)) u_mux_107 (
        .y(_node_69),
        .sel(_node_68),
        .a(_T_347_34),
        .b(_node_67)
    );
    wire _node_70;
    EQ_UNSIGNED #(.width(7)) u_eq_108 (
        .y(_node_70),
        .a(7'd35),
        .b(_value__q)
    );
    wire [4:0] _node_71;
    MUX_UNSIGNED #(.width(5)) u_mux_109 (
        .y(_node_71),
        .sel(_node_70),
        .a(_T_347_35),
        .b(_node_69)
    );
    wire _node_72;
    EQ_UNSIGNED #(.width(7)) u_eq_110 (
        .y(_node_72),
        .a(7'd36),
        .b(_value__q)
    );
    wire [4:0] _node_73;
    MUX_UNSIGNED #(.width(5)) u_mux_111 (
        .y(_node_73),
        .sel(_node_72),
        .a(_T_347_36),
        .b(_node_71)
    );
    wire _node_74;
    EQ_UNSIGNED #(.width(7)) u_eq_112 (
        .y(_node_74),
        .a(7'd37),
        .b(_value__q)
    );
    wire [4:0] _node_75;
    MUX_UNSIGNED #(.width(5)) u_mux_113 (
        .y(_node_75),
        .sel(_node_74),
        .a(_T_347_37),
        .b(_node_73)
    );
    wire _node_76;
    EQ_UNSIGNED #(.width(7)) u_eq_114 (
        .y(_node_76),
        .a(7'd38),
        .b(_value__q)
    );
    wire [4:0] _node_77;
    MUX_UNSIGNED #(.width(5)) u_mux_115 (
        .y(_node_77),
        .sel(_node_76),
        .a(_T_347_38),
        .b(_node_75)
    );
    wire _node_78;
    EQ_UNSIGNED #(.width(7)) u_eq_116 (
        .y(_node_78),
        .a(7'd39),
        .b(_value__q)
    );
    wire [4:0] _node_79;
    MUX_UNSIGNED #(.width(5)) u_mux_117 (
        .y(_node_79),
        .sel(_node_78),
        .a(_T_347_39),
        .b(_node_77)
    );
    wire _node_80;
    EQ_UNSIGNED #(.width(7)) u_eq_118 (
        .y(_node_80),
        .a(7'd40),
        .b(_value__q)
    );
    wire [4:0] _node_81;
    MUX_UNSIGNED #(.width(5)) u_mux_119 (
        .y(_node_81),
        .sel(_node_80),
        .a(_T_347_40),
        .b(_node_79)
    );
    wire _node_82;
    EQ_UNSIGNED #(.width(7)) u_eq_120 (
        .y(_node_82),
        .a(7'd41),
        .b(_value__q)
    );
    wire [4:0] _node_83;
    MUX_UNSIGNED #(.width(5)) u_mux_121 (
        .y(_node_83),
        .sel(_node_82),
        .a(_T_347_41),
        .b(_node_81)
    );
    wire _node_84;
    EQ_UNSIGNED #(.width(7)) u_eq_122 (
        .y(_node_84),
        .a(7'd42),
        .b(_value__q)
    );
    wire [4:0] _node_85;
    MUX_UNSIGNED #(.width(5)) u_mux_123 (
        .y(_node_85),
        .sel(_node_84),
        .a(_T_347_42),
        .b(_node_83)
    );
    wire _node_86;
    EQ_UNSIGNED #(.width(7)) u_eq_124 (
        .y(_node_86),
        .a(7'd43),
        .b(_value__q)
    );
    wire [4:0] _node_87;
    MUX_UNSIGNED #(.width(5)) u_mux_125 (
        .y(_node_87),
        .sel(_node_86),
        .a(_T_347_43),
        .b(_node_85)
    );
    wire _node_88;
    EQ_UNSIGNED #(.width(7)) u_eq_126 (
        .y(_node_88),
        .a(7'd44),
        .b(_value__q)
    );
    wire [4:0] _node_89;
    MUX_UNSIGNED #(.width(5)) u_mux_127 (
        .y(_node_89),
        .sel(_node_88),
        .a(_T_347_44),
        .b(_node_87)
    );
    wire _node_90;
    EQ_UNSIGNED #(.width(7)) u_eq_128 (
        .y(_node_90),
        .a(7'd45),
        .b(_value__q)
    );
    wire [4:0] _node_91;
    MUX_UNSIGNED #(.width(5)) u_mux_129 (
        .y(_node_91),
        .sel(_node_90),
        .a(_T_347_45),
        .b(_node_89)
    );
    wire _node_92;
    EQ_UNSIGNED #(.width(7)) u_eq_130 (
        .y(_node_92),
        .a(7'd46),
        .b(_value__q)
    );
    wire [4:0] _node_93;
    MUX_UNSIGNED #(.width(5)) u_mux_131 (
        .y(_node_93),
        .sel(_node_92),
        .a(_T_347_46),
        .b(_node_91)
    );
    wire _node_94;
    EQ_UNSIGNED #(.width(7)) u_eq_132 (
        .y(_node_94),
        .a(7'd47),
        .b(_value__q)
    );
    wire [4:0] _node_95;
    MUX_UNSIGNED #(.width(5)) u_mux_133 (
        .y(_node_95),
        .sel(_node_94),
        .a(_T_347_47),
        .b(_node_93)
    );
    wire _node_96;
    EQ_UNSIGNED #(.width(7)) u_eq_134 (
        .y(_node_96),
        .a(7'd48),
        .b(_value__q)
    );
    wire [4:0] _node_97;
    MUX_UNSIGNED #(.width(5)) u_mux_135 (
        .y(_node_97),
        .sel(_node_96),
        .a(_T_347_48),
        .b(_node_95)
    );
    wire _node_98;
    EQ_UNSIGNED #(.width(7)) u_eq_136 (
        .y(_node_98),
        .a(7'd49),
        .b(_value__q)
    );
    wire [4:0] _node_99;
    MUX_UNSIGNED #(.width(5)) u_mux_137 (
        .y(_node_99),
        .sel(_node_98),
        .a(_T_347_49),
        .b(_node_97)
    );
    wire _node_100;
    EQ_UNSIGNED #(.width(7)) u_eq_138 (
        .y(_node_100),
        .a(7'd50),
        .b(_value__q)
    );
    wire [4:0] _node_101;
    MUX_UNSIGNED #(.width(5)) u_mux_139 (
        .y(_node_101),
        .sel(_node_100),
        .a(_T_347_50),
        .b(_node_99)
    );
    wire _node_102;
    EQ_UNSIGNED #(.width(7)) u_eq_140 (
        .y(_node_102),
        .a(7'd51),
        .b(_value__q)
    );
    wire [4:0] _node_103;
    MUX_UNSIGNED #(.width(5)) u_mux_141 (
        .y(_node_103),
        .sel(_node_102),
        .a(_T_347_51),
        .b(_node_101)
    );
    wire _node_104;
    EQ_UNSIGNED #(.width(7)) u_eq_142 (
        .y(_node_104),
        .a(7'd52),
        .b(_value__q)
    );
    wire [4:0] _node_105;
    MUX_UNSIGNED #(.width(5)) u_mux_143 (
        .y(_node_105),
        .sel(_node_104),
        .a(_T_347_52),
        .b(_node_103)
    );
    wire _node_106;
    EQ_UNSIGNED #(.width(7)) u_eq_144 (
        .y(_node_106),
        .a(7'd53),
        .b(_value__q)
    );
    wire [4:0] _node_107;
    MUX_UNSIGNED #(.width(5)) u_mux_145 (
        .y(_node_107),
        .sel(_node_106),
        .a(_T_347_53),
        .b(_node_105)
    );
    wire _node_108;
    EQ_UNSIGNED #(.width(7)) u_eq_146 (
        .y(_node_108),
        .a(7'd54),
        .b(_value__q)
    );
    wire [4:0] _node_109;
    MUX_UNSIGNED #(.width(5)) u_mux_147 (
        .y(_node_109),
        .sel(_node_108),
        .a(_T_347_54),
        .b(_node_107)
    );
    wire _node_110;
    EQ_UNSIGNED #(.width(7)) u_eq_148 (
        .y(_node_110),
        .a(7'd55),
        .b(_value__q)
    );
    wire [4:0] _node_111;
    MUX_UNSIGNED #(.width(5)) u_mux_149 (
        .y(_node_111),
        .sel(_node_110),
        .a(_T_347_55),
        .b(_node_109)
    );
    wire _node_112;
    EQ_UNSIGNED #(.width(7)) u_eq_150 (
        .y(_node_112),
        .a(7'd56),
        .b(_value__q)
    );
    wire [4:0] _node_113;
    MUX_UNSIGNED #(.width(5)) u_mux_151 (
        .y(_node_113),
        .sel(_node_112),
        .a(_T_347_56),
        .b(_node_111)
    );
    wire _node_114;
    EQ_UNSIGNED #(.width(7)) u_eq_152 (
        .y(_node_114),
        .a(7'd57),
        .b(_value__q)
    );
    wire [4:0] _node_115;
    MUX_UNSIGNED #(.width(5)) u_mux_153 (
        .y(_node_115),
        .sel(_node_114),
        .a(_T_347_57),
        .b(_node_113)
    );
    wire _node_116;
    EQ_UNSIGNED #(.width(7)) u_eq_154 (
        .y(_node_116),
        .a(7'd58),
        .b(_value__q)
    );
    wire [4:0] _node_117;
    MUX_UNSIGNED #(.width(5)) u_mux_155 (
        .y(_node_117),
        .sel(_node_116),
        .a(_T_347_58),
        .b(_node_115)
    );
    wire _node_118;
    EQ_UNSIGNED #(.width(7)) u_eq_156 (
        .y(_node_118),
        .a(7'd59),
        .b(_value__q)
    );
    wire [4:0] _node_119;
    MUX_UNSIGNED #(.width(5)) u_mux_157 (
        .y(_node_119),
        .sel(_node_118),
        .a(_T_347_59),
        .b(_node_117)
    );
    wire _node_120;
    EQ_UNSIGNED #(.width(7)) u_eq_158 (
        .y(_node_120),
        .a(7'd60),
        .b(_value__q)
    );
    wire [4:0] _node_121;
    MUX_UNSIGNED #(.width(5)) u_mux_159 (
        .y(_node_121),
        .sel(_node_120),
        .a(_T_347_60),
        .b(_node_119)
    );
    wire _node_122;
    EQ_UNSIGNED #(.width(7)) u_eq_160 (
        .y(_node_122),
        .a(7'd61),
        .b(_value__q)
    );
    wire [4:0] _node_123;
    MUX_UNSIGNED #(.width(5)) u_mux_161 (
        .y(_node_123),
        .sel(_node_122),
        .a(_T_347_61),
        .b(_node_121)
    );
    wire _node_124;
    EQ_UNSIGNED #(.width(7)) u_eq_162 (
        .y(_node_124),
        .a(7'd62),
        .b(_value__q)
    );
    wire [4:0] _node_125;
    MUX_UNSIGNED #(.width(5)) u_mux_163 (
        .y(_node_125),
        .sel(_node_124),
        .a(_T_347_62),
        .b(_node_123)
    );
    wire _node_126;
    EQ_UNSIGNED #(.width(7)) u_eq_164 (
        .y(_node_126),
        .a(7'd63),
        .b(_value__q)
    );
    wire [4:0] _node_127;
    MUX_UNSIGNED #(.width(5)) u_mux_165 (
        .y(_node_127),
        .sel(_node_126),
        .a(_T_347_63),
        .b(_node_125)
    );
    wire _node_128;
    EQ_UNSIGNED #(.width(7)) u_eq_166 (
        .y(_node_128),
        .a(7'd64),
        .b(_value__q)
    );
    wire [4:0] _node_129;
    MUX_UNSIGNED #(.width(5)) u_mux_167 (
        .y(_node_129),
        .sel(_node_128),
        .a(_T_347_64),
        .b(_node_127)
    );
    wire _node_130;
    EQ_UNSIGNED #(.width(7)) u_eq_168 (
        .y(_node_130),
        .a(7'd65),
        .b(_value__q)
    );
    wire [4:0] _node_131;
    MUX_UNSIGNED #(.width(5)) u_mux_169 (
        .y(_node_131),
        .sel(_node_130),
        .a(_T_347_65),
        .b(_node_129)
    );
    wire _node_132;
    EQ_UNSIGNED #(.width(7)) u_eq_170 (
        .y(_node_132),
        .a(7'd66),
        .b(_value__q)
    );
    wire [4:0] _node_133;
    MUX_UNSIGNED #(.width(5)) u_mux_171 (
        .y(_node_133),
        .sel(_node_132),
        .a(_T_347_66),
        .b(_node_131)
    );
    wire _node_134;
    EQ_UNSIGNED #(.width(7)) u_eq_172 (
        .y(_node_134),
        .a(7'd67),
        .b(_value__q)
    );
    wire [4:0] _node_135;
    MUX_UNSIGNED #(.width(5)) u_mux_173 (
        .y(_node_135),
        .sel(_node_134),
        .a(_T_347_67),
        .b(_node_133)
    );
    wire _node_136;
    EQ_UNSIGNED #(.width(7)) u_eq_174 (
        .y(_node_136),
        .a(7'd68),
        .b(_value__q)
    );
    wire [4:0] _node_137;
    MUX_UNSIGNED #(.width(5)) u_mux_175 (
        .y(_node_137),
        .sel(_node_136),
        .a(_T_347_68),
        .b(_node_135)
    );
    wire _node_138;
    EQ_UNSIGNED #(.width(7)) u_eq_176 (
        .y(_node_138),
        .a(7'd69),
        .b(_value__q)
    );
    wire [4:0] _node_139;
    MUX_UNSIGNED #(.width(5)) u_mux_177 (
        .y(_node_139),
        .sel(_node_138),
        .a(_T_347_69),
        .b(_node_137)
    );
    wire _node_140;
    EQ_UNSIGNED #(.width(7)) u_eq_178 (
        .y(_node_140),
        .a(7'd70),
        .b(_value__q)
    );
    wire [4:0] _node_141;
    MUX_UNSIGNED #(.width(5)) u_mux_179 (
        .y(_node_141),
        .sel(_node_140),
        .a(_T_347_70),
        .b(_node_139)
    );
    wire _node_142;
    EQ_UNSIGNED #(.width(7)) u_eq_180 (
        .y(_node_142),
        .a(7'd71),
        .b(_value__q)
    );
    wire [4:0] _node_143;
    MUX_UNSIGNED #(.width(5)) u_mux_181 (
        .y(_node_143),
        .sel(_node_142),
        .a(_T_347_71),
        .b(_node_141)
    );
    wire _node_144;
    EQ_UNSIGNED #(.width(7)) u_eq_182 (
        .y(_node_144),
        .a(7'd72),
        .b(_value__q)
    );
    wire [4:0] _node_145;
    MUX_UNSIGNED #(.width(5)) u_mux_183 (
        .y(_node_145),
        .sel(_node_144),
        .a(_T_347_72),
        .b(_node_143)
    );
    wire _node_146;
    EQ_UNSIGNED #(.width(7)) u_eq_184 (
        .y(_node_146),
        .a(7'd73),
        .b(_value__q)
    );
    wire [4:0] _node_147;
    MUX_UNSIGNED #(.width(5)) u_mux_185 (
        .y(_node_147),
        .sel(_node_146),
        .a(_T_347_73),
        .b(_node_145)
    );
    wire _node_148;
    EQ_UNSIGNED #(.width(7)) u_eq_186 (
        .y(_node_148),
        .a(7'd74),
        .b(_value__q)
    );
    wire [4:0] _node_149;
    MUX_UNSIGNED #(.width(5)) u_mux_187 (
        .y(_node_149),
        .sel(_node_148),
        .a(_T_347_74),
        .b(_node_147)
    );
    wire _node_150;
    EQ_UNSIGNED #(.width(7)) u_eq_188 (
        .y(_node_150),
        .a(7'd75),
        .b(_value__q)
    );
    wire [4:0] _node_151;
    MUX_UNSIGNED #(.width(5)) u_mux_189 (
        .y(_node_151),
        .sel(_node_150),
        .a(_T_347_75),
        .b(_node_149)
    );
    wire _node_152;
    EQ_UNSIGNED #(.width(7)) u_eq_190 (
        .y(_node_152),
        .a(7'd76),
        .b(_value__q)
    );
    wire [4:0] _node_153;
    MUX_UNSIGNED #(.width(5)) u_mux_191 (
        .y(_node_153),
        .sel(_node_152),
        .a(_T_347_76),
        .b(_node_151)
    );
    wire _node_154;
    EQ_UNSIGNED #(.width(7)) u_eq_192 (
        .y(_node_154),
        .a(7'd77),
        .b(_value__q)
    );
    wire [4:0] _node_155;
    MUX_UNSIGNED #(.width(5)) u_mux_193 (
        .y(_node_155),
        .sel(_node_154),
        .a(_T_347_77),
        .b(_node_153)
    );
    wire _node_156;
    EQ_UNSIGNED #(.width(7)) u_eq_194 (
        .y(_node_156),
        .a(7'd78),
        .b(_value__q)
    );
    wire [4:0] _node_157;
    MUX_UNSIGNED #(.width(5)) u_mux_195 (
        .y(_node_157),
        .sel(_node_156),
        .a(_T_347_78),
        .b(_node_155)
    );
    wire _node_158;
    EQ_UNSIGNED #(.width(7)) u_eq_196 (
        .y(_node_158),
        .a(7'd79),
        .b(_value__q)
    );
    wire [4:0] _node_159;
    MUX_UNSIGNED #(.width(5)) u_mux_197 (
        .y(_node_159),
        .sel(_node_158),
        .a(_T_347_79),
        .b(_node_157)
    );
    wire _node_160;
    EQ_UNSIGNED #(.width(7)) u_eq_198 (
        .y(_node_160),
        .a(7'd80),
        .b(_value__q)
    );
    wire [4:0] _node_161;
    MUX_UNSIGNED #(.width(5)) u_mux_199 (
        .y(_node_161),
        .sel(_node_160),
        .a(_T_347_80),
        .b(_node_159)
    );
    wire _node_162;
    EQ_UNSIGNED #(.width(7)) u_eq_200 (
        .y(_node_162),
        .a(7'd81),
        .b(_value__q)
    );
    wire [4:0] _node_163;
    MUX_UNSIGNED #(.width(5)) u_mux_201 (
        .y(_node_163),
        .sel(_node_162),
        .a(_T_347_81),
        .b(_node_161)
    );
    wire _node_164;
    EQ_UNSIGNED #(.width(7)) u_eq_202 (
        .y(_node_164),
        .a(7'd82),
        .b(_value__q)
    );
    wire [4:0] _node_165;
    MUX_UNSIGNED #(.width(5)) u_mux_203 (
        .y(_node_165),
        .sel(_node_164),
        .a(_T_347_82),
        .b(_node_163)
    );
    wire _node_166;
    EQ_UNSIGNED #(.width(7)) u_eq_204 (
        .y(_node_166),
        .a(7'd83),
        .b(_value__q)
    );
    wire [4:0] _node_167;
    MUX_UNSIGNED #(.width(5)) u_mux_205 (
        .y(_node_167),
        .sel(_node_166),
        .a(_T_347_83),
        .b(_node_165)
    );
    wire _node_168;
    EQ_UNSIGNED #(.width(7)) u_eq_206 (
        .y(_node_168),
        .a(7'd84),
        .b(_value__q)
    );
    wire [4:0] _node_169;
    MUX_UNSIGNED #(.width(5)) u_mux_207 (
        .y(_node_169),
        .sel(_node_168),
        .a(_T_347_84),
        .b(_node_167)
    );
    wire _node_170;
    EQ_UNSIGNED #(.width(7)) u_eq_208 (
        .y(_node_170),
        .a(7'd85),
        .b(_value__q)
    );
    wire [4:0] _node_171;
    MUX_UNSIGNED #(.width(5)) u_mux_209 (
        .y(_node_171),
        .sel(_node_170),
        .a(_T_347_85),
        .b(_node_169)
    );
    wire _node_172;
    EQ_UNSIGNED #(.width(7)) u_eq_210 (
        .y(_node_172),
        .a(7'd86),
        .b(_value__q)
    );
    wire [4:0] _node_173;
    MUX_UNSIGNED #(.width(5)) u_mux_211 (
        .y(_node_173),
        .sel(_node_172),
        .a(_T_347_86),
        .b(_node_171)
    );
    wire _node_174;
    EQ_UNSIGNED #(.width(7)) u_eq_212 (
        .y(_node_174),
        .a(7'd87),
        .b(_value__q)
    );
    wire [4:0] _node_175;
    MUX_UNSIGNED #(.width(5)) u_mux_213 (
        .y(_node_175),
        .sel(_node_174),
        .a(_T_347_87),
        .b(_node_173)
    );
    wire _node_176;
    EQ_UNSIGNED #(.width(7)) u_eq_214 (
        .y(_node_176),
        .a(7'd88),
        .b(_value__q)
    );
    wire [4:0] _node_177;
    MUX_UNSIGNED #(.width(5)) u_mux_215 (
        .y(_node_177),
        .sel(_node_176),
        .a(_T_347_88),
        .b(_node_175)
    );
    wire _node_178;
    EQ_UNSIGNED #(.width(7)) u_eq_216 (
        .y(_node_178),
        .a(7'd89),
        .b(_value__q)
    );
    wire [4:0] _node_179;
    MUX_UNSIGNED #(.width(5)) u_mux_217 (
        .y(_node_179),
        .sel(_node_178),
        .a(_T_347_89),
        .b(_node_177)
    );
    wire _node_180;
    EQ_UNSIGNED #(.width(7)) u_eq_218 (
        .y(_node_180),
        .a(7'd90),
        .b(_value__q)
    );
    wire [4:0] _node_181;
    MUX_UNSIGNED #(.width(5)) u_mux_219 (
        .y(_node_181),
        .sel(_node_180),
        .a(_T_347_90),
        .b(_node_179)
    );
    wire _node_182;
    EQ_UNSIGNED #(.width(7)) u_eq_220 (
        .y(_node_182),
        .a(7'd91),
        .b(_value__q)
    );
    wire [4:0] _node_183;
    MUX_UNSIGNED #(.width(5)) u_mux_221 (
        .y(_node_183),
        .sel(_node_182),
        .a(_T_347_91),
        .b(_node_181)
    );
    wire _node_184;
    EQ_UNSIGNED #(.width(7)) u_eq_222 (
        .y(_node_184),
        .a(7'd92),
        .b(_value__q)
    );
    wire [4:0] _node_185;
    MUX_UNSIGNED #(.width(5)) u_mux_223 (
        .y(_node_185),
        .sel(_node_184),
        .a(_T_347_92),
        .b(_node_183)
    );
    wire _node_186;
    EQ_UNSIGNED #(.width(7)) u_eq_224 (
        .y(_node_186),
        .a(7'd93),
        .b(_value__q)
    );
    wire [4:0] _node_187;
    MUX_UNSIGNED #(.width(5)) u_mux_225 (
        .y(_node_187),
        .sel(_node_186),
        .a(_T_347_93),
        .b(_node_185)
    );
    wire _node_188;
    EQ_UNSIGNED #(.width(7)) u_eq_226 (
        .y(_node_188),
        .a(7'd94),
        .b(_value__q)
    );
    wire [4:0] _node_189;
    MUX_UNSIGNED #(.width(5)) u_mux_227 (
        .y(_node_189),
        .sel(_node_188),
        .a(_T_347_94),
        .b(_node_187)
    );
    wire _node_190;
    EQ_UNSIGNED #(.width(7)) u_eq_228 (
        .y(_node_190),
        .a(7'd95),
        .b(_value__q)
    );
    wire [4:0] _node_191;
    MUX_UNSIGNED #(.width(5)) u_mux_229 (
        .y(_node_191),
        .sel(_node_190),
        .a(_T_347_95),
        .b(_node_189)
    );
    wire _node_192;
    EQ_UNSIGNED #(.width(7)) u_eq_230 (
        .y(_node_192),
        .a(7'd96),
        .b(_value__q)
    );
    wire [4:0] _node_193;
    MUX_UNSIGNED #(.width(5)) u_mux_231 (
        .y(_node_193),
        .sel(_node_192),
        .a(_T_347_96),
        .b(_node_191)
    );
    wire _node_194;
    EQ_UNSIGNED #(.width(7)) u_eq_232 (
        .y(_node_194),
        .a(7'd97),
        .b(_value__q)
    );
    wire [4:0] _node_195;
    MUX_UNSIGNED #(.width(5)) u_mux_233 (
        .y(_node_195),
        .sel(_node_194),
        .a(_T_347_97),
        .b(_node_193)
    );
    wire _node_196;
    EQ_UNSIGNED #(.width(7)) u_eq_234 (
        .y(_node_196),
        .a(7'd98),
        .b(_value__q)
    );
    wire [4:0] _node_197;
    MUX_UNSIGNED #(.width(5)) u_mux_235 (
        .y(_node_197),
        .sel(_node_196),
        .a(_T_347_98),
        .b(_node_195)
    );
    wire _node_198;
    EQ_UNSIGNED #(.width(7)) u_eq_236 (
        .y(_node_198),
        .a(7'd99),
        .b(_value__q)
    );
    wire [4:0] _node_199;
    MUX_UNSIGNED #(.width(5)) u_mux_237 (
        .y(_node_199),
        .sel(_node_198),
        .a(_T_347_99),
        .b(_node_197)
    );
    wire _node_200;
    EQ_UNSIGNED #(.width(7)) u_eq_238 (
        .y(_node_200),
        .a(7'd100),
        .b(_value__q)
    );
    wire [4:0] _node_201;
    MUX_UNSIGNED #(.width(5)) u_mux_239 (
        .y(_node_201),
        .sel(_node_200),
        .a(_T_347_100),
        .b(_node_199)
    );
    wire _node_202;
    EQ_UNSIGNED #(.width(7)) u_eq_240 (
        .y(_node_202),
        .a(7'd101),
        .b(_value__q)
    );
    wire [4:0] _node_203;
    MUX_UNSIGNED #(.width(5)) u_mux_241 (
        .y(_node_203),
        .sel(_node_202),
        .a(_T_347_101),
        .b(_node_201)
    );
    wire [6:0] _T_454;
    BITS #(.width(9), .high(6), .low(0)) bits_242 (
        .y(_T_454),
        .in(__T_4__q)
    );
    wire _node_204;
    EQ_UNSIGNED #(.width(7)) u_eq_243 (
        .y(_node_204),
        .a(7'd0),
        .b(_T_454)
    );
    wire _node_205;
    assign _node_205 = _T_136_0;
    wire _node_206;
    EQ_UNSIGNED #(.width(7)) u_eq_244 (
        .y(_node_206),
        .a(7'd1),
        .b(_T_454)
    );
    wire _node_207;
    MUX_UNSIGNED #(.width(1)) u_mux_245 (
        .y(_node_207),
        .sel(_node_206),
        .a(_T_136_1),
        .b(_node_205)
    );
    wire _node_208;
    EQ_UNSIGNED #(.width(7)) u_eq_246 (
        .y(_node_208),
        .a(7'd2),
        .b(_T_454)
    );
    wire _node_209;
    MUX_UNSIGNED #(.width(1)) u_mux_247 (
        .y(_node_209),
        .sel(_node_208),
        .a(_T_136_2),
        .b(_node_207)
    );
    wire _node_210;
    EQ_UNSIGNED #(.width(7)) u_eq_248 (
        .y(_node_210),
        .a(7'd3),
        .b(_T_454)
    );
    wire _node_211;
    MUX_UNSIGNED #(.width(1)) u_mux_249 (
        .y(_node_211),
        .sel(_node_210),
        .a(_T_136_3),
        .b(_node_209)
    );
    wire _node_212;
    EQ_UNSIGNED #(.width(7)) u_eq_250 (
        .y(_node_212),
        .a(7'd4),
        .b(_T_454)
    );
    wire _node_213;
    MUX_UNSIGNED #(.width(1)) u_mux_251 (
        .y(_node_213),
        .sel(_node_212),
        .a(_T_136_4),
        .b(_node_211)
    );
    wire _node_214;
    EQ_UNSIGNED #(.width(7)) u_eq_252 (
        .y(_node_214),
        .a(7'd5),
        .b(_T_454)
    );
    wire _node_215;
    MUX_UNSIGNED #(.width(1)) u_mux_253 (
        .y(_node_215),
        .sel(_node_214),
        .a(_T_136_5),
        .b(_node_213)
    );
    wire _node_216;
    EQ_UNSIGNED #(.width(7)) u_eq_254 (
        .y(_node_216),
        .a(7'd6),
        .b(_T_454)
    );
    wire _node_217;
    MUX_UNSIGNED #(.width(1)) u_mux_255 (
        .y(_node_217),
        .sel(_node_216),
        .a(_T_136_6),
        .b(_node_215)
    );
    wire _node_218;
    EQ_UNSIGNED #(.width(7)) u_eq_256 (
        .y(_node_218),
        .a(7'd7),
        .b(_T_454)
    );
    wire _node_219;
    MUX_UNSIGNED #(.width(1)) u_mux_257 (
        .y(_node_219),
        .sel(_node_218),
        .a(_T_136_7),
        .b(_node_217)
    );
    wire _node_220;
    EQ_UNSIGNED #(.width(7)) u_eq_258 (
        .y(_node_220),
        .a(7'd8),
        .b(_T_454)
    );
    wire _node_221;
    MUX_UNSIGNED #(.width(1)) u_mux_259 (
        .y(_node_221),
        .sel(_node_220),
        .a(_T_136_8),
        .b(_node_219)
    );
    wire _node_222;
    EQ_UNSIGNED #(.width(7)) u_eq_260 (
        .y(_node_222),
        .a(7'd9),
        .b(_T_454)
    );
    wire _node_223;
    MUX_UNSIGNED #(.width(1)) u_mux_261 (
        .y(_node_223),
        .sel(_node_222),
        .a(_T_136_9),
        .b(_node_221)
    );
    wire _node_224;
    EQ_UNSIGNED #(.width(7)) u_eq_262 (
        .y(_node_224),
        .a(7'd10),
        .b(_T_454)
    );
    wire _node_225;
    MUX_UNSIGNED #(.width(1)) u_mux_263 (
        .y(_node_225),
        .sel(_node_224),
        .a(_T_136_10),
        .b(_node_223)
    );
    wire _node_226;
    EQ_UNSIGNED #(.width(7)) u_eq_264 (
        .y(_node_226),
        .a(7'd11),
        .b(_T_454)
    );
    wire _node_227;
    MUX_UNSIGNED #(.width(1)) u_mux_265 (
        .y(_node_227),
        .sel(_node_226),
        .a(_T_136_11),
        .b(_node_225)
    );
    wire _node_228;
    EQ_UNSIGNED #(.width(7)) u_eq_266 (
        .y(_node_228),
        .a(7'd12),
        .b(_T_454)
    );
    wire _node_229;
    MUX_UNSIGNED #(.width(1)) u_mux_267 (
        .y(_node_229),
        .sel(_node_228),
        .a(_T_136_12),
        .b(_node_227)
    );
    wire _node_230;
    EQ_UNSIGNED #(.width(7)) u_eq_268 (
        .y(_node_230),
        .a(7'd13),
        .b(_T_454)
    );
    wire _node_231;
    MUX_UNSIGNED #(.width(1)) u_mux_269 (
        .y(_node_231),
        .sel(_node_230),
        .a(_T_136_13),
        .b(_node_229)
    );
    wire _node_232;
    EQ_UNSIGNED #(.width(7)) u_eq_270 (
        .y(_node_232),
        .a(7'd14),
        .b(_T_454)
    );
    wire _node_233;
    MUX_UNSIGNED #(.width(1)) u_mux_271 (
        .y(_node_233),
        .sel(_node_232),
        .a(_T_136_14),
        .b(_node_231)
    );
    wire _node_234;
    EQ_UNSIGNED #(.width(7)) u_eq_272 (
        .y(_node_234),
        .a(7'd15),
        .b(_T_454)
    );
    wire _node_235;
    MUX_UNSIGNED #(.width(1)) u_mux_273 (
        .y(_node_235),
        .sel(_node_234),
        .a(_T_136_15),
        .b(_node_233)
    );
    wire _node_236;
    EQ_UNSIGNED #(.width(7)) u_eq_274 (
        .y(_node_236),
        .a(7'd16),
        .b(_T_454)
    );
    wire _node_237;
    MUX_UNSIGNED #(.width(1)) u_mux_275 (
        .y(_node_237),
        .sel(_node_236),
        .a(_T_136_16),
        .b(_node_235)
    );
    wire _node_238;
    EQ_UNSIGNED #(.width(7)) u_eq_276 (
        .y(_node_238),
        .a(7'd17),
        .b(_T_454)
    );
    wire _node_239;
    MUX_UNSIGNED #(.width(1)) u_mux_277 (
        .y(_node_239),
        .sel(_node_238),
        .a(_T_136_17),
        .b(_node_237)
    );
    wire _node_240;
    EQ_UNSIGNED #(.width(7)) u_eq_278 (
        .y(_node_240),
        .a(7'd18),
        .b(_T_454)
    );
    wire _node_241;
    MUX_UNSIGNED #(.width(1)) u_mux_279 (
        .y(_node_241),
        .sel(_node_240),
        .a(_T_136_18),
        .b(_node_239)
    );
    wire _node_242;
    EQ_UNSIGNED #(.width(7)) u_eq_280 (
        .y(_node_242),
        .a(7'd19),
        .b(_T_454)
    );
    wire _node_243;
    MUX_UNSIGNED #(.width(1)) u_mux_281 (
        .y(_node_243),
        .sel(_node_242),
        .a(_T_136_19),
        .b(_node_241)
    );
    wire _node_244;
    EQ_UNSIGNED #(.width(7)) u_eq_282 (
        .y(_node_244),
        .a(7'd20),
        .b(_T_454)
    );
    wire _node_245;
    MUX_UNSIGNED #(.width(1)) u_mux_283 (
        .y(_node_245),
        .sel(_node_244),
        .a(_T_136_20),
        .b(_node_243)
    );
    wire _node_246;
    EQ_UNSIGNED #(.width(7)) u_eq_284 (
        .y(_node_246),
        .a(7'd21),
        .b(_T_454)
    );
    wire _node_247;
    MUX_UNSIGNED #(.width(1)) u_mux_285 (
        .y(_node_247),
        .sel(_node_246),
        .a(_T_136_21),
        .b(_node_245)
    );
    wire _node_248;
    EQ_UNSIGNED #(.width(7)) u_eq_286 (
        .y(_node_248),
        .a(7'd22),
        .b(_T_454)
    );
    wire _node_249;
    MUX_UNSIGNED #(.width(1)) u_mux_287 (
        .y(_node_249),
        .sel(_node_248),
        .a(_T_136_22),
        .b(_node_247)
    );
    wire _node_250;
    EQ_UNSIGNED #(.width(7)) u_eq_288 (
        .y(_node_250),
        .a(7'd23),
        .b(_T_454)
    );
    wire _node_251;
    MUX_UNSIGNED #(.width(1)) u_mux_289 (
        .y(_node_251),
        .sel(_node_250),
        .a(_T_136_23),
        .b(_node_249)
    );
    wire _node_252;
    EQ_UNSIGNED #(.width(7)) u_eq_290 (
        .y(_node_252),
        .a(7'd24),
        .b(_T_454)
    );
    wire _node_253;
    MUX_UNSIGNED #(.width(1)) u_mux_291 (
        .y(_node_253),
        .sel(_node_252),
        .a(_T_136_24),
        .b(_node_251)
    );
    wire _node_254;
    EQ_UNSIGNED #(.width(7)) u_eq_292 (
        .y(_node_254),
        .a(7'd25),
        .b(_T_454)
    );
    wire _node_255;
    MUX_UNSIGNED #(.width(1)) u_mux_293 (
        .y(_node_255),
        .sel(_node_254),
        .a(_T_136_25),
        .b(_node_253)
    );
    wire _node_256;
    EQ_UNSIGNED #(.width(7)) u_eq_294 (
        .y(_node_256),
        .a(7'd26),
        .b(_T_454)
    );
    wire _node_257;
    MUX_UNSIGNED #(.width(1)) u_mux_295 (
        .y(_node_257),
        .sel(_node_256),
        .a(_T_136_26),
        .b(_node_255)
    );
    wire _node_258;
    EQ_UNSIGNED #(.width(7)) u_eq_296 (
        .y(_node_258),
        .a(7'd27),
        .b(_T_454)
    );
    wire _node_259;
    MUX_UNSIGNED #(.width(1)) u_mux_297 (
        .y(_node_259),
        .sel(_node_258),
        .a(_T_136_27),
        .b(_node_257)
    );
    wire _node_260;
    EQ_UNSIGNED #(.width(7)) u_eq_298 (
        .y(_node_260),
        .a(7'd28),
        .b(_T_454)
    );
    wire _node_261;
    MUX_UNSIGNED #(.width(1)) u_mux_299 (
        .y(_node_261),
        .sel(_node_260),
        .a(_T_136_28),
        .b(_node_259)
    );
    wire _node_262;
    EQ_UNSIGNED #(.width(7)) u_eq_300 (
        .y(_node_262),
        .a(7'd29),
        .b(_T_454)
    );
    wire _node_263;
    MUX_UNSIGNED #(.width(1)) u_mux_301 (
        .y(_node_263),
        .sel(_node_262),
        .a(_T_136_29),
        .b(_node_261)
    );
    wire _node_264;
    EQ_UNSIGNED #(.width(7)) u_eq_302 (
        .y(_node_264),
        .a(7'd30),
        .b(_T_454)
    );
    wire _node_265;
    MUX_UNSIGNED #(.width(1)) u_mux_303 (
        .y(_node_265),
        .sel(_node_264),
        .a(_T_136_30),
        .b(_node_263)
    );
    wire _node_266;
    EQ_UNSIGNED #(.width(7)) u_eq_304 (
        .y(_node_266),
        .a(7'd31),
        .b(_T_454)
    );
    wire _node_267;
    MUX_UNSIGNED #(.width(1)) u_mux_305 (
        .y(_node_267),
        .sel(_node_266),
        .a(_T_136_31),
        .b(_node_265)
    );
    wire _node_268;
    EQ_UNSIGNED #(.width(7)) u_eq_306 (
        .y(_node_268),
        .a(7'd32),
        .b(_T_454)
    );
    wire _node_269;
    MUX_UNSIGNED #(.width(1)) u_mux_307 (
        .y(_node_269),
        .sel(_node_268),
        .a(_T_136_32),
        .b(_node_267)
    );
    wire _node_270;
    EQ_UNSIGNED #(.width(7)) u_eq_308 (
        .y(_node_270),
        .a(7'd33),
        .b(_T_454)
    );
    wire _node_271;
    MUX_UNSIGNED #(.width(1)) u_mux_309 (
        .y(_node_271),
        .sel(_node_270),
        .a(_T_136_33),
        .b(_node_269)
    );
    wire _node_272;
    EQ_UNSIGNED #(.width(7)) u_eq_310 (
        .y(_node_272),
        .a(7'd34),
        .b(_T_454)
    );
    wire _node_273;
    MUX_UNSIGNED #(.width(1)) u_mux_311 (
        .y(_node_273),
        .sel(_node_272),
        .a(_T_136_34),
        .b(_node_271)
    );
    wire _node_274;
    EQ_UNSIGNED #(.width(7)) u_eq_312 (
        .y(_node_274),
        .a(7'd35),
        .b(_T_454)
    );
    wire _node_275;
    MUX_UNSIGNED #(.width(1)) u_mux_313 (
        .y(_node_275),
        .sel(_node_274),
        .a(_T_136_35),
        .b(_node_273)
    );
    wire _node_276;
    EQ_UNSIGNED #(.width(7)) u_eq_314 (
        .y(_node_276),
        .a(7'd36),
        .b(_T_454)
    );
    wire _node_277;
    MUX_UNSIGNED #(.width(1)) u_mux_315 (
        .y(_node_277),
        .sel(_node_276),
        .a(_T_136_36),
        .b(_node_275)
    );
    wire _node_278;
    EQ_UNSIGNED #(.width(7)) u_eq_316 (
        .y(_node_278),
        .a(7'd37),
        .b(_T_454)
    );
    wire _node_279;
    MUX_UNSIGNED #(.width(1)) u_mux_317 (
        .y(_node_279),
        .sel(_node_278),
        .a(_T_136_37),
        .b(_node_277)
    );
    wire _node_280;
    EQ_UNSIGNED #(.width(7)) u_eq_318 (
        .y(_node_280),
        .a(7'd38),
        .b(_T_454)
    );
    wire _node_281;
    MUX_UNSIGNED #(.width(1)) u_mux_319 (
        .y(_node_281),
        .sel(_node_280),
        .a(_T_136_38),
        .b(_node_279)
    );
    wire _node_282;
    EQ_UNSIGNED #(.width(7)) u_eq_320 (
        .y(_node_282),
        .a(7'd39),
        .b(_T_454)
    );
    wire _node_283;
    MUX_UNSIGNED #(.width(1)) u_mux_321 (
        .y(_node_283),
        .sel(_node_282),
        .a(_T_136_39),
        .b(_node_281)
    );
    wire _node_284;
    EQ_UNSIGNED #(.width(7)) u_eq_322 (
        .y(_node_284),
        .a(7'd40),
        .b(_T_454)
    );
    wire _node_285;
    MUX_UNSIGNED #(.width(1)) u_mux_323 (
        .y(_node_285),
        .sel(_node_284),
        .a(_T_136_40),
        .b(_node_283)
    );
    wire _node_286;
    EQ_UNSIGNED #(.width(7)) u_eq_324 (
        .y(_node_286),
        .a(7'd41),
        .b(_T_454)
    );
    wire _node_287;
    MUX_UNSIGNED #(.width(1)) u_mux_325 (
        .y(_node_287),
        .sel(_node_286),
        .a(_T_136_41),
        .b(_node_285)
    );
    wire _node_288;
    EQ_UNSIGNED #(.width(7)) u_eq_326 (
        .y(_node_288),
        .a(7'd42),
        .b(_T_454)
    );
    wire _node_289;
    MUX_UNSIGNED #(.width(1)) u_mux_327 (
        .y(_node_289),
        .sel(_node_288),
        .a(_T_136_42),
        .b(_node_287)
    );
    wire _node_290;
    EQ_UNSIGNED #(.width(7)) u_eq_328 (
        .y(_node_290),
        .a(7'd43),
        .b(_T_454)
    );
    wire _node_291;
    MUX_UNSIGNED #(.width(1)) u_mux_329 (
        .y(_node_291),
        .sel(_node_290),
        .a(_T_136_43),
        .b(_node_289)
    );
    wire _node_292;
    EQ_UNSIGNED #(.width(7)) u_eq_330 (
        .y(_node_292),
        .a(7'd44),
        .b(_T_454)
    );
    wire _node_293;
    MUX_UNSIGNED #(.width(1)) u_mux_331 (
        .y(_node_293),
        .sel(_node_292),
        .a(_T_136_44),
        .b(_node_291)
    );
    wire _node_294;
    EQ_UNSIGNED #(.width(7)) u_eq_332 (
        .y(_node_294),
        .a(7'd45),
        .b(_T_454)
    );
    wire _node_295;
    MUX_UNSIGNED #(.width(1)) u_mux_333 (
        .y(_node_295),
        .sel(_node_294),
        .a(_T_136_45),
        .b(_node_293)
    );
    wire _node_296;
    EQ_UNSIGNED #(.width(7)) u_eq_334 (
        .y(_node_296),
        .a(7'd46),
        .b(_T_454)
    );
    wire _node_297;
    MUX_UNSIGNED #(.width(1)) u_mux_335 (
        .y(_node_297),
        .sel(_node_296),
        .a(_T_136_46),
        .b(_node_295)
    );
    wire _node_298;
    EQ_UNSIGNED #(.width(7)) u_eq_336 (
        .y(_node_298),
        .a(7'd47),
        .b(_T_454)
    );
    wire _node_299;
    MUX_UNSIGNED #(.width(1)) u_mux_337 (
        .y(_node_299),
        .sel(_node_298),
        .a(_T_136_47),
        .b(_node_297)
    );
    wire _node_300;
    EQ_UNSIGNED #(.width(7)) u_eq_338 (
        .y(_node_300),
        .a(7'd48),
        .b(_T_454)
    );
    wire _node_301;
    MUX_UNSIGNED #(.width(1)) u_mux_339 (
        .y(_node_301),
        .sel(_node_300),
        .a(_T_136_48),
        .b(_node_299)
    );
    wire _node_302;
    EQ_UNSIGNED #(.width(7)) u_eq_340 (
        .y(_node_302),
        .a(7'd49),
        .b(_T_454)
    );
    wire _node_303;
    MUX_UNSIGNED #(.width(1)) u_mux_341 (
        .y(_node_303),
        .sel(_node_302),
        .a(_T_136_49),
        .b(_node_301)
    );
    wire _node_304;
    EQ_UNSIGNED #(.width(7)) u_eq_342 (
        .y(_node_304),
        .a(7'd50),
        .b(_T_454)
    );
    wire _node_305;
    MUX_UNSIGNED #(.width(1)) u_mux_343 (
        .y(_node_305),
        .sel(_node_304),
        .a(_T_136_50),
        .b(_node_303)
    );
    wire _node_306;
    EQ_UNSIGNED #(.width(7)) u_eq_344 (
        .y(_node_306),
        .a(7'd51),
        .b(_T_454)
    );
    wire _node_307;
    MUX_UNSIGNED #(.width(1)) u_mux_345 (
        .y(_node_307),
        .sel(_node_306),
        .a(_T_136_51),
        .b(_node_305)
    );
    wire _node_308;
    EQ_UNSIGNED #(.width(7)) u_eq_346 (
        .y(_node_308),
        .a(7'd52),
        .b(_T_454)
    );
    wire _node_309;
    MUX_UNSIGNED #(.width(1)) u_mux_347 (
        .y(_node_309),
        .sel(_node_308),
        .a(_T_136_52),
        .b(_node_307)
    );
    wire _node_310;
    EQ_UNSIGNED #(.width(7)) u_eq_348 (
        .y(_node_310),
        .a(7'd53),
        .b(_T_454)
    );
    wire _node_311;
    MUX_UNSIGNED #(.width(1)) u_mux_349 (
        .y(_node_311),
        .sel(_node_310),
        .a(_T_136_53),
        .b(_node_309)
    );
    wire _node_312;
    EQ_UNSIGNED #(.width(7)) u_eq_350 (
        .y(_node_312),
        .a(7'd54),
        .b(_T_454)
    );
    wire _node_313;
    MUX_UNSIGNED #(.width(1)) u_mux_351 (
        .y(_node_313),
        .sel(_node_312),
        .a(_T_136_54),
        .b(_node_311)
    );
    wire _node_314;
    EQ_UNSIGNED #(.width(7)) u_eq_352 (
        .y(_node_314),
        .a(7'd55),
        .b(_T_454)
    );
    wire _node_315;
    MUX_UNSIGNED #(.width(1)) u_mux_353 (
        .y(_node_315),
        .sel(_node_314),
        .a(_T_136_55),
        .b(_node_313)
    );
    wire _node_316;
    EQ_UNSIGNED #(.width(7)) u_eq_354 (
        .y(_node_316),
        .a(7'd56),
        .b(_T_454)
    );
    wire _node_317;
    MUX_UNSIGNED #(.width(1)) u_mux_355 (
        .y(_node_317),
        .sel(_node_316),
        .a(_T_136_56),
        .b(_node_315)
    );
    wire _node_318;
    EQ_UNSIGNED #(.width(7)) u_eq_356 (
        .y(_node_318),
        .a(7'd57),
        .b(_T_454)
    );
    wire _node_319;
    MUX_UNSIGNED #(.width(1)) u_mux_357 (
        .y(_node_319),
        .sel(_node_318),
        .a(_T_136_57),
        .b(_node_317)
    );
    wire _node_320;
    EQ_UNSIGNED #(.width(7)) u_eq_358 (
        .y(_node_320),
        .a(7'd58),
        .b(_T_454)
    );
    wire _node_321;
    MUX_UNSIGNED #(.width(1)) u_mux_359 (
        .y(_node_321),
        .sel(_node_320),
        .a(_T_136_58),
        .b(_node_319)
    );
    wire _node_322;
    EQ_UNSIGNED #(.width(7)) u_eq_360 (
        .y(_node_322),
        .a(7'd59),
        .b(_T_454)
    );
    wire _node_323;
    MUX_UNSIGNED #(.width(1)) u_mux_361 (
        .y(_node_323),
        .sel(_node_322),
        .a(_T_136_59),
        .b(_node_321)
    );
    wire _node_324;
    EQ_UNSIGNED #(.width(7)) u_eq_362 (
        .y(_node_324),
        .a(7'd60),
        .b(_T_454)
    );
    wire _node_325;
    MUX_UNSIGNED #(.width(1)) u_mux_363 (
        .y(_node_325),
        .sel(_node_324),
        .a(_T_136_60),
        .b(_node_323)
    );
    wire _node_326;
    EQ_UNSIGNED #(.width(7)) u_eq_364 (
        .y(_node_326),
        .a(7'd61),
        .b(_T_454)
    );
    wire _node_327;
    MUX_UNSIGNED #(.width(1)) u_mux_365 (
        .y(_node_327),
        .sel(_node_326),
        .a(_T_136_61),
        .b(_node_325)
    );
    wire _node_328;
    EQ_UNSIGNED #(.width(7)) u_eq_366 (
        .y(_node_328),
        .a(7'd62),
        .b(_T_454)
    );
    wire _node_329;
    MUX_UNSIGNED #(.width(1)) u_mux_367 (
        .y(_node_329),
        .sel(_node_328),
        .a(_T_136_62),
        .b(_node_327)
    );
    wire _node_330;
    EQ_UNSIGNED #(.width(7)) u_eq_368 (
        .y(_node_330),
        .a(7'd63),
        .b(_T_454)
    );
    wire _node_331;
    MUX_UNSIGNED #(.width(1)) u_mux_369 (
        .y(_node_331),
        .sel(_node_330),
        .a(_T_136_63),
        .b(_node_329)
    );
    wire _node_332;
    EQ_UNSIGNED #(.width(7)) u_eq_370 (
        .y(_node_332),
        .a(7'd64),
        .b(_T_454)
    );
    wire _node_333;
    MUX_UNSIGNED #(.width(1)) u_mux_371 (
        .y(_node_333),
        .sel(_node_332),
        .a(_T_136_64),
        .b(_node_331)
    );
    wire _node_334;
    EQ_UNSIGNED #(.width(7)) u_eq_372 (
        .y(_node_334),
        .a(7'd65),
        .b(_T_454)
    );
    wire _node_335;
    MUX_UNSIGNED #(.width(1)) u_mux_373 (
        .y(_node_335),
        .sel(_node_334),
        .a(_T_136_65),
        .b(_node_333)
    );
    wire _node_336;
    EQ_UNSIGNED #(.width(7)) u_eq_374 (
        .y(_node_336),
        .a(7'd66),
        .b(_T_454)
    );
    wire _node_337;
    MUX_UNSIGNED #(.width(1)) u_mux_375 (
        .y(_node_337),
        .sel(_node_336),
        .a(_T_136_66),
        .b(_node_335)
    );
    wire _node_338;
    EQ_UNSIGNED #(.width(7)) u_eq_376 (
        .y(_node_338),
        .a(7'd67),
        .b(_T_454)
    );
    wire _node_339;
    MUX_UNSIGNED #(.width(1)) u_mux_377 (
        .y(_node_339),
        .sel(_node_338),
        .a(_T_136_67),
        .b(_node_337)
    );
    wire _node_340;
    EQ_UNSIGNED #(.width(7)) u_eq_378 (
        .y(_node_340),
        .a(7'd68),
        .b(_T_454)
    );
    wire _node_341;
    MUX_UNSIGNED #(.width(1)) u_mux_379 (
        .y(_node_341),
        .sel(_node_340),
        .a(_T_136_68),
        .b(_node_339)
    );
    wire _node_342;
    EQ_UNSIGNED #(.width(7)) u_eq_380 (
        .y(_node_342),
        .a(7'd69),
        .b(_T_454)
    );
    wire _node_343;
    MUX_UNSIGNED #(.width(1)) u_mux_381 (
        .y(_node_343),
        .sel(_node_342),
        .a(_T_136_69),
        .b(_node_341)
    );
    wire _node_344;
    EQ_UNSIGNED #(.width(7)) u_eq_382 (
        .y(_node_344),
        .a(7'd70),
        .b(_T_454)
    );
    wire _node_345;
    MUX_UNSIGNED #(.width(1)) u_mux_383 (
        .y(_node_345),
        .sel(_node_344),
        .a(_T_136_70),
        .b(_node_343)
    );
    wire _node_346;
    EQ_UNSIGNED #(.width(7)) u_eq_384 (
        .y(_node_346),
        .a(7'd71),
        .b(_T_454)
    );
    wire _node_347;
    MUX_UNSIGNED #(.width(1)) u_mux_385 (
        .y(_node_347),
        .sel(_node_346),
        .a(_T_136_71),
        .b(_node_345)
    );
    wire _node_348;
    EQ_UNSIGNED #(.width(7)) u_eq_386 (
        .y(_node_348),
        .a(7'd72),
        .b(_T_454)
    );
    wire _node_349;
    MUX_UNSIGNED #(.width(1)) u_mux_387 (
        .y(_node_349),
        .sel(_node_348),
        .a(_T_136_72),
        .b(_node_347)
    );
    wire _node_350;
    EQ_UNSIGNED #(.width(7)) u_eq_388 (
        .y(_node_350),
        .a(7'd73),
        .b(_T_454)
    );
    wire _node_351;
    MUX_UNSIGNED #(.width(1)) u_mux_389 (
        .y(_node_351),
        .sel(_node_350),
        .a(_T_136_73),
        .b(_node_349)
    );
    wire _node_352;
    EQ_UNSIGNED #(.width(7)) u_eq_390 (
        .y(_node_352),
        .a(7'd74),
        .b(_T_454)
    );
    wire _node_353;
    MUX_UNSIGNED #(.width(1)) u_mux_391 (
        .y(_node_353),
        .sel(_node_352),
        .a(_T_136_74),
        .b(_node_351)
    );
    wire _node_354;
    EQ_UNSIGNED #(.width(7)) u_eq_392 (
        .y(_node_354),
        .a(7'd75),
        .b(_T_454)
    );
    wire _node_355;
    MUX_UNSIGNED #(.width(1)) u_mux_393 (
        .y(_node_355),
        .sel(_node_354),
        .a(_T_136_75),
        .b(_node_353)
    );
    wire _node_356;
    EQ_UNSIGNED #(.width(7)) u_eq_394 (
        .y(_node_356),
        .a(7'd76),
        .b(_T_454)
    );
    wire _node_357;
    MUX_UNSIGNED #(.width(1)) u_mux_395 (
        .y(_node_357),
        .sel(_node_356),
        .a(_T_136_76),
        .b(_node_355)
    );
    wire _node_358;
    EQ_UNSIGNED #(.width(7)) u_eq_396 (
        .y(_node_358),
        .a(7'd77),
        .b(_T_454)
    );
    wire _node_359;
    MUX_UNSIGNED #(.width(1)) u_mux_397 (
        .y(_node_359),
        .sel(_node_358),
        .a(_T_136_77),
        .b(_node_357)
    );
    wire _node_360;
    EQ_UNSIGNED #(.width(7)) u_eq_398 (
        .y(_node_360),
        .a(7'd78),
        .b(_T_454)
    );
    wire _node_361;
    MUX_UNSIGNED #(.width(1)) u_mux_399 (
        .y(_node_361),
        .sel(_node_360),
        .a(_T_136_78),
        .b(_node_359)
    );
    wire _node_362;
    EQ_UNSIGNED #(.width(7)) u_eq_400 (
        .y(_node_362),
        .a(7'd79),
        .b(_T_454)
    );
    wire _node_363;
    MUX_UNSIGNED #(.width(1)) u_mux_401 (
        .y(_node_363),
        .sel(_node_362),
        .a(_T_136_79),
        .b(_node_361)
    );
    wire _node_364;
    EQ_UNSIGNED #(.width(7)) u_eq_402 (
        .y(_node_364),
        .a(7'd80),
        .b(_T_454)
    );
    wire _node_365;
    MUX_UNSIGNED #(.width(1)) u_mux_403 (
        .y(_node_365),
        .sel(_node_364),
        .a(_T_136_80),
        .b(_node_363)
    );
    wire _node_366;
    EQ_UNSIGNED #(.width(7)) u_eq_404 (
        .y(_node_366),
        .a(7'd81),
        .b(_T_454)
    );
    wire _node_367;
    MUX_UNSIGNED #(.width(1)) u_mux_405 (
        .y(_node_367),
        .sel(_node_366),
        .a(_T_136_81),
        .b(_node_365)
    );
    wire _node_368;
    EQ_UNSIGNED #(.width(7)) u_eq_406 (
        .y(_node_368),
        .a(7'd82),
        .b(_T_454)
    );
    wire _node_369;
    MUX_UNSIGNED #(.width(1)) u_mux_407 (
        .y(_node_369),
        .sel(_node_368),
        .a(_T_136_82),
        .b(_node_367)
    );
    wire _node_370;
    EQ_UNSIGNED #(.width(7)) u_eq_408 (
        .y(_node_370),
        .a(7'd83),
        .b(_T_454)
    );
    wire _node_371;
    MUX_UNSIGNED #(.width(1)) u_mux_409 (
        .y(_node_371),
        .sel(_node_370),
        .a(_T_136_83),
        .b(_node_369)
    );
    wire _node_372;
    EQ_UNSIGNED #(.width(7)) u_eq_410 (
        .y(_node_372),
        .a(7'd84),
        .b(_T_454)
    );
    wire _node_373;
    MUX_UNSIGNED #(.width(1)) u_mux_411 (
        .y(_node_373),
        .sel(_node_372),
        .a(_T_136_84),
        .b(_node_371)
    );
    wire _node_374;
    EQ_UNSIGNED #(.width(7)) u_eq_412 (
        .y(_node_374),
        .a(7'd85),
        .b(_T_454)
    );
    wire _node_375;
    MUX_UNSIGNED #(.width(1)) u_mux_413 (
        .y(_node_375),
        .sel(_node_374),
        .a(_T_136_85),
        .b(_node_373)
    );
    wire _node_376;
    EQ_UNSIGNED #(.width(7)) u_eq_414 (
        .y(_node_376),
        .a(7'd86),
        .b(_T_454)
    );
    wire _node_377;
    MUX_UNSIGNED #(.width(1)) u_mux_415 (
        .y(_node_377),
        .sel(_node_376),
        .a(_T_136_86),
        .b(_node_375)
    );
    wire _node_378;
    EQ_UNSIGNED #(.width(7)) u_eq_416 (
        .y(_node_378),
        .a(7'd87),
        .b(_T_454)
    );
    wire _node_379;
    MUX_UNSIGNED #(.width(1)) u_mux_417 (
        .y(_node_379),
        .sel(_node_378),
        .a(_T_136_87),
        .b(_node_377)
    );
    wire _node_380;
    EQ_UNSIGNED #(.width(7)) u_eq_418 (
        .y(_node_380),
        .a(7'd88),
        .b(_T_454)
    );
    wire _node_381;
    MUX_UNSIGNED #(.width(1)) u_mux_419 (
        .y(_node_381),
        .sel(_node_380),
        .a(_T_136_88),
        .b(_node_379)
    );
    wire _node_382;
    EQ_UNSIGNED #(.width(7)) u_eq_420 (
        .y(_node_382),
        .a(7'd89),
        .b(_T_454)
    );
    wire _node_383;
    MUX_UNSIGNED #(.width(1)) u_mux_421 (
        .y(_node_383),
        .sel(_node_382),
        .a(_T_136_89),
        .b(_node_381)
    );
    wire _node_384;
    EQ_UNSIGNED #(.width(7)) u_eq_422 (
        .y(_node_384),
        .a(7'd90),
        .b(_T_454)
    );
    wire _node_385;
    MUX_UNSIGNED #(.width(1)) u_mux_423 (
        .y(_node_385),
        .sel(_node_384),
        .a(_T_136_90),
        .b(_node_383)
    );
    wire _node_386;
    EQ_UNSIGNED #(.width(7)) u_eq_424 (
        .y(_node_386),
        .a(7'd91),
        .b(_T_454)
    );
    wire _node_387;
    MUX_UNSIGNED #(.width(1)) u_mux_425 (
        .y(_node_387),
        .sel(_node_386),
        .a(_T_136_91),
        .b(_node_385)
    );
    wire _node_388;
    EQ_UNSIGNED #(.width(7)) u_eq_426 (
        .y(_node_388),
        .a(7'd92),
        .b(_T_454)
    );
    wire _node_389;
    MUX_UNSIGNED #(.width(1)) u_mux_427 (
        .y(_node_389),
        .sel(_node_388),
        .a(_T_136_92),
        .b(_node_387)
    );
    wire _node_390;
    EQ_UNSIGNED #(.width(7)) u_eq_428 (
        .y(_node_390),
        .a(7'd93),
        .b(_T_454)
    );
    wire _node_391;
    MUX_UNSIGNED #(.width(1)) u_mux_429 (
        .y(_node_391),
        .sel(_node_390),
        .a(_T_136_93),
        .b(_node_389)
    );
    wire _node_392;
    EQ_UNSIGNED #(.width(7)) u_eq_430 (
        .y(_node_392),
        .a(7'd94),
        .b(_T_454)
    );
    wire _node_393;
    MUX_UNSIGNED #(.width(1)) u_mux_431 (
        .y(_node_393),
        .sel(_node_392),
        .a(_T_136_94),
        .b(_node_391)
    );
    wire _node_394;
    EQ_UNSIGNED #(.width(7)) u_eq_432 (
        .y(_node_394),
        .a(7'd95),
        .b(_T_454)
    );
    wire _node_395;
    MUX_UNSIGNED #(.width(1)) u_mux_433 (
        .y(_node_395),
        .sel(_node_394),
        .a(_T_136_95),
        .b(_node_393)
    );
    wire _node_396;
    EQ_UNSIGNED #(.width(7)) u_eq_434 (
        .y(_node_396),
        .a(7'd96),
        .b(_T_454)
    );
    wire _node_397;
    MUX_UNSIGNED #(.width(1)) u_mux_435 (
        .y(_node_397),
        .sel(_node_396),
        .a(_T_136_96),
        .b(_node_395)
    );
    wire _node_398;
    EQ_UNSIGNED #(.width(7)) u_eq_436 (
        .y(_node_398),
        .a(7'd97),
        .b(_T_454)
    );
    wire _node_399;
    MUX_UNSIGNED #(.width(1)) u_mux_437 (
        .y(_node_399),
        .sel(_node_398),
        .a(_T_136_97),
        .b(_node_397)
    );
    wire _node_400;
    EQ_UNSIGNED #(.width(7)) u_eq_438 (
        .y(_node_400),
        .a(7'd98),
        .b(_T_454)
    );
    wire _node_401;
    MUX_UNSIGNED #(.width(1)) u_mux_439 (
        .y(_node_401),
        .sel(_node_400),
        .a(_T_136_98),
        .b(_node_399)
    );
    wire _node_402;
    EQ_UNSIGNED #(.width(7)) u_eq_440 (
        .y(_node_402),
        .a(7'd99),
        .b(_T_454)
    );
    wire _node_403;
    MUX_UNSIGNED #(.width(1)) u_mux_441 (
        .y(_node_403),
        .sel(_node_402),
        .a(_T_136_99),
        .b(_node_401)
    );
    wire _node_404;
    EQ_UNSIGNED #(.width(7)) u_eq_442 (
        .y(_node_404),
        .a(7'd100),
        .b(_T_454)
    );
    wire _node_405;
    MUX_UNSIGNED #(.width(1)) u_mux_443 (
        .y(_node_405),
        .sel(_node_404),
        .a(_T_136_100),
        .b(_node_403)
    );
    wire _node_406;
    EQ_UNSIGNED #(.width(7)) u_eq_444 (
        .y(_node_406),
        .a(7'd101),
        .b(_T_454)
    );
    wire _node_407;
    MUX_UNSIGNED #(.width(1)) u_mux_445 (
        .y(_node_407),
        .sel(_node_406),
        .a(_T_136_101),
        .b(_node_405)
    );
    wire _T_455;
    BITWISEAND #(.width(1)) bitwiseand_446 (
        .y(_T_455),
        .a(_device_under_test__io_in_valid),
        .b(_device_under_test__io_in_ready)
    );
    wire _T_457;
    EQ_UNSIGNED #(.width(7)) u_eq_447 (
        .y(_T_457),
        .a(_value__q),
        .b(7'h64)
    );
    wire [7:0] _T_459;
    wire [6:0] _WTEMP_11;
    PAD_UNSIGNED #(.width(1), .n(7)) u_pad_448 (
        .y(_WTEMP_11),
        .in(1'h1)
    );
    ADD_UNSIGNED #(.width(7)) u_add_449 (
        .y(_T_459),
        .a(_value__q),
        .b(_WTEMP_11)
    );
    wire [6:0] _T_460;
    TAIL #(.width(8), .n(1)) tail_450 (
        .y(_T_460),
        .in(_T_459)
    );
    wire _T_463;
    EQ_UNSIGNED #(.width(1)) u_eq_451 (
        .y(_T_463),
        .a(__T_7__q),
        .b(1'h0)
    );
    wire _T_465;
    wire [8:0] _WTEMP_12;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_452 (
        .y(_WTEMP_12),
        .in(7'h64)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_453 (
        .y(_T_465),
        .a(__T_4__q),
        .b(_WTEMP_12)
    );
    wire [9:0] _T_468;
    wire [8:0] _WTEMP_13;
    PAD_UNSIGNED #(.width(1), .n(9)) u_pad_454 (
        .y(_WTEMP_13),
        .in(1'h1)
    );
    ADD_UNSIGNED #(.width(9)) u_add_455 (
        .y(_T_468),
        .a(__T_4__q),
        .b(_WTEMP_13)
    );
    wire [8:0] _T_469;
    TAIL #(.width(10), .n(1)) tail_456 (
        .y(_T_469),
        .in(_T_468)
    );
    wire _node_408;
    MUX_UNSIGNED #(.width(1)) u_mux_457 (
        .y(_node_408),
        .sel(_T_465),
        .a(1'h1),
        .b(__T_7__q)
    );
    wire [8:0] _node_409;
    MUX_UNSIGNED #(.width(9)) u_mux_458 (
        .y(_node_409),
        .sel(_T_463),
        .a(_T_469),
        .b(__T_4__q)
    );
    wire _node_410;
    MUX_UNSIGNED #(.width(1)) u_mux_459 (
        .y(_node_410),
        .sel(_T_463),
        .a(_node_408),
        .b(__T_7__q)
    );
    wire [6:0] _node_411;
    wire [6:0] _WTEMP_14;
    PAD_UNSIGNED #(.width(1), .n(7)) u_pad_460 (
        .y(_WTEMP_14),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(7)) u_mux_461 (
        .y(_node_411),
        .sel(_T_457),
        .a(_WTEMP_14),
        .b(_T_460)
    );
    wire _T_574_0;
    wire _T_574_1;
    wire _T_574_2;
    wire _T_574_3;
    wire _T_574_4;
    wire _T_574_5;
    wire _T_574_6;
    wire _T_574_7;
    wire _T_574_8;
    wire _T_574_9;
    wire _T_574_10;
    wire _T_574_11;
    wire _T_574_12;
    wire _T_574_13;
    wire _T_574_14;
    wire _T_574_15;
    wire _T_574_16;
    wire _T_574_17;
    wire _T_574_18;
    wire _T_574_19;
    wire _T_574_20;
    wire _T_574_21;
    wire _T_574_22;
    wire _T_574_23;
    wire _T_574_24;
    wire _T_574_25;
    wire _T_574_26;
    wire _T_574_27;
    wire _T_574_28;
    wire _T_574_29;
    wire _T_574_30;
    wire _T_574_31;
    wire _T_574_32;
    wire _T_574_33;
    wire _T_574_34;
    wire _T_574_35;
    wire _T_574_36;
    wire _T_574_37;
    wire _T_574_38;
    wire _T_574_39;
    wire _T_574_40;
    wire _T_574_41;
    wire _T_574_42;
    wire _T_574_43;
    wire _T_574_44;
    wire _T_574_45;
    wire _T_574_46;
    wire _T_574_47;
    wire _T_574_48;
    wire _T_574_49;
    wire _T_574_50;
    wire _T_574_51;
    wire _T_574_52;
    wire _T_574_53;
    wire _T_574_54;
    wire _T_574_55;
    wire _T_574_56;
    wire _T_574_57;
    wire _T_574_58;
    wire _T_574_59;
    wire _T_574_60;
    wire _T_574_61;
    wire _T_574_62;
    wire _T_574_63;
    wire _T_574_64;
    wire _T_574_65;
    wire _T_574_66;
    wire _T_574_67;
    wire _T_574_68;
    wire _T_574_69;
    wire _T_574_70;
    wire _T_574_71;
    wire _T_574_72;
    wire _T_574_73;
    wire _T_574_74;
    wire _T_574_75;
    wire _T_574_76;
    wire _T_574_77;
    wire _T_574_78;
    wire _T_574_79;
    wire _T_574_80;
    wire _T_574_81;
    wire _T_574_82;
    wire _T_574_83;
    wire _T_574_84;
    wire _T_574_85;
    wire _T_574_86;
    wire _T_574_87;
    wire _T_574_88;
    wire _T_574_89;
    wire _T_574_90;
    wire _T_574_91;
    wire _T_574_92;
    wire _T_574_93;
    wire _T_574_94;
    wire _T_574_95;
    wire _T_574_96;
    wire _T_574_97;
    wire _T_574_98;
    wire _T_574_99;
    wire _T_574_100;
    wire _T_574_101;
    wire [4:0] _value_1__q;
    wire [4:0] _value_1__d;
    DFF_POSCLK #(.width(5)) value_1 (
        .q(_value_1__q),
        .d(_value_1__d),
        .clk(clock)
    );
    wire [4:0] _WTEMP_15;
    MUX_UNSIGNED #(.width(5)) u_mux_462 (
        .y(_value_1__d),
        .sel(reset),
        .a(5'h0),
        .b(_WTEMP_15)
    );
    wire [3:0] _T_711_0;
    wire [3:0] _T_711_1;
    wire [3:0] _T_711_2;
    wire [3:0] _T_711_3;
    wire [3:0] _T_711_4;
    wire [3:0] _T_711_5;
    wire [3:0] _T_711_6;
    wire [3:0] _T_711_7;
    wire [3:0] _T_711_8;
    wire [3:0] _T_711_9;
    wire [3:0] _T_711_10;
    wire [3:0] _T_711_11;
    wire [3:0] _T_711_12;
    wire [3:0] _T_711_13;
    wire [3:0] _T_711_14;
    wire [3:0] _T_711_15;
    wire [3:0] _T_711_16;
    wire [3:0] _T_711_17;
    wire [3:0] _T_711_18;
    wire [3:0] _T_711_19;
    wire [3:0] _T_711_20;
    wire [3:0] _T_711_21;
    wire [3:0] _T_711_22;
    wire [3:0] _T_711_23;
    wire [3:0] _T_711_24;
    wire [3:0] _T_711_25;
    wire [3:0] _T_711_26;
    wire [3:0] _T_711_27;
    wire _node_412;
    EQ_UNSIGNED #(.width(7)) u_eq_463 (
        .y(_node_412),
        .a(7'd0),
        .b(__T_10__q)
    );
    wire _node_413;
    assign _node_413 = _T_574_0;
    wire _node_414;
    EQ_UNSIGNED #(.width(7)) u_eq_464 (
        .y(_node_414),
        .a(7'd1),
        .b(__T_10__q)
    );
    wire _node_415;
    MUX_UNSIGNED #(.width(1)) u_mux_465 (
        .y(_node_415),
        .sel(_node_414),
        .a(_T_574_1),
        .b(_node_413)
    );
    wire _node_416;
    EQ_UNSIGNED #(.width(7)) u_eq_466 (
        .y(_node_416),
        .a(7'd2),
        .b(__T_10__q)
    );
    wire _node_417;
    MUX_UNSIGNED #(.width(1)) u_mux_467 (
        .y(_node_417),
        .sel(_node_416),
        .a(_T_574_2),
        .b(_node_415)
    );
    wire _node_418;
    EQ_UNSIGNED #(.width(7)) u_eq_468 (
        .y(_node_418),
        .a(7'd3),
        .b(__T_10__q)
    );
    wire _node_419;
    MUX_UNSIGNED #(.width(1)) u_mux_469 (
        .y(_node_419),
        .sel(_node_418),
        .a(_T_574_3),
        .b(_node_417)
    );
    wire _node_420;
    EQ_UNSIGNED #(.width(7)) u_eq_470 (
        .y(_node_420),
        .a(7'd4),
        .b(__T_10__q)
    );
    wire _node_421;
    MUX_UNSIGNED #(.width(1)) u_mux_471 (
        .y(_node_421),
        .sel(_node_420),
        .a(_T_574_4),
        .b(_node_419)
    );
    wire _node_422;
    EQ_UNSIGNED #(.width(7)) u_eq_472 (
        .y(_node_422),
        .a(7'd5),
        .b(__T_10__q)
    );
    wire _node_423;
    MUX_UNSIGNED #(.width(1)) u_mux_473 (
        .y(_node_423),
        .sel(_node_422),
        .a(_T_574_5),
        .b(_node_421)
    );
    wire _node_424;
    EQ_UNSIGNED #(.width(7)) u_eq_474 (
        .y(_node_424),
        .a(7'd6),
        .b(__T_10__q)
    );
    wire _node_425;
    MUX_UNSIGNED #(.width(1)) u_mux_475 (
        .y(_node_425),
        .sel(_node_424),
        .a(_T_574_6),
        .b(_node_423)
    );
    wire _node_426;
    EQ_UNSIGNED #(.width(7)) u_eq_476 (
        .y(_node_426),
        .a(7'd7),
        .b(__T_10__q)
    );
    wire _node_427;
    MUX_UNSIGNED #(.width(1)) u_mux_477 (
        .y(_node_427),
        .sel(_node_426),
        .a(_T_574_7),
        .b(_node_425)
    );
    wire _node_428;
    EQ_UNSIGNED #(.width(7)) u_eq_478 (
        .y(_node_428),
        .a(7'd8),
        .b(__T_10__q)
    );
    wire _node_429;
    MUX_UNSIGNED #(.width(1)) u_mux_479 (
        .y(_node_429),
        .sel(_node_428),
        .a(_T_574_8),
        .b(_node_427)
    );
    wire _node_430;
    EQ_UNSIGNED #(.width(7)) u_eq_480 (
        .y(_node_430),
        .a(7'd9),
        .b(__T_10__q)
    );
    wire _node_431;
    MUX_UNSIGNED #(.width(1)) u_mux_481 (
        .y(_node_431),
        .sel(_node_430),
        .a(_T_574_9),
        .b(_node_429)
    );
    wire _node_432;
    EQ_UNSIGNED #(.width(7)) u_eq_482 (
        .y(_node_432),
        .a(7'd10),
        .b(__T_10__q)
    );
    wire _node_433;
    MUX_UNSIGNED #(.width(1)) u_mux_483 (
        .y(_node_433),
        .sel(_node_432),
        .a(_T_574_10),
        .b(_node_431)
    );
    wire _node_434;
    EQ_UNSIGNED #(.width(7)) u_eq_484 (
        .y(_node_434),
        .a(7'd11),
        .b(__T_10__q)
    );
    wire _node_435;
    MUX_UNSIGNED #(.width(1)) u_mux_485 (
        .y(_node_435),
        .sel(_node_434),
        .a(_T_574_11),
        .b(_node_433)
    );
    wire _node_436;
    EQ_UNSIGNED #(.width(7)) u_eq_486 (
        .y(_node_436),
        .a(7'd12),
        .b(__T_10__q)
    );
    wire _node_437;
    MUX_UNSIGNED #(.width(1)) u_mux_487 (
        .y(_node_437),
        .sel(_node_436),
        .a(_T_574_12),
        .b(_node_435)
    );
    wire _node_438;
    EQ_UNSIGNED #(.width(7)) u_eq_488 (
        .y(_node_438),
        .a(7'd13),
        .b(__T_10__q)
    );
    wire _node_439;
    MUX_UNSIGNED #(.width(1)) u_mux_489 (
        .y(_node_439),
        .sel(_node_438),
        .a(_T_574_13),
        .b(_node_437)
    );
    wire _node_440;
    EQ_UNSIGNED #(.width(7)) u_eq_490 (
        .y(_node_440),
        .a(7'd14),
        .b(__T_10__q)
    );
    wire _node_441;
    MUX_UNSIGNED #(.width(1)) u_mux_491 (
        .y(_node_441),
        .sel(_node_440),
        .a(_T_574_14),
        .b(_node_439)
    );
    wire _node_442;
    EQ_UNSIGNED #(.width(7)) u_eq_492 (
        .y(_node_442),
        .a(7'd15),
        .b(__T_10__q)
    );
    wire _node_443;
    MUX_UNSIGNED #(.width(1)) u_mux_493 (
        .y(_node_443),
        .sel(_node_442),
        .a(_T_574_15),
        .b(_node_441)
    );
    wire _node_444;
    EQ_UNSIGNED #(.width(7)) u_eq_494 (
        .y(_node_444),
        .a(7'd16),
        .b(__T_10__q)
    );
    wire _node_445;
    MUX_UNSIGNED #(.width(1)) u_mux_495 (
        .y(_node_445),
        .sel(_node_444),
        .a(_T_574_16),
        .b(_node_443)
    );
    wire _node_446;
    EQ_UNSIGNED #(.width(7)) u_eq_496 (
        .y(_node_446),
        .a(7'd17),
        .b(__T_10__q)
    );
    wire _node_447;
    MUX_UNSIGNED #(.width(1)) u_mux_497 (
        .y(_node_447),
        .sel(_node_446),
        .a(_T_574_17),
        .b(_node_445)
    );
    wire _node_448;
    EQ_UNSIGNED #(.width(7)) u_eq_498 (
        .y(_node_448),
        .a(7'd18),
        .b(__T_10__q)
    );
    wire _node_449;
    MUX_UNSIGNED #(.width(1)) u_mux_499 (
        .y(_node_449),
        .sel(_node_448),
        .a(_T_574_18),
        .b(_node_447)
    );
    wire _node_450;
    EQ_UNSIGNED #(.width(7)) u_eq_500 (
        .y(_node_450),
        .a(7'd19),
        .b(__T_10__q)
    );
    wire _node_451;
    MUX_UNSIGNED #(.width(1)) u_mux_501 (
        .y(_node_451),
        .sel(_node_450),
        .a(_T_574_19),
        .b(_node_449)
    );
    wire _node_452;
    EQ_UNSIGNED #(.width(7)) u_eq_502 (
        .y(_node_452),
        .a(7'd20),
        .b(__T_10__q)
    );
    wire _node_453;
    MUX_UNSIGNED #(.width(1)) u_mux_503 (
        .y(_node_453),
        .sel(_node_452),
        .a(_T_574_20),
        .b(_node_451)
    );
    wire _node_454;
    EQ_UNSIGNED #(.width(7)) u_eq_504 (
        .y(_node_454),
        .a(7'd21),
        .b(__T_10__q)
    );
    wire _node_455;
    MUX_UNSIGNED #(.width(1)) u_mux_505 (
        .y(_node_455),
        .sel(_node_454),
        .a(_T_574_21),
        .b(_node_453)
    );
    wire _node_456;
    EQ_UNSIGNED #(.width(7)) u_eq_506 (
        .y(_node_456),
        .a(7'd22),
        .b(__T_10__q)
    );
    wire _node_457;
    MUX_UNSIGNED #(.width(1)) u_mux_507 (
        .y(_node_457),
        .sel(_node_456),
        .a(_T_574_22),
        .b(_node_455)
    );
    wire _node_458;
    EQ_UNSIGNED #(.width(7)) u_eq_508 (
        .y(_node_458),
        .a(7'd23),
        .b(__T_10__q)
    );
    wire _node_459;
    MUX_UNSIGNED #(.width(1)) u_mux_509 (
        .y(_node_459),
        .sel(_node_458),
        .a(_T_574_23),
        .b(_node_457)
    );
    wire _node_460;
    EQ_UNSIGNED #(.width(7)) u_eq_510 (
        .y(_node_460),
        .a(7'd24),
        .b(__T_10__q)
    );
    wire _node_461;
    MUX_UNSIGNED #(.width(1)) u_mux_511 (
        .y(_node_461),
        .sel(_node_460),
        .a(_T_574_24),
        .b(_node_459)
    );
    wire _node_462;
    EQ_UNSIGNED #(.width(7)) u_eq_512 (
        .y(_node_462),
        .a(7'd25),
        .b(__T_10__q)
    );
    wire _node_463;
    MUX_UNSIGNED #(.width(1)) u_mux_513 (
        .y(_node_463),
        .sel(_node_462),
        .a(_T_574_25),
        .b(_node_461)
    );
    wire _node_464;
    EQ_UNSIGNED #(.width(7)) u_eq_514 (
        .y(_node_464),
        .a(7'd26),
        .b(__T_10__q)
    );
    wire _node_465;
    MUX_UNSIGNED #(.width(1)) u_mux_515 (
        .y(_node_465),
        .sel(_node_464),
        .a(_T_574_26),
        .b(_node_463)
    );
    wire _node_466;
    EQ_UNSIGNED #(.width(7)) u_eq_516 (
        .y(_node_466),
        .a(7'd27),
        .b(__T_10__q)
    );
    wire _node_467;
    MUX_UNSIGNED #(.width(1)) u_mux_517 (
        .y(_node_467),
        .sel(_node_466),
        .a(_T_574_27),
        .b(_node_465)
    );
    wire _node_468;
    EQ_UNSIGNED #(.width(7)) u_eq_518 (
        .y(_node_468),
        .a(7'd28),
        .b(__T_10__q)
    );
    wire _node_469;
    MUX_UNSIGNED #(.width(1)) u_mux_519 (
        .y(_node_469),
        .sel(_node_468),
        .a(_T_574_28),
        .b(_node_467)
    );
    wire _node_470;
    EQ_UNSIGNED #(.width(7)) u_eq_520 (
        .y(_node_470),
        .a(7'd29),
        .b(__T_10__q)
    );
    wire _node_471;
    MUX_UNSIGNED #(.width(1)) u_mux_521 (
        .y(_node_471),
        .sel(_node_470),
        .a(_T_574_29),
        .b(_node_469)
    );
    wire _node_472;
    EQ_UNSIGNED #(.width(7)) u_eq_522 (
        .y(_node_472),
        .a(7'd30),
        .b(__T_10__q)
    );
    wire _node_473;
    MUX_UNSIGNED #(.width(1)) u_mux_523 (
        .y(_node_473),
        .sel(_node_472),
        .a(_T_574_30),
        .b(_node_471)
    );
    wire _node_474;
    EQ_UNSIGNED #(.width(7)) u_eq_524 (
        .y(_node_474),
        .a(7'd31),
        .b(__T_10__q)
    );
    wire _node_475;
    MUX_UNSIGNED #(.width(1)) u_mux_525 (
        .y(_node_475),
        .sel(_node_474),
        .a(_T_574_31),
        .b(_node_473)
    );
    wire _node_476;
    EQ_UNSIGNED #(.width(7)) u_eq_526 (
        .y(_node_476),
        .a(7'd32),
        .b(__T_10__q)
    );
    wire _node_477;
    MUX_UNSIGNED #(.width(1)) u_mux_527 (
        .y(_node_477),
        .sel(_node_476),
        .a(_T_574_32),
        .b(_node_475)
    );
    wire _node_478;
    EQ_UNSIGNED #(.width(7)) u_eq_528 (
        .y(_node_478),
        .a(7'd33),
        .b(__T_10__q)
    );
    wire _node_479;
    MUX_UNSIGNED #(.width(1)) u_mux_529 (
        .y(_node_479),
        .sel(_node_478),
        .a(_T_574_33),
        .b(_node_477)
    );
    wire _node_480;
    EQ_UNSIGNED #(.width(7)) u_eq_530 (
        .y(_node_480),
        .a(7'd34),
        .b(__T_10__q)
    );
    wire _node_481;
    MUX_UNSIGNED #(.width(1)) u_mux_531 (
        .y(_node_481),
        .sel(_node_480),
        .a(_T_574_34),
        .b(_node_479)
    );
    wire _node_482;
    EQ_UNSIGNED #(.width(7)) u_eq_532 (
        .y(_node_482),
        .a(7'd35),
        .b(__T_10__q)
    );
    wire _node_483;
    MUX_UNSIGNED #(.width(1)) u_mux_533 (
        .y(_node_483),
        .sel(_node_482),
        .a(_T_574_35),
        .b(_node_481)
    );
    wire _node_484;
    EQ_UNSIGNED #(.width(7)) u_eq_534 (
        .y(_node_484),
        .a(7'd36),
        .b(__T_10__q)
    );
    wire _node_485;
    MUX_UNSIGNED #(.width(1)) u_mux_535 (
        .y(_node_485),
        .sel(_node_484),
        .a(_T_574_36),
        .b(_node_483)
    );
    wire _node_486;
    EQ_UNSIGNED #(.width(7)) u_eq_536 (
        .y(_node_486),
        .a(7'd37),
        .b(__T_10__q)
    );
    wire _node_487;
    MUX_UNSIGNED #(.width(1)) u_mux_537 (
        .y(_node_487),
        .sel(_node_486),
        .a(_T_574_37),
        .b(_node_485)
    );
    wire _node_488;
    EQ_UNSIGNED #(.width(7)) u_eq_538 (
        .y(_node_488),
        .a(7'd38),
        .b(__T_10__q)
    );
    wire _node_489;
    MUX_UNSIGNED #(.width(1)) u_mux_539 (
        .y(_node_489),
        .sel(_node_488),
        .a(_T_574_38),
        .b(_node_487)
    );
    wire _node_490;
    EQ_UNSIGNED #(.width(7)) u_eq_540 (
        .y(_node_490),
        .a(7'd39),
        .b(__T_10__q)
    );
    wire _node_491;
    MUX_UNSIGNED #(.width(1)) u_mux_541 (
        .y(_node_491),
        .sel(_node_490),
        .a(_T_574_39),
        .b(_node_489)
    );
    wire _node_492;
    EQ_UNSIGNED #(.width(7)) u_eq_542 (
        .y(_node_492),
        .a(7'd40),
        .b(__T_10__q)
    );
    wire _node_493;
    MUX_UNSIGNED #(.width(1)) u_mux_543 (
        .y(_node_493),
        .sel(_node_492),
        .a(_T_574_40),
        .b(_node_491)
    );
    wire _node_494;
    EQ_UNSIGNED #(.width(7)) u_eq_544 (
        .y(_node_494),
        .a(7'd41),
        .b(__T_10__q)
    );
    wire _node_495;
    MUX_UNSIGNED #(.width(1)) u_mux_545 (
        .y(_node_495),
        .sel(_node_494),
        .a(_T_574_41),
        .b(_node_493)
    );
    wire _node_496;
    EQ_UNSIGNED #(.width(7)) u_eq_546 (
        .y(_node_496),
        .a(7'd42),
        .b(__T_10__q)
    );
    wire _node_497;
    MUX_UNSIGNED #(.width(1)) u_mux_547 (
        .y(_node_497),
        .sel(_node_496),
        .a(_T_574_42),
        .b(_node_495)
    );
    wire _node_498;
    EQ_UNSIGNED #(.width(7)) u_eq_548 (
        .y(_node_498),
        .a(7'd43),
        .b(__T_10__q)
    );
    wire _node_499;
    MUX_UNSIGNED #(.width(1)) u_mux_549 (
        .y(_node_499),
        .sel(_node_498),
        .a(_T_574_43),
        .b(_node_497)
    );
    wire _node_500;
    EQ_UNSIGNED #(.width(7)) u_eq_550 (
        .y(_node_500),
        .a(7'd44),
        .b(__T_10__q)
    );
    wire _node_501;
    MUX_UNSIGNED #(.width(1)) u_mux_551 (
        .y(_node_501),
        .sel(_node_500),
        .a(_T_574_44),
        .b(_node_499)
    );
    wire _node_502;
    EQ_UNSIGNED #(.width(7)) u_eq_552 (
        .y(_node_502),
        .a(7'd45),
        .b(__T_10__q)
    );
    wire _node_503;
    MUX_UNSIGNED #(.width(1)) u_mux_553 (
        .y(_node_503),
        .sel(_node_502),
        .a(_T_574_45),
        .b(_node_501)
    );
    wire _node_504;
    EQ_UNSIGNED #(.width(7)) u_eq_554 (
        .y(_node_504),
        .a(7'd46),
        .b(__T_10__q)
    );
    wire _node_505;
    MUX_UNSIGNED #(.width(1)) u_mux_555 (
        .y(_node_505),
        .sel(_node_504),
        .a(_T_574_46),
        .b(_node_503)
    );
    wire _node_506;
    EQ_UNSIGNED #(.width(7)) u_eq_556 (
        .y(_node_506),
        .a(7'd47),
        .b(__T_10__q)
    );
    wire _node_507;
    MUX_UNSIGNED #(.width(1)) u_mux_557 (
        .y(_node_507),
        .sel(_node_506),
        .a(_T_574_47),
        .b(_node_505)
    );
    wire _node_508;
    EQ_UNSIGNED #(.width(7)) u_eq_558 (
        .y(_node_508),
        .a(7'd48),
        .b(__T_10__q)
    );
    wire _node_509;
    MUX_UNSIGNED #(.width(1)) u_mux_559 (
        .y(_node_509),
        .sel(_node_508),
        .a(_T_574_48),
        .b(_node_507)
    );
    wire _node_510;
    EQ_UNSIGNED #(.width(7)) u_eq_560 (
        .y(_node_510),
        .a(7'd49),
        .b(__T_10__q)
    );
    wire _node_511;
    MUX_UNSIGNED #(.width(1)) u_mux_561 (
        .y(_node_511),
        .sel(_node_510),
        .a(_T_574_49),
        .b(_node_509)
    );
    wire _node_512;
    EQ_UNSIGNED #(.width(7)) u_eq_562 (
        .y(_node_512),
        .a(7'd50),
        .b(__T_10__q)
    );
    wire _node_513;
    MUX_UNSIGNED #(.width(1)) u_mux_563 (
        .y(_node_513),
        .sel(_node_512),
        .a(_T_574_50),
        .b(_node_511)
    );
    wire _node_514;
    EQ_UNSIGNED #(.width(7)) u_eq_564 (
        .y(_node_514),
        .a(7'd51),
        .b(__T_10__q)
    );
    wire _node_515;
    MUX_UNSIGNED #(.width(1)) u_mux_565 (
        .y(_node_515),
        .sel(_node_514),
        .a(_T_574_51),
        .b(_node_513)
    );
    wire _node_516;
    EQ_UNSIGNED #(.width(7)) u_eq_566 (
        .y(_node_516),
        .a(7'd52),
        .b(__T_10__q)
    );
    wire _node_517;
    MUX_UNSIGNED #(.width(1)) u_mux_567 (
        .y(_node_517),
        .sel(_node_516),
        .a(_T_574_52),
        .b(_node_515)
    );
    wire _node_518;
    EQ_UNSIGNED #(.width(7)) u_eq_568 (
        .y(_node_518),
        .a(7'd53),
        .b(__T_10__q)
    );
    wire _node_519;
    MUX_UNSIGNED #(.width(1)) u_mux_569 (
        .y(_node_519),
        .sel(_node_518),
        .a(_T_574_53),
        .b(_node_517)
    );
    wire _node_520;
    EQ_UNSIGNED #(.width(7)) u_eq_570 (
        .y(_node_520),
        .a(7'd54),
        .b(__T_10__q)
    );
    wire _node_521;
    MUX_UNSIGNED #(.width(1)) u_mux_571 (
        .y(_node_521),
        .sel(_node_520),
        .a(_T_574_54),
        .b(_node_519)
    );
    wire _node_522;
    EQ_UNSIGNED #(.width(7)) u_eq_572 (
        .y(_node_522),
        .a(7'd55),
        .b(__T_10__q)
    );
    wire _node_523;
    MUX_UNSIGNED #(.width(1)) u_mux_573 (
        .y(_node_523),
        .sel(_node_522),
        .a(_T_574_55),
        .b(_node_521)
    );
    wire _node_524;
    EQ_UNSIGNED #(.width(7)) u_eq_574 (
        .y(_node_524),
        .a(7'd56),
        .b(__T_10__q)
    );
    wire _node_525;
    MUX_UNSIGNED #(.width(1)) u_mux_575 (
        .y(_node_525),
        .sel(_node_524),
        .a(_T_574_56),
        .b(_node_523)
    );
    wire _node_526;
    EQ_UNSIGNED #(.width(7)) u_eq_576 (
        .y(_node_526),
        .a(7'd57),
        .b(__T_10__q)
    );
    wire _node_527;
    MUX_UNSIGNED #(.width(1)) u_mux_577 (
        .y(_node_527),
        .sel(_node_526),
        .a(_T_574_57),
        .b(_node_525)
    );
    wire _node_528;
    EQ_UNSIGNED #(.width(7)) u_eq_578 (
        .y(_node_528),
        .a(7'd58),
        .b(__T_10__q)
    );
    wire _node_529;
    MUX_UNSIGNED #(.width(1)) u_mux_579 (
        .y(_node_529),
        .sel(_node_528),
        .a(_T_574_58),
        .b(_node_527)
    );
    wire _node_530;
    EQ_UNSIGNED #(.width(7)) u_eq_580 (
        .y(_node_530),
        .a(7'd59),
        .b(__T_10__q)
    );
    wire _node_531;
    MUX_UNSIGNED #(.width(1)) u_mux_581 (
        .y(_node_531),
        .sel(_node_530),
        .a(_T_574_59),
        .b(_node_529)
    );
    wire _node_532;
    EQ_UNSIGNED #(.width(7)) u_eq_582 (
        .y(_node_532),
        .a(7'd60),
        .b(__T_10__q)
    );
    wire _node_533;
    MUX_UNSIGNED #(.width(1)) u_mux_583 (
        .y(_node_533),
        .sel(_node_532),
        .a(_T_574_60),
        .b(_node_531)
    );
    wire _node_534;
    EQ_UNSIGNED #(.width(7)) u_eq_584 (
        .y(_node_534),
        .a(7'd61),
        .b(__T_10__q)
    );
    wire _node_535;
    MUX_UNSIGNED #(.width(1)) u_mux_585 (
        .y(_node_535),
        .sel(_node_534),
        .a(_T_574_61),
        .b(_node_533)
    );
    wire _node_536;
    EQ_UNSIGNED #(.width(7)) u_eq_586 (
        .y(_node_536),
        .a(7'd62),
        .b(__T_10__q)
    );
    wire _node_537;
    MUX_UNSIGNED #(.width(1)) u_mux_587 (
        .y(_node_537),
        .sel(_node_536),
        .a(_T_574_62),
        .b(_node_535)
    );
    wire _node_538;
    EQ_UNSIGNED #(.width(7)) u_eq_588 (
        .y(_node_538),
        .a(7'd63),
        .b(__T_10__q)
    );
    wire _node_539;
    MUX_UNSIGNED #(.width(1)) u_mux_589 (
        .y(_node_539),
        .sel(_node_538),
        .a(_T_574_63),
        .b(_node_537)
    );
    wire _node_540;
    EQ_UNSIGNED #(.width(7)) u_eq_590 (
        .y(_node_540),
        .a(7'd64),
        .b(__T_10__q)
    );
    wire _node_541;
    MUX_UNSIGNED #(.width(1)) u_mux_591 (
        .y(_node_541),
        .sel(_node_540),
        .a(_T_574_64),
        .b(_node_539)
    );
    wire _node_542;
    EQ_UNSIGNED #(.width(7)) u_eq_592 (
        .y(_node_542),
        .a(7'd65),
        .b(__T_10__q)
    );
    wire _node_543;
    MUX_UNSIGNED #(.width(1)) u_mux_593 (
        .y(_node_543),
        .sel(_node_542),
        .a(_T_574_65),
        .b(_node_541)
    );
    wire _node_544;
    EQ_UNSIGNED #(.width(7)) u_eq_594 (
        .y(_node_544),
        .a(7'd66),
        .b(__T_10__q)
    );
    wire _node_545;
    MUX_UNSIGNED #(.width(1)) u_mux_595 (
        .y(_node_545),
        .sel(_node_544),
        .a(_T_574_66),
        .b(_node_543)
    );
    wire _node_546;
    EQ_UNSIGNED #(.width(7)) u_eq_596 (
        .y(_node_546),
        .a(7'd67),
        .b(__T_10__q)
    );
    wire _node_547;
    MUX_UNSIGNED #(.width(1)) u_mux_597 (
        .y(_node_547),
        .sel(_node_546),
        .a(_T_574_67),
        .b(_node_545)
    );
    wire _node_548;
    EQ_UNSIGNED #(.width(7)) u_eq_598 (
        .y(_node_548),
        .a(7'd68),
        .b(__T_10__q)
    );
    wire _node_549;
    MUX_UNSIGNED #(.width(1)) u_mux_599 (
        .y(_node_549),
        .sel(_node_548),
        .a(_T_574_68),
        .b(_node_547)
    );
    wire _node_550;
    EQ_UNSIGNED #(.width(7)) u_eq_600 (
        .y(_node_550),
        .a(7'd69),
        .b(__T_10__q)
    );
    wire _node_551;
    MUX_UNSIGNED #(.width(1)) u_mux_601 (
        .y(_node_551),
        .sel(_node_550),
        .a(_T_574_69),
        .b(_node_549)
    );
    wire _node_552;
    EQ_UNSIGNED #(.width(7)) u_eq_602 (
        .y(_node_552),
        .a(7'd70),
        .b(__T_10__q)
    );
    wire _node_553;
    MUX_UNSIGNED #(.width(1)) u_mux_603 (
        .y(_node_553),
        .sel(_node_552),
        .a(_T_574_70),
        .b(_node_551)
    );
    wire _node_554;
    EQ_UNSIGNED #(.width(7)) u_eq_604 (
        .y(_node_554),
        .a(7'd71),
        .b(__T_10__q)
    );
    wire _node_555;
    MUX_UNSIGNED #(.width(1)) u_mux_605 (
        .y(_node_555),
        .sel(_node_554),
        .a(_T_574_71),
        .b(_node_553)
    );
    wire _node_556;
    EQ_UNSIGNED #(.width(7)) u_eq_606 (
        .y(_node_556),
        .a(7'd72),
        .b(__T_10__q)
    );
    wire _node_557;
    MUX_UNSIGNED #(.width(1)) u_mux_607 (
        .y(_node_557),
        .sel(_node_556),
        .a(_T_574_72),
        .b(_node_555)
    );
    wire _node_558;
    EQ_UNSIGNED #(.width(7)) u_eq_608 (
        .y(_node_558),
        .a(7'd73),
        .b(__T_10__q)
    );
    wire _node_559;
    MUX_UNSIGNED #(.width(1)) u_mux_609 (
        .y(_node_559),
        .sel(_node_558),
        .a(_T_574_73),
        .b(_node_557)
    );
    wire _node_560;
    EQ_UNSIGNED #(.width(7)) u_eq_610 (
        .y(_node_560),
        .a(7'd74),
        .b(__T_10__q)
    );
    wire _node_561;
    MUX_UNSIGNED #(.width(1)) u_mux_611 (
        .y(_node_561),
        .sel(_node_560),
        .a(_T_574_74),
        .b(_node_559)
    );
    wire _node_562;
    EQ_UNSIGNED #(.width(7)) u_eq_612 (
        .y(_node_562),
        .a(7'd75),
        .b(__T_10__q)
    );
    wire _node_563;
    MUX_UNSIGNED #(.width(1)) u_mux_613 (
        .y(_node_563),
        .sel(_node_562),
        .a(_T_574_75),
        .b(_node_561)
    );
    wire _node_564;
    EQ_UNSIGNED #(.width(7)) u_eq_614 (
        .y(_node_564),
        .a(7'd76),
        .b(__T_10__q)
    );
    wire _node_565;
    MUX_UNSIGNED #(.width(1)) u_mux_615 (
        .y(_node_565),
        .sel(_node_564),
        .a(_T_574_76),
        .b(_node_563)
    );
    wire _node_566;
    EQ_UNSIGNED #(.width(7)) u_eq_616 (
        .y(_node_566),
        .a(7'd77),
        .b(__T_10__q)
    );
    wire _node_567;
    MUX_UNSIGNED #(.width(1)) u_mux_617 (
        .y(_node_567),
        .sel(_node_566),
        .a(_T_574_77),
        .b(_node_565)
    );
    wire _node_568;
    EQ_UNSIGNED #(.width(7)) u_eq_618 (
        .y(_node_568),
        .a(7'd78),
        .b(__T_10__q)
    );
    wire _node_569;
    MUX_UNSIGNED #(.width(1)) u_mux_619 (
        .y(_node_569),
        .sel(_node_568),
        .a(_T_574_78),
        .b(_node_567)
    );
    wire _node_570;
    EQ_UNSIGNED #(.width(7)) u_eq_620 (
        .y(_node_570),
        .a(7'd79),
        .b(__T_10__q)
    );
    wire _node_571;
    MUX_UNSIGNED #(.width(1)) u_mux_621 (
        .y(_node_571),
        .sel(_node_570),
        .a(_T_574_79),
        .b(_node_569)
    );
    wire _node_572;
    EQ_UNSIGNED #(.width(7)) u_eq_622 (
        .y(_node_572),
        .a(7'd80),
        .b(__T_10__q)
    );
    wire _node_573;
    MUX_UNSIGNED #(.width(1)) u_mux_623 (
        .y(_node_573),
        .sel(_node_572),
        .a(_T_574_80),
        .b(_node_571)
    );
    wire _node_574;
    EQ_UNSIGNED #(.width(7)) u_eq_624 (
        .y(_node_574),
        .a(7'd81),
        .b(__T_10__q)
    );
    wire _node_575;
    MUX_UNSIGNED #(.width(1)) u_mux_625 (
        .y(_node_575),
        .sel(_node_574),
        .a(_T_574_81),
        .b(_node_573)
    );
    wire _node_576;
    EQ_UNSIGNED #(.width(7)) u_eq_626 (
        .y(_node_576),
        .a(7'd82),
        .b(__T_10__q)
    );
    wire _node_577;
    MUX_UNSIGNED #(.width(1)) u_mux_627 (
        .y(_node_577),
        .sel(_node_576),
        .a(_T_574_82),
        .b(_node_575)
    );
    wire _node_578;
    EQ_UNSIGNED #(.width(7)) u_eq_628 (
        .y(_node_578),
        .a(7'd83),
        .b(__T_10__q)
    );
    wire _node_579;
    MUX_UNSIGNED #(.width(1)) u_mux_629 (
        .y(_node_579),
        .sel(_node_578),
        .a(_T_574_83),
        .b(_node_577)
    );
    wire _node_580;
    EQ_UNSIGNED #(.width(7)) u_eq_630 (
        .y(_node_580),
        .a(7'd84),
        .b(__T_10__q)
    );
    wire _node_581;
    MUX_UNSIGNED #(.width(1)) u_mux_631 (
        .y(_node_581),
        .sel(_node_580),
        .a(_T_574_84),
        .b(_node_579)
    );
    wire _node_582;
    EQ_UNSIGNED #(.width(7)) u_eq_632 (
        .y(_node_582),
        .a(7'd85),
        .b(__T_10__q)
    );
    wire _node_583;
    MUX_UNSIGNED #(.width(1)) u_mux_633 (
        .y(_node_583),
        .sel(_node_582),
        .a(_T_574_85),
        .b(_node_581)
    );
    wire _node_584;
    EQ_UNSIGNED #(.width(7)) u_eq_634 (
        .y(_node_584),
        .a(7'd86),
        .b(__T_10__q)
    );
    wire _node_585;
    MUX_UNSIGNED #(.width(1)) u_mux_635 (
        .y(_node_585),
        .sel(_node_584),
        .a(_T_574_86),
        .b(_node_583)
    );
    wire _node_586;
    EQ_UNSIGNED #(.width(7)) u_eq_636 (
        .y(_node_586),
        .a(7'd87),
        .b(__T_10__q)
    );
    wire _node_587;
    MUX_UNSIGNED #(.width(1)) u_mux_637 (
        .y(_node_587),
        .sel(_node_586),
        .a(_T_574_87),
        .b(_node_585)
    );
    wire _node_588;
    EQ_UNSIGNED #(.width(7)) u_eq_638 (
        .y(_node_588),
        .a(7'd88),
        .b(__T_10__q)
    );
    wire _node_589;
    MUX_UNSIGNED #(.width(1)) u_mux_639 (
        .y(_node_589),
        .sel(_node_588),
        .a(_T_574_88),
        .b(_node_587)
    );
    wire _node_590;
    EQ_UNSIGNED #(.width(7)) u_eq_640 (
        .y(_node_590),
        .a(7'd89),
        .b(__T_10__q)
    );
    wire _node_591;
    MUX_UNSIGNED #(.width(1)) u_mux_641 (
        .y(_node_591),
        .sel(_node_590),
        .a(_T_574_89),
        .b(_node_589)
    );
    wire _node_592;
    EQ_UNSIGNED #(.width(7)) u_eq_642 (
        .y(_node_592),
        .a(7'd90),
        .b(__T_10__q)
    );
    wire _node_593;
    MUX_UNSIGNED #(.width(1)) u_mux_643 (
        .y(_node_593),
        .sel(_node_592),
        .a(_T_574_90),
        .b(_node_591)
    );
    wire _node_594;
    EQ_UNSIGNED #(.width(7)) u_eq_644 (
        .y(_node_594),
        .a(7'd91),
        .b(__T_10__q)
    );
    wire _node_595;
    MUX_UNSIGNED #(.width(1)) u_mux_645 (
        .y(_node_595),
        .sel(_node_594),
        .a(_T_574_91),
        .b(_node_593)
    );
    wire _node_596;
    EQ_UNSIGNED #(.width(7)) u_eq_646 (
        .y(_node_596),
        .a(7'd92),
        .b(__T_10__q)
    );
    wire _node_597;
    MUX_UNSIGNED #(.width(1)) u_mux_647 (
        .y(_node_597),
        .sel(_node_596),
        .a(_T_574_92),
        .b(_node_595)
    );
    wire _node_598;
    EQ_UNSIGNED #(.width(7)) u_eq_648 (
        .y(_node_598),
        .a(7'd93),
        .b(__T_10__q)
    );
    wire _node_599;
    MUX_UNSIGNED #(.width(1)) u_mux_649 (
        .y(_node_599),
        .sel(_node_598),
        .a(_T_574_93),
        .b(_node_597)
    );
    wire _node_600;
    EQ_UNSIGNED #(.width(7)) u_eq_650 (
        .y(_node_600),
        .a(7'd94),
        .b(__T_10__q)
    );
    wire _node_601;
    MUX_UNSIGNED #(.width(1)) u_mux_651 (
        .y(_node_601),
        .sel(_node_600),
        .a(_T_574_94),
        .b(_node_599)
    );
    wire _node_602;
    EQ_UNSIGNED #(.width(7)) u_eq_652 (
        .y(_node_602),
        .a(7'd95),
        .b(__T_10__q)
    );
    wire _node_603;
    MUX_UNSIGNED #(.width(1)) u_mux_653 (
        .y(_node_603),
        .sel(_node_602),
        .a(_T_574_95),
        .b(_node_601)
    );
    wire _node_604;
    EQ_UNSIGNED #(.width(7)) u_eq_654 (
        .y(_node_604),
        .a(7'd96),
        .b(__T_10__q)
    );
    wire _node_605;
    MUX_UNSIGNED #(.width(1)) u_mux_655 (
        .y(_node_605),
        .sel(_node_604),
        .a(_T_574_96),
        .b(_node_603)
    );
    wire _node_606;
    EQ_UNSIGNED #(.width(7)) u_eq_656 (
        .y(_node_606),
        .a(7'd97),
        .b(__T_10__q)
    );
    wire _node_607;
    MUX_UNSIGNED #(.width(1)) u_mux_657 (
        .y(_node_607),
        .sel(_node_606),
        .a(_T_574_97),
        .b(_node_605)
    );
    wire _node_608;
    EQ_UNSIGNED #(.width(7)) u_eq_658 (
        .y(_node_608),
        .a(7'd98),
        .b(__T_10__q)
    );
    wire _node_609;
    MUX_UNSIGNED #(.width(1)) u_mux_659 (
        .y(_node_609),
        .sel(_node_608),
        .a(_T_574_98),
        .b(_node_607)
    );
    wire _node_610;
    EQ_UNSIGNED #(.width(7)) u_eq_660 (
        .y(_node_610),
        .a(7'd99),
        .b(__T_10__q)
    );
    wire _node_611;
    MUX_UNSIGNED #(.width(1)) u_mux_661 (
        .y(_node_611),
        .sel(_node_610),
        .a(_T_574_99),
        .b(_node_609)
    );
    wire _node_612;
    EQ_UNSIGNED #(.width(7)) u_eq_662 (
        .y(_node_612),
        .a(7'd100),
        .b(__T_10__q)
    );
    wire _node_613;
    MUX_UNSIGNED #(.width(1)) u_mux_663 (
        .y(_node_613),
        .sel(_node_612),
        .a(_T_574_100),
        .b(_node_611)
    );
    wire _node_614;
    EQ_UNSIGNED #(.width(7)) u_eq_664 (
        .y(_node_614),
        .a(7'd101),
        .b(__T_10__q)
    );
    wire _node_615;
    MUX_UNSIGNED #(.width(1)) u_mux_665 (
        .y(_node_615),
        .sel(_node_614),
        .a(_T_574_101),
        .b(_node_613)
    );
    wire _T_743;
    BITWISEAND #(.width(1)) bitwiseand_666 (
        .y(_T_743),
        .a(_device_under_test__io_out_ready),
        .b(_device_under_test__io_out_valid)
    );
    wire _T_746;
    EQ_UNSIGNED #(.width(1)) u_eq_667 (
        .y(_T_746),
        .a(reset),
        .b(1'h0)
    );
    wire _node_616;
    EQ_UNSIGNED #(.width(5)) u_eq_668 (
        .y(_node_616),
        .a(5'd0),
        .b(_value_1__q)
    );
    wire [3:0] _node_617;
    assign _node_617 = _T_711_0;
    wire _node_618;
    EQ_UNSIGNED #(.width(5)) u_eq_669 (
        .y(_node_618),
        .a(5'd1),
        .b(_value_1__q)
    );
    wire [3:0] _node_619;
    MUX_UNSIGNED #(.width(4)) u_mux_670 (
        .y(_node_619),
        .sel(_node_618),
        .a(_T_711_1),
        .b(_node_617)
    );
    wire _node_620;
    EQ_UNSIGNED #(.width(5)) u_eq_671 (
        .y(_node_620),
        .a(5'd2),
        .b(_value_1__q)
    );
    wire [3:0] _node_621;
    MUX_UNSIGNED #(.width(4)) u_mux_672 (
        .y(_node_621),
        .sel(_node_620),
        .a(_T_711_2),
        .b(_node_619)
    );
    wire _node_622;
    EQ_UNSIGNED #(.width(5)) u_eq_673 (
        .y(_node_622),
        .a(5'd3),
        .b(_value_1__q)
    );
    wire [3:0] _node_623;
    MUX_UNSIGNED #(.width(4)) u_mux_674 (
        .y(_node_623),
        .sel(_node_622),
        .a(_T_711_3),
        .b(_node_621)
    );
    wire _node_624;
    EQ_UNSIGNED #(.width(5)) u_eq_675 (
        .y(_node_624),
        .a(5'd4),
        .b(_value_1__q)
    );
    wire [3:0] _node_625;
    MUX_UNSIGNED #(.width(4)) u_mux_676 (
        .y(_node_625),
        .sel(_node_624),
        .a(_T_711_4),
        .b(_node_623)
    );
    wire _node_626;
    EQ_UNSIGNED #(.width(5)) u_eq_677 (
        .y(_node_626),
        .a(5'd5),
        .b(_value_1__q)
    );
    wire [3:0] _node_627;
    MUX_UNSIGNED #(.width(4)) u_mux_678 (
        .y(_node_627),
        .sel(_node_626),
        .a(_T_711_5),
        .b(_node_625)
    );
    wire _node_628;
    EQ_UNSIGNED #(.width(5)) u_eq_679 (
        .y(_node_628),
        .a(5'd6),
        .b(_value_1__q)
    );
    wire [3:0] _node_629;
    MUX_UNSIGNED #(.width(4)) u_mux_680 (
        .y(_node_629),
        .sel(_node_628),
        .a(_T_711_6),
        .b(_node_627)
    );
    wire _node_630;
    EQ_UNSIGNED #(.width(5)) u_eq_681 (
        .y(_node_630),
        .a(5'd7),
        .b(_value_1__q)
    );
    wire [3:0] _node_631;
    MUX_UNSIGNED #(.width(4)) u_mux_682 (
        .y(_node_631),
        .sel(_node_630),
        .a(_T_711_7),
        .b(_node_629)
    );
    wire _node_632;
    EQ_UNSIGNED #(.width(5)) u_eq_683 (
        .y(_node_632),
        .a(5'd8),
        .b(_value_1__q)
    );
    wire [3:0] _node_633;
    MUX_UNSIGNED #(.width(4)) u_mux_684 (
        .y(_node_633),
        .sel(_node_632),
        .a(_T_711_8),
        .b(_node_631)
    );
    wire _node_634;
    EQ_UNSIGNED #(.width(5)) u_eq_685 (
        .y(_node_634),
        .a(5'd9),
        .b(_value_1__q)
    );
    wire [3:0] _node_635;
    MUX_UNSIGNED #(.width(4)) u_mux_686 (
        .y(_node_635),
        .sel(_node_634),
        .a(_T_711_9),
        .b(_node_633)
    );
    wire _node_636;
    EQ_UNSIGNED #(.width(5)) u_eq_687 (
        .y(_node_636),
        .a(5'd10),
        .b(_value_1__q)
    );
    wire [3:0] _node_637;
    MUX_UNSIGNED #(.width(4)) u_mux_688 (
        .y(_node_637),
        .sel(_node_636),
        .a(_T_711_10),
        .b(_node_635)
    );
    wire _node_638;
    EQ_UNSIGNED #(.width(5)) u_eq_689 (
        .y(_node_638),
        .a(5'd11),
        .b(_value_1__q)
    );
    wire [3:0] _node_639;
    MUX_UNSIGNED #(.width(4)) u_mux_690 (
        .y(_node_639),
        .sel(_node_638),
        .a(_T_711_11),
        .b(_node_637)
    );
    wire _node_640;
    EQ_UNSIGNED #(.width(5)) u_eq_691 (
        .y(_node_640),
        .a(5'd12),
        .b(_value_1__q)
    );
    wire [3:0] _node_641;
    MUX_UNSIGNED #(.width(4)) u_mux_692 (
        .y(_node_641),
        .sel(_node_640),
        .a(_T_711_12),
        .b(_node_639)
    );
    wire _node_642;
    EQ_UNSIGNED #(.width(5)) u_eq_693 (
        .y(_node_642),
        .a(5'd13),
        .b(_value_1__q)
    );
    wire [3:0] _node_643;
    MUX_UNSIGNED #(.width(4)) u_mux_694 (
        .y(_node_643),
        .sel(_node_642),
        .a(_T_711_13),
        .b(_node_641)
    );
    wire _node_644;
    EQ_UNSIGNED #(.width(5)) u_eq_695 (
        .y(_node_644),
        .a(5'd14),
        .b(_value_1__q)
    );
    wire [3:0] _node_645;
    MUX_UNSIGNED #(.width(4)) u_mux_696 (
        .y(_node_645),
        .sel(_node_644),
        .a(_T_711_14),
        .b(_node_643)
    );
    wire _node_646;
    EQ_UNSIGNED #(.width(5)) u_eq_697 (
        .y(_node_646),
        .a(5'd15),
        .b(_value_1__q)
    );
    wire [3:0] _node_647;
    MUX_UNSIGNED #(.width(4)) u_mux_698 (
        .y(_node_647),
        .sel(_node_646),
        .a(_T_711_15),
        .b(_node_645)
    );
    wire _node_648;
    EQ_UNSIGNED #(.width(5)) u_eq_699 (
        .y(_node_648),
        .a(5'd16),
        .b(_value_1__q)
    );
    wire [3:0] _node_649;
    MUX_UNSIGNED #(.width(4)) u_mux_700 (
        .y(_node_649),
        .sel(_node_648),
        .a(_T_711_16),
        .b(_node_647)
    );
    wire _node_650;
    EQ_UNSIGNED #(.width(5)) u_eq_701 (
        .y(_node_650),
        .a(5'd17),
        .b(_value_1__q)
    );
    wire [3:0] _node_651;
    MUX_UNSIGNED #(.width(4)) u_mux_702 (
        .y(_node_651),
        .sel(_node_650),
        .a(_T_711_17),
        .b(_node_649)
    );
    wire _node_652;
    EQ_UNSIGNED #(.width(5)) u_eq_703 (
        .y(_node_652),
        .a(5'd18),
        .b(_value_1__q)
    );
    wire [3:0] _node_653;
    MUX_UNSIGNED #(.width(4)) u_mux_704 (
        .y(_node_653),
        .sel(_node_652),
        .a(_T_711_18),
        .b(_node_651)
    );
    wire _node_654;
    EQ_UNSIGNED #(.width(5)) u_eq_705 (
        .y(_node_654),
        .a(5'd19),
        .b(_value_1__q)
    );
    wire [3:0] _node_655;
    MUX_UNSIGNED #(.width(4)) u_mux_706 (
        .y(_node_655),
        .sel(_node_654),
        .a(_T_711_19),
        .b(_node_653)
    );
    wire _node_656;
    EQ_UNSIGNED #(.width(5)) u_eq_707 (
        .y(_node_656),
        .a(5'd20),
        .b(_value_1__q)
    );
    wire [3:0] _node_657;
    MUX_UNSIGNED #(.width(4)) u_mux_708 (
        .y(_node_657),
        .sel(_node_656),
        .a(_T_711_20),
        .b(_node_655)
    );
    wire _node_658;
    EQ_UNSIGNED #(.width(5)) u_eq_709 (
        .y(_node_658),
        .a(5'd21),
        .b(_value_1__q)
    );
    wire [3:0] _node_659;
    MUX_UNSIGNED #(.width(4)) u_mux_710 (
        .y(_node_659),
        .sel(_node_658),
        .a(_T_711_21),
        .b(_node_657)
    );
    wire _node_660;
    EQ_UNSIGNED #(.width(5)) u_eq_711 (
        .y(_node_660),
        .a(5'd22),
        .b(_value_1__q)
    );
    wire [3:0] _node_661;
    MUX_UNSIGNED #(.width(4)) u_mux_712 (
        .y(_node_661),
        .sel(_node_660),
        .a(_T_711_22),
        .b(_node_659)
    );
    wire _node_662;
    EQ_UNSIGNED #(.width(5)) u_eq_713 (
        .y(_node_662),
        .a(5'd23),
        .b(_value_1__q)
    );
    wire [3:0] _node_663;
    MUX_UNSIGNED #(.width(4)) u_mux_714 (
        .y(_node_663),
        .sel(_node_662),
        .a(_T_711_23),
        .b(_node_661)
    );
    wire _node_664;
    EQ_UNSIGNED #(.width(5)) u_eq_715 (
        .y(_node_664),
        .a(5'd24),
        .b(_value_1__q)
    );
    wire [3:0] _node_665;
    MUX_UNSIGNED #(.width(4)) u_mux_716 (
        .y(_node_665),
        .sel(_node_664),
        .a(_T_711_24),
        .b(_node_663)
    );
    wire _node_666;
    EQ_UNSIGNED #(.width(5)) u_eq_717 (
        .y(_node_666),
        .a(5'd25),
        .b(_value_1__q)
    );
    wire [3:0] _node_667;
    MUX_UNSIGNED #(.width(4)) u_mux_718 (
        .y(_node_667),
        .sel(_node_666),
        .a(_T_711_25),
        .b(_node_665)
    );
    wire _node_668;
    EQ_UNSIGNED #(.width(5)) u_eq_719 (
        .y(_node_668),
        .a(5'd26),
        .b(_value_1__q)
    );
    wire [3:0] _node_669;
    MUX_UNSIGNED #(.width(4)) u_mux_720 (
        .y(_node_669),
        .sel(_node_668),
        .a(_T_711_26),
        .b(_node_667)
    );
    wire _node_670;
    EQ_UNSIGNED #(.width(5)) u_eq_721 (
        .y(_node_670),
        .a(5'd27),
        .b(_value_1__q)
    );
    wire [3:0] _node_671;
    MUX_UNSIGNED #(.width(4)) u_mux_722 (
        .y(_node_671),
        .sel(_node_670),
        .a(_T_711_27),
        .b(_node_669)
    );
    wire _T_748;
    wire [31:0] _WTEMP_16;
    PAD_UNSIGNED #(.width(4), .n(32)) u_pad_723 (
        .y(_WTEMP_16),
        .in(_node_671)
    );
    NEQ_UNSIGNED #(.width(32)) u_neq_724 (
        .y(_T_748),
        .a(_device_under_test__io_out_bits),
        .b(_WTEMP_16)
    );
    wire _T_751;
    EQ_UNSIGNED #(.width(1)) u_eq_725 (
        .y(_T_751),
        .a(reset),
        .b(1'h0)
    );
    wire _T_753;
    BITWISEOR #(.width(1)) bitwiseor_726 (
        .y(_T_753),
        .a(1'h0),
        .b(reset)
    );
    wire _T_755;
    EQ_UNSIGNED #(.width(1)) u_eq_727 (
        .y(_T_755),
        .a(_T_753),
        .b(1'h0)
    );
    wire _T_757;
    EQ_UNSIGNED #(.width(1)) u_eq_728 (
        .y(_T_757),
        .a(reset),
        .b(1'h0)
    );
    wire _T_759;
    EQ_UNSIGNED #(.width(5)) u_eq_729 (
        .y(_T_759),
        .a(_value_1__q),
        .b(5'h1A)
    );
    wire [5:0] _T_761;
    wire [4:0] _WTEMP_17;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_730 (
        .y(_WTEMP_17),
        .in(1'h1)
    );
    ADD_UNSIGNED #(.width(5)) u_add_731 (
        .y(_T_761),
        .a(_value_1__q),
        .b(_WTEMP_17)
    );
    wire [4:0] _T_762;
    TAIL #(.width(6), .n(1)) tail_732 (
        .y(_T_762),
        .in(_T_761)
    );
    wire _T_765;
    EQ_UNSIGNED #(.width(1)) u_eq_733 (
        .y(_T_765),
        .a(__T_13__q),
        .b(1'h0)
    );
    wire _T_767;
    wire [6:0] _WTEMP_18;
    PAD_UNSIGNED #(.width(5), .n(7)) u_pad_734 (
        .y(_WTEMP_18),
        .in(5'h1A)
    );
    EQ_UNSIGNED #(.width(7)) u_eq_735 (
        .y(_T_767),
        .a(__T_10__q),
        .b(_WTEMP_18)
    );
    wire [7:0] _T_770;
    wire [6:0] _WTEMP_19;
    PAD_UNSIGNED #(.width(1), .n(7)) u_pad_736 (
        .y(_WTEMP_19),
        .in(1'h1)
    );
    ADD_UNSIGNED #(.width(7)) u_add_737 (
        .y(_T_770),
        .a(__T_10__q),
        .b(_WTEMP_19)
    );
    wire [6:0] _T_771;
    TAIL #(.width(8), .n(1)) tail_738 (
        .y(_T_771),
        .in(_T_770)
    );
    wire _node_672;
    MUX_UNSIGNED #(.width(1)) u_mux_739 (
        .y(_node_672),
        .sel(_T_767),
        .a(1'h1),
        .b(__T_13__q)
    );
    wire [6:0] _node_673;
    MUX_UNSIGNED #(.width(7)) u_mux_740 (
        .y(_node_673),
        .sel(_T_765),
        .a(_T_771),
        .b(__T_10__q)
    );
    wire _node_674;
    MUX_UNSIGNED #(.width(1)) u_mux_741 (
        .y(_node_674),
        .sel(_T_765),
        .a(_node_672),
        .b(__T_13__q)
    );
    wire [4:0] _node_675;
    wire [4:0] _WTEMP_20;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_742 (
        .y(_WTEMP_20),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(5)) u_mux_743 (
        .y(_node_675),
        .sel(_T_759),
        .a(_WTEMP_20),
        .b(_T_762)
    );
    MUX_UNSIGNED #(.width(7)) u_mux_744 (
        .y(_WTEMP_6),
        .sel(_T_743),
        .a(_node_673),
        .b(__T_10__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_745 (
        .y(_WTEMP_7),
        .sel(_T_743),
        .a(_node_674),
        .b(__T_13__q)
    );
    assign _T_136_0 = 1'h1;
    assign _T_136_1 = 1'h1;
    assign _T_136_10 = 1'h1;
    assign _T_136_100 = 1'h1;
    assign _T_136_101 = 1'h0;
    assign _T_136_11 = 1'h1;
    assign _T_136_12 = 1'h1;
    assign _T_136_13 = 1'h1;
    assign _T_136_14 = 1'h1;
    assign _T_136_15 = 1'h1;
    assign _T_136_16 = 1'h1;
    assign _T_136_17 = 1'h1;
    assign _T_136_18 = 1'h1;
    assign _T_136_19 = 1'h1;
    assign _T_136_2 = 1'h1;
    assign _T_136_20 = 1'h1;
    assign _T_136_21 = 1'h1;
    assign _T_136_22 = 1'h1;
    assign _T_136_23 = 1'h1;
    assign _T_136_24 = 1'h1;
    assign _T_136_25 = 1'h1;
    assign _T_136_26 = 1'h1;
    assign _T_136_27 = 1'h1;
    assign _T_136_28 = 1'h1;
    assign _T_136_29 = 1'h1;
    assign _T_136_3 = 1'h1;
    assign _T_136_30 = 1'h1;
    assign _T_136_31 = 1'h1;
    assign _T_136_32 = 1'h1;
    assign _T_136_33 = 1'h1;
    assign _T_136_34 = 1'h1;
    assign _T_136_35 = 1'h1;
    assign _T_136_36 = 1'h1;
    assign _T_136_37 = 1'h1;
    assign _T_136_38 = 1'h1;
    assign _T_136_39 = 1'h1;
    assign _T_136_4 = 1'h1;
    assign _T_136_40 = 1'h1;
    assign _T_136_41 = 1'h1;
    assign _T_136_42 = 1'h1;
    assign _T_136_43 = 1'h1;
    assign _T_136_44 = 1'h1;
    assign _T_136_45 = 1'h1;
    assign _T_136_46 = 1'h1;
    assign _T_136_47 = 1'h1;
    assign _T_136_48 = 1'h1;
    assign _T_136_49 = 1'h1;
    assign _T_136_5 = 1'h1;
    assign _T_136_50 = 1'h1;
    assign _T_136_51 = 1'h1;
    assign _T_136_52 = 1'h1;
    assign _T_136_53 = 1'h1;
    assign _T_136_54 = 1'h1;
    assign _T_136_55 = 1'h1;
    assign _T_136_56 = 1'h1;
    assign _T_136_57 = 1'h1;
    assign _T_136_58 = 1'h1;
    assign _T_136_59 = 1'h1;
    assign _T_136_6 = 1'h1;
    assign _T_136_60 = 1'h1;
    assign _T_136_61 = 1'h1;
    assign _T_136_62 = 1'h1;
    assign _T_136_63 = 1'h1;
    assign _T_136_64 = 1'h1;
    assign _T_136_65 = 1'h1;
    assign _T_136_66 = 1'h1;
    assign _T_136_67 = 1'h1;
    assign _T_136_68 = 1'h1;
    assign _T_136_69 = 1'h1;
    assign _T_136_7 = 1'h1;
    assign _T_136_70 = 1'h1;
    assign _T_136_71 = 1'h1;
    assign _T_136_72 = 1'h1;
    assign _T_136_73 = 1'h1;
    assign _T_136_74 = 1'h1;
    assign _T_136_75 = 1'h1;
    assign _T_136_76 = 1'h1;
    assign _T_136_77 = 1'h1;
    assign _T_136_78 = 1'h1;
    assign _T_136_79 = 1'h1;
    assign _T_136_8 = 1'h1;
    assign _T_136_80 = 1'h1;
    assign _T_136_81 = 1'h1;
    assign _T_136_82 = 1'h1;
    assign _T_136_83 = 1'h1;
    assign _T_136_84 = 1'h1;
    assign _T_136_85 = 1'h1;
    assign _T_136_86 = 1'h1;
    assign _T_136_87 = 1'h1;
    assign _T_136_88 = 1'h1;
    assign _T_136_89 = 1'h1;
    assign _T_136_9 = 1'h1;
    assign _T_136_90 = 1'h1;
    assign _T_136_91 = 1'h1;
    assign _T_136_92 = 1'h1;
    assign _T_136_93 = 1'h1;
    assign _T_136_94 = 1'h1;
    assign _T_136_95 = 1'h1;
    assign _T_136_96 = 1'h1;
    assign _T_136_97 = 1'h1;
    assign _T_136_98 = 1'h1;
    assign _T_136_99 = 1'h1;
    assign _WTEMP_8 = _T_24;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_746 (
        .y(_T_347_0),
        .in(1'h0)
    );
    PAD_UNSIGNED #(.width(4), .n(5)) u_pad_747 (
        .y(_T_347_1),
        .in(4'h8)
    );
    assign _T_347_10 = 5'h11;
    assign _T_347_100 = 5'h10;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_748 (
        .y(_T_347_101),
        .in(1'h0)
    );
    assign _T_347_11 = 5'h11;
    PAD_UNSIGNED #(.width(4), .n(5)) u_pad_749 (
        .y(_T_347_12),
        .in(4'hD)
    );
    PAD_UNSIGNED #(.width(2), .n(5)) u_pad_750 (
        .y(_T_347_13),
        .in(2'h2)
    );
    PAD_UNSIGNED #(.width(4), .n(5)) u_pad_751 (
        .y(_T_347_14),
        .in(4'hF)
    );
    PAD_UNSIGNED #(.width(3), .n(5)) u_pad_752 (
        .y(_T_347_15),
        .in(3'h4)
    );
    PAD_UNSIGNED #(.width(3), .n(5)) u_pad_753 (
        .y(_T_347_16),
        .in(3'h4)
    );
    PAD_UNSIGNED #(.width(4), .n(5)) u_pad_754 (
        .y(_T_347_17),
        .in(4'hF)
    );
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_755 (
        .y(_T_347_18),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_756 (
        .y(_T_347_19),
        .in(1'h0)
    );
    PAD_UNSIGNED #(.width(4), .n(5)) u_pad_757 (
        .y(_T_347_2),
        .in(4'h9)
    );
    PAD_UNSIGNED #(.width(2), .n(5)) u_pad_758 (
        .y(_T_347_20),
        .in(2'h3)
    );
    PAD_UNSIGNED #(.width(4), .n(5)) u_pad_759 (
        .y(_T_347_21),
        .in(4'h8)
    );
    PAD_UNSIGNED #(.width(3), .n(5)) u_pad_760 (
        .y(_T_347_22),
        .in(3'h4)
    );
    PAD_UNSIGNED #(.width(3), .n(5)) u_pad_761 (
        .y(_T_347_23),
        .in(3'h7)
    );
    PAD_UNSIGNED #(.width(4), .n(5)) u_pad_762 (
        .y(_T_347_24),
        .in(4'hC)
    );
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_763 (
        .y(_T_347_25),
        .in(1'h0)
    );
    PAD_UNSIGNED #(.width(2), .n(5)) u_pad_764 (
        .y(_T_347_26),
        .in(2'h3)
    );
    PAD_UNSIGNED #(.width(2), .n(5)) u_pad_765 (
        .y(_T_347_27),
        .in(2'h2)
    );
    PAD_UNSIGNED #(.width(4), .n(5)) u_pad_766 (
        .y(_T_347_28),
        .in(4'hC)
    );
    PAD_UNSIGNED #(.width(2), .n(5)) u_pad_767 (
        .y(_T_347_29),
        .in(2'h3)
    );
    PAD_UNSIGNED #(.width(3), .n(5)) u_pad_768 (
        .y(_T_347_3),
        .in(3'h7)
    );
    PAD_UNSIGNED #(.width(3), .n(5)) u_pad_769 (
        .y(_T_347_30),
        .in(3'h5)
    );
    PAD_UNSIGNED #(.width(3), .n(5)) u_pad_770 (
        .y(_T_347_31),
        .in(3'h5)
    );
    assign _T_347_32 = 5'h11;
    PAD_UNSIGNED #(.width(3), .n(5)) u_pad_771 (
        .y(_T_347_33),
        .in(3'h7)
    );
    PAD_UNSIGNED #(.width(2), .n(5)) u_pad_772 (
        .y(_T_347_34),
        .in(2'h2)
    );
    PAD_UNSIGNED #(.width(2), .n(5)) u_pad_773 (
        .y(_T_347_35),
        .in(2'h2)
    );
    PAD_UNSIGNED #(.width(3), .n(5)) u_pad_774 (
        .y(_T_347_36),
        .in(3'h5)
    );
    PAD_UNSIGNED #(.width(4), .n(5)) u_pad_775 (
        .y(_T_347_37),
        .in(4'hD)
    );
    assign _T_347_38 = 5'h12;
    PAD_UNSIGNED #(.width(4), .n(5)) u_pad_776 (
        .y(_T_347_39),
        .in(4'hF)
    );
    PAD_UNSIGNED #(.width(4), .n(5)) u_pad_777 (
        .y(_T_347_4),
        .in(4'hF)
    );
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_778 (
        .y(_T_347_40),
        .in(1'h0)
    );
    PAD_UNSIGNED #(.width(4), .n(5)) u_pad_779 (
        .y(_T_347_41),
        .in(4'hF)
    );
    PAD_UNSIGNED #(.width(4), .n(5)) u_pad_780 (
        .y(_T_347_42),
        .in(4'hF)
    );
    PAD_UNSIGNED #(.width(4), .n(5)) u_pad_781 (
        .y(_T_347_43),
        .in(4'hA)
    );
    assign _T_347_44 = 5'h12;
    PAD_UNSIGNED #(.width(4), .n(5)) u_pad_782 (
        .y(_T_347_45),
        .in(4'hB)
    );
    PAD_UNSIGNED #(.width(4), .n(5)) u_pad_783 (
        .y(_T_347_46),
        .in(4'hE)
    );
    assign _T_347_47 = 5'h10;
    PAD_UNSIGNED #(.width(4), .n(5)) u_pad_784 (
        .y(_T_347_48),
        .in(4'hC)
    );
    PAD_UNSIGNED #(.width(2), .n(5)) u_pad_785 (
        .y(_T_347_49),
        .in(2'h2)
    );
    PAD_UNSIGNED #(.width(4), .n(5)) u_pad_786 (
        .y(_T_347_5),
        .in(4'hD)
    );
    assign _T_347_50 = 5'h13;
    assign _T_347_51 = 5'h11;
    assign _T_347_52 = 5'h10;
    PAD_UNSIGNED #(.width(3), .n(5)) u_pad_787 (
        .y(_T_347_53),
        .in(3'h6)
    );
    PAD_UNSIGNED #(.width(3), .n(5)) u_pad_788 (
        .y(_T_347_54),
        .in(3'h7)
    );
    assign _T_347_55 = 5'h10;
    PAD_UNSIGNED #(.width(4), .n(5)) u_pad_789 (
        .y(_T_347_56),
        .in(4'h8)
    );
    assign _T_347_57 = 5'h11;
    PAD_UNSIGNED #(.width(2), .n(5)) u_pad_790 (
        .y(_T_347_58),
        .in(2'h3)
    );
    PAD_UNSIGNED #(.width(3), .n(5)) u_pad_791 (
        .y(_T_347_59),
        .in(3'h7)
    );
    PAD_UNSIGNED #(.width(4), .n(5)) u_pad_792 (
        .y(_T_347_6),
        .in(4'hB)
    );
    PAD_UNSIGNED #(.width(3), .n(5)) u_pad_793 (
        .y(_T_347_60),
        .in(3'h7)
    );
    PAD_UNSIGNED #(.width(4), .n(5)) u_pad_794 (
        .y(_T_347_61),
        .in(4'h8)
    );
    PAD_UNSIGNED #(.width(3), .n(5)) u_pad_795 (
        .y(_T_347_62),
        .in(3'h5)
    );
    assign _T_347_63 = 5'h12;
    PAD_UNSIGNED #(.width(4), .n(5)) u_pad_796 (
        .y(_T_347_64),
        .in(4'h8)
    );
    assign _T_347_65 = 5'h11;
    PAD_UNSIGNED #(.width(4), .n(5)) u_pad_797 (
        .y(_T_347_66),
        .in(4'hB)
    );
    assign _T_347_67 = 5'h12;
    assign _T_347_68 = 5'h12;
    assign _T_347_69 = 5'h12;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_798 (
        .y(_T_347_7),
        .in(1'h1)
    );
    assign _T_347_70 = 5'h12;
    PAD_UNSIGNED #(.width(4), .n(5)) u_pad_799 (
        .y(_T_347_71),
        .in(4'hC)
    );
    assign _T_347_72 = 5'h11;
    PAD_UNSIGNED #(.width(4), .n(5)) u_pad_800 (
        .y(_T_347_73),
        .in(4'hB)
    );
    PAD_UNSIGNED #(.width(3), .n(5)) u_pad_801 (
        .y(_T_347_74),
        .in(3'h6)
    );
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_802 (
        .y(_T_347_75),
        .in(1'h0)
    );
    assign _T_347_76 = 5'h11;
    PAD_UNSIGNED #(.width(2), .n(5)) u_pad_803 (
        .y(_T_347_77),
        .in(2'h2)
    );
    PAD_UNSIGNED #(.width(4), .n(5)) u_pad_804 (
        .y(_T_347_78),
        .in(4'hF)
    );
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_805 (
        .y(_T_347_79),
        .in(1'h0)
    );
    assign _T_347_8 = 5'h13;
    PAD_UNSIGNED #(.width(3), .n(5)) u_pad_806 (
        .y(_T_347_80),
        .in(3'h7)
    );
    PAD_UNSIGNED #(.width(4), .n(5)) u_pad_807 (
        .y(_T_347_81),
        .in(4'hD)
    );
    assign _T_347_82 = 5'h11;
    PAD_UNSIGNED #(.width(4), .n(5)) u_pad_808 (
        .y(_T_347_83),
        .in(4'h9)
    );
    PAD_UNSIGNED #(.width(3), .n(5)) u_pad_809 (
        .y(_T_347_84),
        .in(3'h5)
    );
    PAD_UNSIGNED #(.width(4), .n(5)) u_pad_810 (
        .y(_T_347_85),
        .in(4'hC)
    );
    PAD_UNSIGNED #(.width(4), .n(5)) u_pad_811 (
        .y(_T_347_86),
        .in(4'h9)
    );
    PAD_UNSIGNED #(.width(2), .n(5)) u_pad_812 (
        .y(_T_347_87),
        .in(2'h3)
    );
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_813 (
        .y(_T_347_88),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_814 (
        .y(_T_347_89),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(4), .n(5)) u_pad_815 (
        .y(_T_347_9),
        .in(4'hE)
    );
    PAD_UNSIGNED #(.width(2), .n(5)) u_pad_816 (
        .y(_T_347_90),
        .in(2'h3)
    );
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_817 (
        .y(_T_347_91),
        .in(1'h0)
    );
    PAD_UNSIGNED #(.width(4), .n(5)) u_pad_818 (
        .y(_T_347_92),
        .in(4'h8)
    );
    PAD_UNSIGNED #(.width(4), .n(5)) u_pad_819 (
        .y(_T_347_93),
        .in(4'hE)
    );
    assign _T_347_94 = 5'h10;
    PAD_UNSIGNED #(.width(2), .n(5)) u_pad_820 (
        .y(_T_347_95),
        .in(2'h3)
    );
    assign _T_347_96 = 5'h11;
    PAD_UNSIGNED #(.width(2), .n(5)) u_pad_821 (
        .y(_T_347_97),
        .in(2'h2)
    );
    PAD_UNSIGNED #(.width(3), .n(5)) u_pad_822 (
        .y(_T_347_98),
        .in(3'h5)
    );
    PAD_UNSIGNED #(.width(4), .n(5)) u_pad_823 (
        .y(_T_347_99),
        .in(4'hB)
    );
    MUX_UNSIGNED #(.width(9)) u_mux_824 (
        .y(_WTEMP_4),
        .sel(_T_455),
        .a(_node_409),
        .b(__T_4__q)
    );
    assign _T_574_0 = 1'h1;
    assign _T_574_1 = 1'h1;
    assign _T_574_10 = 1'h1;
    assign _T_574_100 = 1'h0;
    assign _T_574_101 = 1'h0;
    assign _T_574_11 = 1'h1;
    assign _T_574_12 = 1'h1;
    assign _T_574_13 = 1'h1;
    assign _T_574_14 = 1'h1;
    assign _T_574_15 = 1'h1;
    assign _T_574_16 = 1'h1;
    assign _T_574_17 = 1'h1;
    assign _T_574_18 = 1'h1;
    assign _T_574_19 = 1'h1;
    assign _T_574_2 = 1'h1;
    assign _T_574_20 = 1'h1;
    assign _T_574_21 = 1'h1;
    assign _T_574_22 = 1'h1;
    assign _T_574_23 = 1'h1;
    assign _T_574_24 = 1'h1;
    assign _T_574_25 = 1'h1;
    assign _T_574_26 = 1'h1;
    assign _T_574_27 = 1'h0;
    assign _T_574_28 = 1'h0;
    assign _T_574_29 = 1'h0;
    assign _T_574_3 = 1'h1;
    assign _T_574_30 = 1'h0;
    assign _T_574_31 = 1'h0;
    assign _T_574_32 = 1'h0;
    assign _T_574_33 = 1'h0;
    assign _T_574_34 = 1'h0;
    assign _T_574_35 = 1'h0;
    assign _T_574_36 = 1'h0;
    assign _T_574_37 = 1'h0;
    assign _T_574_38 = 1'h0;
    assign _T_574_39 = 1'h0;
    assign _T_574_4 = 1'h1;
    assign _T_574_40 = 1'h0;
    assign _T_574_41 = 1'h0;
    assign _T_574_42 = 1'h0;
    assign _T_574_43 = 1'h0;
    assign _T_574_44 = 1'h0;
    assign _T_574_45 = 1'h0;
    assign _T_574_46 = 1'h0;
    assign _T_574_47 = 1'h0;
    assign _T_574_48 = 1'h0;
    assign _T_574_49 = 1'h0;
    assign _T_574_5 = 1'h1;
    assign _T_574_50 = 1'h0;
    assign _T_574_51 = 1'h0;
    assign _T_574_52 = 1'h0;
    assign _T_574_53 = 1'h0;
    assign _T_574_54 = 1'h0;
    assign _T_574_55 = 1'h0;
    assign _T_574_56 = 1'h0;
    assign _T_574_57 = 1'h0;
    assign _T_574_58 = 1'h0;
    assign _T_574_59 = 1'h0;
    assign _T_574_6 = 1'h1;
    assign _T_574_60 = 1'h0;
    assign _T_574_61 = 1'h0;
    assign _T_574_62 = 1'h0;
    assign _T_574_63 = 1'h0;
    assign _T_574_64 = 1'h0;
    assign _T_574_65 = 1'h0;
    assign _T_574_66 = 1'h0;
    assign _T_574_67 = 1'h0;
    assign _T_574_68 = 1'h0;
    assign _T_574_69 = 1'h0;
    assign _T_574_7 = 1'h1;
    assign _T_574_70 = 1'h0;
    assign _T_574_71 = 1'h0;
    assign _T_574_72 = 1'h0;
    assign _T_574_73 = 1'h0;
    assign _T_574_74 = 1'h0;
    assign _T_574_75 = 1'h0;
    assign _T_574_76 = 1'h0;
    assign _T_574_77 = 1'h0;
    assign _T_574_78 = 1'h0;
    assign _T_574_79 = 1'h0;
    assign _T_574_8 = 1'h1;
    assign _T_574_80 = 1'h0;
    assign _T_574_81 = 1'h0;
    assign _T_574_82 = 1'h0;
    assign _T_574_83 = 1'h0;
    assign _T_574_84 = 1'h0;
    assign _T_574_85 = 1'h0;
    assign _T_574_86 = 1'h0;
    assign _T_574_87 = 1'h0;
    assign _T_574_88 = 1'h0;
    assign _T_574_89 = 1'h0;
    assign _T_574_9 = 1'h1;
    assign _T_574_90 = 1'h0;
    assign _T_574_91 = 1'h0;
    assign _T_574_92 = 1'h0;
    assign _T_574_93 = 1'h0;
    assign _T_574_94 = 1'h0;
    assign _T_574_95 = 1'h0;
    assign _T_574_96 = 1'h0;
    assign _T_574_97 = 1'h0;
    assign _T_574_98 = 1'h0;
    assign _T_574_99 = 1'h0;
    MUX_UNSIGNED #(.width(1)) u_mux_825 (
        .y(_WTEMP_5),
        .sel(_T_455),
        .a(_node_410),
        .b(__T_7__q)
    );
    assign _T_711_0 = 4'h9;
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_826 (
        .y(_T_711_1),
        .in(3'h7)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_827 (
        .y(_T_711_10),
        .in(3'h7)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_828 (
        .y(_T_711_11),
        .in(3'h5)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_829 (
        .y(_T_711_12),
        .in(3'h7)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_830 (
        .y(_T_711_13),
        .in(2'h3)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_831 (
        .y(_T_711_14),
        .in(3'h7)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_832 (
        .y(_T_711_15),
        .in(3'h7)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_833 (
        .y(_T_711_16),
        .in(3'h5)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_834 (
        .y(_T_711_17),
        .in(3'h7)
    );
    assign _T_711_18 = 4'h9;
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_835 (
        .y(_T_711_19),
        .in(3'h5)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_836 (
        .y(_T_711_2),
        .in(1'h1)
    );
    assign _T_711_20 = 4'h9;
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_837 (
        .y(_T_711_21),
        .in(2'h3)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_838 (
        .y(_T_711_22),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_839 (
        .y(_T_711_23),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_840 (
        .y(_T_711_24),
        .in(2'h3)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_841 (
        .y(_T_711_25),
        .in(2'h3)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_842 (
        .y(_T_711_26),
        .in(3'h5)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_843 (
        .y(_T_711_27),
        .in(1'h0)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_844 (
        .y(_T_711_3),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_845 (
        .y(_T_711_4),
        .in(2'h3)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_846 (
        .y(_T_711_5),
        .in(3'h7)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_847 (
        .y(_T_711_6),
        .in(2'h3)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_848 (
        .y(_T_711_7),
        .in(2'h3)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_849 (
        .y(_T_711_8),
        .in(3'h5)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_850 (
        .y(_T_711_9),
        .in(3'h5)
    );
    assign _device_under_test__clock = clock;
    PAD_UNSIGNED #(.width(5), .n(32)) u_pad_851 (
        .y(_device_under_test__io_in_bits),
        .in(_node_203)
    );
    assign _device_under_test__io_in_valid = _node_407;
    assign _device_under_test__io_out_ready = _node_615;
    assign _device_under_test__reset = reset;
    MUX_UNSIGNED #(.width(7)) u_mux_852 (
        .y(_WTEMP_10),
        .sel(_T_455),
        .a(_node_411),
        .b(_value__q)
    );
    MUX_UNSIGNED #(.width(5)) u_mux_853 (
        .y(_WTEMP_15),
        .sel(_T_743),
        .a(_node_675),
        .b(_value_1__q)
    );
endmodule //SmallOdds3Tester
module SmallOdds3(
    input clock,
    input reset,
    output io_in_ready,
    input io_in_valid,
    input [31:0] io_in_bits,
    input io_out_ready,
    output io_out_valid,
    output [31:0] io_out_bits
);
    wire _SmallOdds3Filter__clock;
    wire _SmallOdds3Filter__reset;
    wire _SmallOdds3Filter__io_in_ready;
    wire _SmallOdds3Filter__io_in_valid;
    wire [31:0] _SmallOdds3Filter__io_in_bits;
    wire _SmallOdds3Filter__io_out_ready;
    wire _SmallOdds3Filter__io_out_valid;
    wire [31:0] _SmallOdds3Filter__io_out_bits;
    SmallOdds3Filter SmallOdds3Filter (
        .clock(_SmallOdds3Filter__clock),
        .reset(_SmallOdds3Filter__reset),
        .io_in_ready(_SmallOdds3Filter__io_in_ready),
        .io_in_valid(_SmallOdds3Filter__io_in_valid),
        .io_in_bits(_SmallOdds3Filter__io_in_bits),
        .io_out_ready(_SmallOdds3Filter__io_out_ready),
        .io_out_valid(_SmallOdds3Filter__io_out_valid),
        .io_out_bits(_SmallOdds3Filter__io_out_bits)
    );
    wire _Queue__clock;
    wire _Queue__reset;
    wire _Queue__io_enq_ready;
    wire _Queue__io_enq_valid;
    wire [31:0] _Queue__io_enq_bits;
    wire _Queue__io_deq_ready;
    wire _Queue__io_deq_valid;
    wire [31:0] _Queue__io_deq_bits;
    wire _Queue__io_count;
    Queue Queue (
        .clock(_Queue__clock),
        .reset(_Queue__reset),
        .io_enq_ready(_Queue__io_enq_ready),
        .io_enq_valid(_Queue__io_enq_valid),
        .io_enq_bits(_Queue__io_enq_bits),
        .io_deq_ready(_Queue__io_deq_ready),
        .io_deq_valid(_Queue__io_deq_valid),
        .io_deq_bits(_Queue__io_deq_bits),
        .io_count(_Queue__io_count)
    );
    wire _SmallOdds3Filter_1__clock;
    wire _SmallOdds3Filter_1__reset;
    wire _SmallOdds3Filter_1__io_in_ready;
    wire _SmallOdds3Filter_1__io_in_valid;
    wire [31:0] _SmallOdds3Filter_1__io_in_bits;
    wire _SmallOdds3Filter_1__io_out_ready;
    wire _SmallOdds3Filter_1__io_out_valid;
    wire [31:0] _SmallOdds3Filter_1__io_out_bits;
    SmallOdds3Filter_1 SmallOdds3Filter_1 (
        .clock(_SmallOdds3Filter_1__clock),
        .reset(_SmallOdds3Filter_1__reset),
        .io_in_ready(_SmallOdds3Filter_1__io_in_ready),
        .io_in_valid(_SmallOdds3Filter_1__io_in_valid),
        .io_in_bits(_SmallOdds3Filter_1__io_in_bits),
        .io_out_ready(_SmallOdds3Filter_1__io_out_ready),
        .io_out_valid(_SmallOdds3Filter_1__io_out_valid),
        .io_out_bits(_SmallOdds3Filter_1__io_out_bits)
    );
    assign _Queue__clock = clock;
    assign _Queue__io_deq_ready = _SmallOdds3Filter_1__io_in_ready;
    assign _Queue__io_enq_bits = _SmallOdds3Filter__io_out_bits;
    assign _Queue__io_enq_valid = _SmallOdds3Filter__io_out_valid;
    assign _Queue__reset = reset;
    assign _SmallOdds3Filter__clock = clock;
    assign _SmallOdds3Filter__io_in_bits = io_in_bits;
    assign _SmallOdds3Filter__io_in_valid = io_in_valid;
    assign _SmallOdds3Filter__io_out_ready = _Queue__io_enq_ready;
    assign _SmallOdds3Filter__reset = reset;
    assign _SmallOdds3Filter_1__clock = clock;
    assign _SmallOdds3Filter_1__io_in_bits = _Queue__io_deq_bits;
    assign _SmallOdds3Filter_1__io_in_valid = _Queue__io_deq_valid;
    assign _SmallOdds3Filter_1__io_out_ready = io_out_ready;
    assign _SmallOdds3Filter_1__reset = reset;
    assign io_in_ready = _SmallOdds3Filter__io_in_ready;
    assign io_out_bits = _SmallOdds3Filter_1__io_out_bits;
    assign io_out_valid = _SmallOdds3Filter_1__io_out_valid;
endmodule //SmallOdds3
module SmallOdds3Filter(
    input clock,
    input reset,
    output io_in_ready,
    input io_in_valid,
    input [31:0] io_in_bits,
    input io_out_ready,
    output io_out_valid,
    output [31:0] io_out_bits
);
    wire _T_14;
    BITWISEAND #(.width(1)) bitwiseand_1 (
        .y(_T_14),
        .a(io_out_ready),
        .b(io_in_valid)
    );
    wire _T_16;
    wire [31:0] _WTEMP_0;
    PAD_UNSIGNED #(.width(4), .n(32)) u_pad_2 (
        .y(_WTEMP_0),
        .in(4'hA)
    );
    LT_UNSIGNED #(.width(32)) u_lt_3 (
        .y(_T_16),
        .a(io_in_bits),
        .b(_WTEMP_0)
    );
    wire _T_17;
    BITWISEAND #(.width(1)) bitwiseand_4 (
        .y(_T_17),
        .a(_T_14),
        .b(_T_16)
    );
    assign io_in_ready = io_out_ready;
    assign io_out_bits = io_in_bits;
    assign io_out_valid = _T_17;
endmodule //SmallOdds3Filter
module BITWISEAND(y, a, b);
    parameter width = 4;
    output [width-1:0] y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a & b;
endmodule // BITWISEAND
module PAD_UNSIGNED(y, in);
    parameter width = 4;
    parameter n = 4;
    output [(n > width ? n : width)-1:0] y;
    input [width-1:0] in;
    assign y = (n > width) ? {{(n - width){1'b0}}, in} : in;
endmodule // PAD_UNSIGNED
module LT_UNSIGNED(y, a, b);
    parameter width = 4;
    output y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a < b;
endmodule // LT_UNSIGNED
module Queue(
    input clock,
    input reset,
    output io_enq_ready,
    input io_enq_valid,
    input [31:0] io_enq_bits,
    input io_deq_ready,
    output io_deq_valid,
    output [31:0] io_deq_bits,
    output io_count
);
    wire ram__T_34_clk;
    wire ram__T_34_en;
    wire ram__T_34_mask;
    wire ram__T_34_addr;
    wire [31:0] ram__T_34_data;
    wire [31:0] ram__T_43_data;
    wire ram__T_43_clk;
    wire ram__T_43_en;
    wire ram__T_43_addr;
    RAMMEM #(.depth(1), .addrbits(1), .width(32), .isSyncRead(0)) ram (
        .read_data(ram__T_43_data),
        .read_clk(ram__T_43_clk),
        .read_en(ram__T_43_en),
        .read_addr(ram__T_43_addr),
        .write_clk(ram__T_34_clk),
        .write_en(ram__T_34_en),
        .write_mask(ram__T_34_mask),
        .write_addr(ram__T_34_addr),
        .write_data(ram__T_34_data)
    );
    wire _maybe_full__q;
    wire _maybe_full__d;
    DFF_POSCLK #(.width(1)) maybe_full (
        .q(_maybe_full__q),
        .d(_maybe_full__d),
        .clk(clock)
    );
    wire _WTEMP_1;
    MUX_UNSIGNED #(.width(1)) u_mux_5 (
        .y(_maybe_full__d),
        .sel(reset),
        .a(1'h0),
        .b(_WTEMP_1)
    );
    wire _T_24;
    assign _T_24 = 1'h1;
    wire _T_26;
    EQ_UNSIGNED #(.width(1)) u_eq_6 (
        .y(_T_26),
        .a(_maybe_full__q),
        .b(1'h0)
    );
    wire _T_27;
    BITWISEAND #(.width(1)) bitwiseand_7 (
        .y(_T_27),
        .a(_T_24),
        .b(_T_26)
    );
    wire _T_28;
    BITWISEAND #(.width(1)) bitwiseand_8 (
        .y(_T_28),
        .a(_T_24),
        .b(_maybe_full__q)
    );
    wire _T_29;
    BITWISEAND #(.width(1)) bitwiseand_9 (
        .y(_T_29),
        .a(io_enq_ready),
        .b(io_enq_valid)
    );
    wire do_enq;
    wire _T_31;
    BITWISEAND #(.width(1)) bitwiseand_10 (
        .y(_T_31),
        .a(io_deq_ready),
        .b(io_deq_valid)
    );
    wire do_deq;
    assign ram__T_34_addr = 1'h0;
    assign ram__T_34_en = do_enq;
    assign ram__T_34_clk = clock;
    assign ram__T_34_mask = 1'h1;
    wire _T_37;
    NEQ_UNSIGNED #(.width(1)) u_neq_11 (
        .y(_T_37),
        .a(do_enq),
        .b(do_deq)
    );
    wire _T_39;
    EQ_UNSIGNED #(.width(1)) u_eq_12 (
        .y(_T_39),
        .a(_T_27),
        .b(1'h0)
    );
    wire _T_41;
    EQ_UNSIGNED #(.width(1)) u_eq_13 (
        .y(_T_41),
        .a(_T_28),
        .b(1'h0)
    );
    assign ram__T_43_addr = 1'h0;
    assign ram__T_43_en = 1'h1;
    assign ram__T_43_clk = clock;
    wire [1:0] _T_44;
    assign _T_44 = 2'h0;
    wire [1:0] _T_45;
    assign _T_45 = 2'h0;
    wire _T_46;
    assign _T_46 = 1'h0;
    wire _T_47;
    BITWISEAND #(.width(1)) bitwiseand_14 (
        .y(_T_47),
        .a(_maybe_full__q),
        .b(_T_24)
    );
    wire [1:0] _T_48;
    CAT #(.width_a(1), .width_b(1)) cat_15 (
        .y(_T_48),
        .a(_T_47),
        .b(_T_46)
    );
    assign do_deq = _T_31;
    assign do_enq = _T_29;
    BITS #(.width(2), .high(0), .low(0)) bits_16 (
        .y(io_count),
        .in(_T_48)
    );
    assign io_deq_bits = ram__T_43_data;
    assign io_deq_valid = _T_39;
    assign io_enq_ready = _T_41;
    MUX_UNSIGNED #(.width(1)) u_mux_17 (
        .y(_WTEMP_1),
        .sel(_T_37),
        .a(do_enq),
        .b(_maybe_full__q)
    );
    assign ram__T_34_data = io_enq_bits;
endmodule //Queue
module RAMMEM(read_data, read_clk, read_en, read_addr, write_clk, write_en, write_mask, write_addr, write_data);
    parameter depth = 16;
    parameter addrbits = 4;
    parameter width = 32;
    parameter isSyncRead = 0;
    output [width-1:0] read_data;
    input read_clk;
    input read_en;
    input [addrbits-1:0] read_addr;
    input write_clk;
    input write_en;
    input write_mask;
    input [addrbits-1:0] write_addr;
    input [width-1:0] write_data;
    reg [width-1:0] memcore [0:depth-1];
    wire [addrbits-1:0] final_read_addr;
    generate
        if (isSyncRead) begin: raddr_processor
            reg [addrbits-1:0] read_addr_pipe_0;
            always @(posedge read_clk) begin
                if (read_en) begin
                    read_addr_pipe_0 <= read_addr;
                end
            end
            assign final_read_addr = read_addr_pipe_0;
        end else begin: raddr_processor
            assign final_read_addr = read_addr;
        end
    endgenerate
    assign read_data = memcore[final_read_addr];
    always @(posedge write_clk) begin
        if (write_en & write_mask) begin
            memcore[write_addr] <= write_data;
        end
    end
endmodule // RAMMEM
module DFF_POSCLK(q, d, clk);
    parameter width = 4;
    output reg [width-1:0] q;
    input [width-1:0] d;
    input clk;
    always @(posedge clk) begin
        q <= d;
    end
endmodule // DFF_POSCLK
module MUX_UNSIGNED(y, sel, a, b);
    parameter width = 4;
    output [width-1:0] y;
    input sel;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = sel ? a : b;
endmodule // MUX_UNSIGNED
module EQ_UNSIGNED(y, a, b);
    parameter width = 4;
    output y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a == b;
endmodule // EQ_UNSIGNED
module NEQ_UNSIGNED(y, a, b);
    parameter width = 4;
    output y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a != b;
endmodule // NEQ_UNSIGNED
module CAT(y, a, b);
    parameter width_a = 4;
    parameter width_b = 4;
    output [width_a+width_b-1:0] y;
    input [width_a-1:0] a;
    input [width_b-1:0] b;
    assign y = {a, b};
endmodule // CAT
module BITS(y, in);
    parameter width = 4;
    parameter high = 2;
    parameter low = 0;
    output [high-low:0] y;
    input [width-1:0] in;
    assign y = in[high:low];
endmodule // BITS
module SmallOdds3Filter_1(
    input clock,
    input reset,
    output io_in_ready,
    input io_in_valid,
    input [31:0] io_in_bits,
    input io_out_ready,
    output io_out_valid,
    output [31:0] io_out_bits
);
    wire _T_14;
    BITWISEAND #(.width(1)) bitwiseand_18 (
        .y(_T_14),
        .a(io_out_ready),
        .b(io_in_valid)
    );
    wire [31:0] _T_16;
    wire [31:0] _WTEMP_2;
    PAD_UNSIGNED #(.width(1), .n(32)) u_pad_19 (
        .y(_WTEMP_2),
        .in(1'h1)
    );
    BITWISEAND #(.width(32)) bitwiseand_20 (
        .y(_T_16),
        .a(io_in_bits),
        .b(_WTEMP_2)
    );
    wire _T_18;
    wire [31:0] _WTEMP_3;
    PAD_UNSIGNED #(.width(1), .n(32)) u_pad_21 (
        .y(_WTEMP_3),
        .in(1'h1)
    );
    EQ_UNSIGNED #(.width(32)) u_eq_22 (
        .y(_T_18),
        .a(_T_16),
        .b(_WTEMP_3)
    );
    wire _T_19;
    BITWISEAND #(.width(1)) bitwiseand_23 (
        .y(_T_19),
        .a(_T_14),
        .b(_T_18)
    );
    assign io_in_ready = io_out_ready;
    assign io_out_bits = io_in_bits;
    assign io_out_valid = _T_19;
endmodule //SmallOdds3Filter_1
module ADD_UNSIGNED(y, a, b);
    parameter width = 4;
    output [width:0] y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a + b;
endmodule // ADD_UNSIGNED
module TAIL(y, in);
    parameter width = 4;
    parameter n = 2;
    output [width-n-1:0] y;
    input [width-1:0] in;
    assign y = in[width-n-1:0];
endmodule // TAIL
module GT_UNSIGNED(y, a, b);
    parameter width = 4;
    output y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a > b;
endmodule // GT_UNSIGNED
module BITWISEOR(y, a, b);
    parameter width = 4;
    output [width-1:0] y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a | b;
endmodule // BITWISEOR
