module Queue(
    input clock
);
endmodule //Queue
