module NodeType(
  input   clock
);
endmodule
