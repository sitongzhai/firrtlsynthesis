module DecoupledRealGCDTests4(
    input clock,
    input reset
);
    wire _c__clock;
    wire _c__reset;
    wire _c__io_in_ready;
    wire _c__io_in_valid;
    wire [15:0] _c__io_in_bits_a;
    wire [15:0] _c__io_in_bits_b;
    wire _c__io_out_valid;
    wire [15:0] _c__io_out_bits;
    RealGCD c (
        .clock(_c__clock),
        .reset(_c__reset),
        .io_in_ready(_c__io_in_ready),
        .io_in_valid(_c__io_in_valid),
        .io_in_bits_a(_c__io_in_bits_a),
        .io_in_bits_b(_c__io_in_bits_b),
        .io_out_valid(_c__io_out_valid),
        .io_out_bits(_c__io_out_bits)
    );
    wire [8:0] __T_4__q;
    wire [8:0] __T_4__d;
    DFF_POSCLK #(.width(9)) _T_4 (
        .q(__T_4__q),
        .d(__T_4__d),
        .clk(clock)
    );
    wire [8:0] _WTEMP_4;
    MUX_UNSIGNED #(.width(9)) u_mux_29 (
        .y(__T_4__d),
        .sel(reset),
        .a(9'h0),
        .b(_WTEMP_4)
    );
    wire __T_7__q;
    wire __T_7__d;
    DFF_POSCLK #(.width(1)) _T_7 (
        .q(__T_7__q),
        .d(__T_7__d),
        .clk(clock)
    );
    wire _WTEMP_5;
    MUX_UNSIGNED #(.width(1)) u_mux_30 (
        .y(__T_7__d),
        .sel(reset),
        .a(1'h0),
        .b(_WTEMP_5)
    );
    wire [8:0] __T_10__q;
    wire [8:0] __T_10__d;
    DFF_POSCLK #(.width(9)) _T_10 (
        .q(__T_10__q),
        .d(__T_10__d),
        .clk(clock)
    );
    wire [8:0] _WTEMP_6;
    MUX_UNSIGNED #(.width(9)) u_mux_31 (
        .y(__T_10__d),
        .sel(reset),
        .a(9'h0),
        .b(_WTEMP_6)
    );
    wire __T_13__q;
    wire __T_13__d;
    DFF_POSCLK #(.width(1)) _T_13 (
        .q(__T_13__q),
        .d(__T_13__d),
        .clk(clock)
    );
    wire _WTEMP_7;
    MUX_UNSIGNED #(.width(1)) u_mux_32 (
        .y(__T_13__d),
        .sel(reset),
        .a(1'h0),
        .b(_WTEMP_7)
    );
    wire _T_14;
    BITWISEAND #(.width(1)) bitwiseand_33 (
        .y(_T_14),
        .a(__T_7__q),
        .b(__T_13__q)
    );
    wire _T_16;
    EQ_UNSIGNED #(.width(1)) u_eq_34 (
        .y(_T_16),
        .a(reset),
        .b(1'h0)
    );
    wire _T_18;
    EQ_UNSIGNED #(.width(1)) u_eq_35 (
        .y(_T_18),
        .a(reset),
        .b(1'h0)
    );
    wire [11:0] __T_21__q;
    wire [11:0] __T_21__d;
    DFF_POSCLK #(.width(12)) _T_21 (
        .q(__T_21__q),
        .d(__T_21__d),
        .clk(clock)
    );
    wire [11:0] _WTEMP_8;
    MUX_UNSIGNED #(.width(12)) u_mux_36 (
        .y(__T_21__d),
        .sel(reset),
        .a(12'h0),
        .b(_WTEMP_8)
    );
    wire [12:0] _T_23;
    wire [11:0] _WTEMP_9;
    PAD_UNSIGNED #(.width(1), .n(12)) u_pad_37 (
        .y(_WTEMP_9),
        .in(1'h1)
    );
    ADD_UNSIGNED #(.width(12)) u_add_38 (
        .y(_T_23),
        .a(__T_21__q),
        .b(_WTEMP_9)
    );
    wire [11:0] _T_24;
    TAIL #(.width(13), .n(1)) tail_39 (
        .y(_T_24),
        .in(_T_23)
    );
    wire _T_26;
    GT_UNSIGNED #(.width(12)) u_gt_40 (
        .y(_T_26),
        .a(__T_21__q),
        .b(12'hFA0)
    );
    wire _T_29;
    EQ_UNSIGNED #(.width(1)) u_eq_41 (
        .y(_T_29),
        .a(reset),
        .b(1'h0)
    );
    wire _T_31;
    EQ_UNSIGNED #(.width(1)) u_eq_42 (
        .y(_T_31),
        .a(reset),
        .b(1'h0)
    );
    wire _T_135_0;
    wire _T_135_1;
    wire _T_135_2;
    wire _T_135_3;
    wire _T_135_4;
    wire _T_135_5;
    wire _T_135_6;
    wire _T_135_7;
    wire _T_135_8;
    wire _T_135_9;
    wire _T_135_10;
    wire _T_135_11;
    wire _T_135_12;
    wire _T_135_13;
    wire _T_135_14;
    wire _T_135_15;
    wire _T_135_16;
    wire _T_135_17;
    wire _T_135_18;
    wire _T_135_19;
    wire _T_135_20;
    wire _T_135_21;
    wire _T_135_22;
    wire _T_135_23;
    wire _T_135_24;
    wire _T_135_25;
    wire _T_135_26;
    wire _T_135_27;
    wire _T_135_28;
    wire _T_135_29;
    wire _T_135_30;
    wire _T_135_31;
    wire _T_135_32;
    wire _T_135_33;
    wire _T_135_34;
    wire _T_135_35;
    wire _T_135_36;
    wire _T_135_37;
    wire _T_135_38;
    wire _T_135_39;
    wire _T_135_40;
    wire _T_135_41;
    wire _T_135_42;
    wire _T_135_43;
    wire _T_135_44;
    wire _T_135_45;
    wire _T_135_46;
    wire _T_135_47;
    wire _T_135_48;
    wire _T_135_49;
    wire _T_135_50;
    wire _T_135_51;
    wire _T_135_52;
    wire _T_135_53;
    wire _T_135_54;
    wire _T_135_55;
    wire _T_135_56;
    wire _T_135_57;
    wire _T_135_58;
    wire _T_135_59;
    wire _T_135_60;
    wire _T_135_61;
    wire _T_135_62;
    wire _T_135_63;
    wire _T_135_64;
    wire _T_135_65;
    wire _T_135_66;
    wire _T_135_67;
    wire _T_135_68;
    wire _T_135_69;
    wire _T_135_70;
    wire _T_135_71;
    wire _T_135_72;
    wire _T_135_73;
    wire _T_135_74;
    wire _T_135_75;
    wire _T_135_76;
    wire _T_135_77;
    wire _T_135_78;
    wire _T_135_79;
    wire _T_135_80;
    wire _T_135_81;
    wire _T_135_82;
    wire _T_135_83;
    wire _T_135_84;
    wire _T_135_85;
    wire _T_135_86;
    wire _T_135_87;
    wire _T_135_88;
    wire _T_135_89;
    wire _T_135_90;
    wire _T_135_91;
    wire _T_135_92;
    wire _T_135_93;
    wire _T_135_94;
    wire _T_135_95;
    wire _T_135_96;
    wire _T_135_97;
    wire _T_135_98;
    wire _T_135_99;
    wire _T_135_100;
    wire [6:0] _value__q;
    wire [6:0] _value__d;
    DFF_POSCLK #(.width(7)) value (
        .q(_value__q),
        .d(_value__d),
        .clk(clock)
    );
    wire [6:0] _WTEMP_10;
    MUX_UNSIGNED #(.width(7)) u_mux_43 (
        .y(_value__d),
        .sel(reset),
        .a(7'h0),
        .b(_WTEMP_10)
    );
    wire [3:0] _T_344_0;
    wire [3:0] _T_344_1;
    wire [3:0] _T_344_2;
    wire [3:0] _T_344_3;
    wire [3:0] _T_344_4;
    wire [3:0] _T_344_5;
    wire [3:0] _T_344_6;
    wire [3:0] _T_344_7;
    wire [3:0] _T_344_8;
    wire [3:0] _T_344_9;
    wire [3:0] _T_344_10;
    wire [3:0] _T_344_11;
    wire [3:0] _T_344_12;
    wire [3:0] _T_344_13;
    wire [3:0] _T_344_14;
    wire [3:0] _T_344_15;
    wire [3:0] _T_344_16;
    wire [3:0] _T_344_17;
    wire [3:0] _T_344_18;
    wire [3:0] _T_344_19;
    wire [3:0] _T_344_20;
    wire [3:0] _T_344_21;
    wire [3:0] _T_344_22;
    wire [3:0] _T_344_23;
    wire [3:0] _T_344_24;
    wire [3:0] _T_344_25;
    wire [3:0] _T_344_26;
    wire [3:0] _T_344_27;
    wire [3:0] _T_344_28;
    wire [3:0] _T_344_29;
    wire [3:0] _T_344_30;
    wire [3:0] _T_344_31;
    wire [3:0] _T_344_32;
    wire [3:0] _T_344_33;
    wire [3:0] _T_344_34;
    wire [3:0] _T_344_35;
    wire [3:0] _T_344_36;
    wire [3:0] _T_344_37;
    wire [3:0] _T_344_38;
    wire [3:0] _T_344_39;
    wire [3:0] _T_344_40;
    wire [3:0] _T_344_41;
    wire [3:0] _T_344_42;
    wire [3:0] _T_344_43;
    wire [3:0] _T_344_44;
    wire [3:0] _T_344_45;
    wire [3:0] _T_344_46;
    wire [3:0] _T_344_47;
    wire [3:0] _T_344_48;
    wire [3:0] _T_344_49;
    wire [3:0] _T_344_50;
    wire [3:0] _T_344_51;
    wire [3:0] _T_344_52;
    wire [3:0] _T_344_53;
    wire [3:0] _T_344_54;
    wire [3:0] _T_344_55;
    wire [3:0] _T_344_56;
    wire [3:0] _T_344_57;
    wire [3:0] _T_344_58;
    wire [3:0] _T_344_59;
    wire [3:0] _T_344_60;
    wire [3:0] _T_344_61;
    wire [3:0] _T_344_62;
    wire [3:0] _T_344_63;
    wire [3:0] _T_344_64;
    wire [3:0] _T_344_65;
    wire [3:0] _T_344_66;
    wire [3:0] _T_344_67;
    wire [3:0] _T_344_68;
    wire [3:0] _T_344_69;
    wire [3:0] _T_344_70;
    wire [3:0] _T_344_71;
    wire [3:0] _T_344_72;
    wire [3:0] _T_344_73;
    wire [3:0] _T_344_74;
    wire [3:0] _T_344_75;
    wire [3:0] _T_344_76;
    wire [3:0] _T_344_77;
    wire [3:0] _T_344_78;
    wire [3:0] _T_344_79;
    wire [3:0] _T_344_80;
    wire [3:0] _T_344_81;
    wire [3:0] _T_344_82;
    wire [3:0] _T_344_83;
    wire [3:0] _T_344_84;
    wire [3:0] _T_344_85;
    wire [3:0] _T_344_86;
    wire [3:0] _T_344_87;
    wire [3:0] _T_344_88;
    wire [3:0] _T_344_89;
    wire [3:0] _T_344_90;
    wire [3:0] _T_344_91;
    wire [3:0] _T_344_92;
    wire [3:0] _T_344_93;
    wire [3:0] _T_344_94;
    wire [3:0] _T_344_95;
    wire [3:0] _T_344_96;
    wire [3:0] _T_344_97;
    wire [3:0] _T_344_98;
    wire [3:0] _T_344_99;
    wire [3:0] _T_344_100;
    wire [3:0] _T_551_0;
    wire [3:0] _T_551_1;
    wire [3:0] _T_551_2;
    wire [3:0] _T_551_3;
    wire [3:0] _T_551_4;
    wire [3:0] _T_551_5;
    wire [3:0] _T_551_6;
    wire [3:0] _T_551_7;
    wire [3:0] _T_551_8;
    wire [3:0] _T_551_9;
    wire [3:0] _T_551_10;
    wire [3:0] _T_551_11;
    wire [3:0] _T_551_12;
    wire [3:0] _T_551_13;
    wire [3:0] _T_551_14;
    wire [3:0] _T_551_15;
    wire [3:0] _T_551_16;
    wire [3:0] _T_551_17;
    wire [3:0] _T_551_18;
    wire [3:0] _T_551_19;
    wire [3:0] _T_551_20;
    wire [3:0] _T_551_21;
    wire [3:0] _T_551_22;
    wire [3:0] _T_551_23;
    wire [3:0] _T_551_24;
    wire [3:0] _T_551_25;
    wire [3:0] _T_551_26;
    wire [3:0] _T_551_27;
    wire [3:0] _T_551_28;
    wire [3:0] _T_551_29;
    wire [3:0] _T_551_30;
    wire [3:0] _T_551_31;
    wire [3:0] _T_551_32;
    wire [3:0] _T_551_33;
    wire [3:0] _T_551_34;
    wire [3:0] _T_551_35;
    wire [3:0] _T_551_36;
    wire [3:0] _T_551_37;
    wire [3:0] _T_551_38;
    wire [3:0] _T_551_39;
    wire [3:0] _T_551_40;
    wire [3:0] _T_551_41;
    wire [3:0] _T_551_42;
    wire [3:0] _T_551_43;
    wire [3:0] _T_551_44;
    wire [3:0] _T_551_45;
    wire [3:0] _T_551_46;
    wire [3:0] _T_551_47;
    wire [3:0] _T_551_48;
    wire [3:0] _T_551_49;
    wire [3:0] _T_551_50;
    wire [3:0] _T_551_51;
    wire [3:0] _T_551_52;
    wire [3:0] _T_551_53;
    wire [3:0] _T_551_54;
    wire [3:0] _T_551_55;
    wire [3:0] _T_551_56;
    wire [3:0] _T_551_57;
    wire [3:0] _T_551_58;
    wire [3:0] _T_551_59;
    wire [3:0] _T_551_60;
    wire [3:0] _T_551_61;
    wire [3:0] _T_551_62;
    wire [3:0] _T_551_63;
    wire [3:0] _T_551_64;
    wire [3:0] _T_551_65;
    wire [3:0] _T_551_66;
    wire [3:0] _T_551_67;
    wire [3:0] _T_551_68;
    wire [3:0] _T_551_69;
    wire [3:0] _T_551_70;
    wire [3:0] _T_551_71;
    wire [3:0] _T_551_72;
    wire [3:0] _T_551_73;
    wire [3:0] _T_551_74;
    wire [3:0] _T_551_75;
    wire [3:0] _T_551_76;
    wire [3:0] _T_551_77;
    wire [3:0] _T_551_78;
    wire [3:0] _T_551_79;
    wire [3:0] _T_551_80;
    wire [3:0] _T_551_81;
    wire [3:0] _T_551_82;
    wire [3:0] _T_551_83;
    wire [3:0] _T_551_84;
    wire [3:0] _T_551_85;
    wire [3:0] _T_551_86;
    wire [3:0] _T_551_87;
    wire [3:0] _T_551_88;
    wire [3:0] _T_551_89;
    wire [3:0] _T_551_90;
    wire [3:0] _T_551_91;
    wire [3:0] _T_551_92;
    wire [3:0] _T_551_93;
    wire [3:0] _T_551_94;
    wire [3:0] _T_551_95;
    wire [3:0] _T_551_96;
    wire [3:0] _T_551_97;
    wire [3:0] _T_551_98;
    wire [3:0] _T_551_99;
    wire [3:0] _T_551_100;
    wire _node_8;
    EQ_UNSIGNED #(.width(7)) u_eq_44 (
        .y(_node_8),
        .a(7'd0),
        .b(_value__q)
    );
    wire [3:0] _node_9;
    assign _node_9 = _T_344_0;
    wire _node_10;
    EQ_UNSIGNED #(.width(7)) u_eq_45 (
        .y(_node_10),
        .a(7'd1),
        .b(_value__q)
    );
    wire [3:0] _node_11;
    MUX_UNSIGNED #(.width(4)) u_mux_46 (
        .y(_node_11),
        .sel(_node_10),
        .a(_T_344_1),
        .b(_node_9)
    );
    wire _node_12;
    EQ_UNSIGNED #(.width(7)) u_eq_47 (
        .y(_node_12),
        .a(7'd2),
        .b(_value__q)
    );
    wire [3:0] _node_13;
    MUX_UNSIGNED #(.width(4)) u_mux_48 (
        .y(_node_13),
        .sel(_node_12),
        .a(_T_344_2),
        .b(_node_11)
    );
    wire _node_14;
    EQ_UNSIGNED #(.width(7)) u_eq_49 (
        .y(_node_14),
        .a(7'd3),
        .b(_value__q)
    );
    wire [3:0] _node_15;
    MUX_UNSIGNED #(.width(4)) u_mux_50 (
        .y(_node_15),
        .sel(_node_14),
        .a(_T_344_3),
        .b(_node_13)
    );
    wire _node_16;
    EQ_UNSIGNED #(.width(7)) u_eq_51 (
        .y(_node_16),
        .a(7'd4),
        .b(_value__q)
    );
    wire [3:0] _node_17;
    MUX_UNSIGNED #(.width(4)) u_mux_52 (
        .y(_node_17),
        .sel(_node_16),
        .a(_T_344_4),
        .b(_node_15)
    );
    wire _node_18;
    EQ_UNSIGNED #(.width(7)) u_eq_53 (
        .y(_node_18),
        .a(7'd5),
        .b(_value__q)
    );
    wire [3:0] _node_19;
    MUX_UNSIGNED #(.width(4)) u_mux_54 (
        .y(_node_19),
        .sel(_node_18),
        .a(_T_344_5),
        .b(_node_17)
    );
    wire _node_20;
    EQ_UNSIGNED #(.width(7)) u_eq_55 (
        .y(_node_20),
        .a(7'd6),
        .b(_value__q)
    );
    wire [3:0] _node_21;
    MUX_UNSIGNED #(.width(4)) u_mux_56 (
        .y(_node_21),
        .sel(_node_20),
        .a(_T_344_6),
        .b(_node_19)
    );
    wire _node_22;
    EQ_UNSIGNED #(.width(7)) u_eq_57 (
        .y(_node_22),
        .a(7'd7),
        .b(_value__q)
    );
    wire [3:0] _node_23;
    MUX_UNSIGNED #(.width(4)) u_mux_58 (
        .y(_node_23),
        .sel(_node_22),
        .a(_T_344_7),
        .b(_node_21)
    );
    wire _node_24;
    EQ_UNSIGNED #(.width(7)) u_eq_59 (
        .y(_node_24),
        .a(7'd8),
        .b(_value__q)
    );
    wire [3:0] _node_25;
    MUX_UNSIGNED #(.width(4)) u_mux_60 (
        .y(_node_25),
        .sel(_node_24),
        .a(_T_344_8),
        .b(_node_23)
    );
    wire _node_26;
    EQ_UNSIGNED #(.width(7)) u_eq_61 (
        .y(_node_26),
        .a(7'd9),
        .b(_value__q)
    );
    wire [3:0] _node_27;
    MUX_UNSIGNED #(.width(4)) u_mux_62 (
        .y(_node_27),
        .sel(_node_26),
        .a(_T_344_9),
        .b(_node_25)
    );
    wire _node_28;
    EQ_UNSIGNED #(.width(7)) u_eq_63 (
        .y(_node_28),
        .a(7'd10),
        .b(_value__q)
    );
    wire [3:0] _node_29;
    MUX_UNSIGNED #(.width(4)) u_mux_64 (
        .y(_node_29),
        .sel(_node_28),
        .a(_T_344_10),
        .b(_node_27)
    );
    wire _node_30;
    EQ_UNSIGNED #(.width(7)) u_eq_65 (
        .y(_node_30),
        .a(7'd11),
        .b(_value__q)
    );
    wire [3:0] _node_31;
    MUX_UNSIGNED #(.width(4)) u_mux_66 (
        .y(_node_31),
        .sel(_node_30),
        .a(_T_344_11),
        .b(_node_29)
    );
    wire _node_32;
    EQ_UNSIGNED #(.width(7)) u_eq_67 (
        .y(_node_32),
        .a(7'd12),
        .b(_value__q)
    );
    wire [3:0] _node_33;
    MUX_UNSIGNED #(.width(4)) u_mux_68 (
        .y(_node_33),
        .sel(_node_32),
        .a(_T_344_12),
        .b(_node_31)
    );
    wire _node_34;
    EQ_UNSIGNED #(.width(7)) u_eq_69 (
        .y(_node_34),
        .a(7'd13),
        .b(_value__q)
    );
    wire [3:0] _node_35;
    MUX_UNSIGNED #(.width(4)) u_mux_70 (
        .y(_node_35),
        .sel(_node_34),
        .a(_T_344_13),
        .b(_node_33)
    );
    wire _node_36;
    EQ_UNSIGNED #(.width(7)) u_eq_71 (
        .y(_node_36),
        .a(7'd14),
        .b(_value__q)
    );
    wire [3:0] _node_37;
    MUX_UNSIGNED #(.width(4)) u_mux_72 (
        .y(_node_37),
        .sel(_node_36),
        .a(_T_344_14),
        .b(_node_35)
    );
    wire _node_38;
    EQ_UNSIGNED #(.width(7)) u_eq_73 (
        .y(_node_38),
        .a(7'd15),
        .b(_value__q)
    );
    wire [3:0] _node_39;
    MUX_UNSIGNED #(.width(4)) u_mux_74 (
        .y(_node_39),
        .sel(_node_38),
        .a(_T_344_15),
        .b(_node_37)
    );
    wire _node_40;
    EQ_UNSIGNED #(.width(7)) u_eq_75 (
        .y(_node_40),
        .a(7'd16),
        .b(_value__q)
    );
    wire [3:0] _node_41;
    MUX_UNSIGNED #(.width(4)) u_mux_76 (
        .y(_node_41),
        .sel(_node_40),
        .a(_T_344_16),
        .b(_node_39)
    );
    wire _node_42;
    EQ_UNSIGNED #(.width(7)) u_eq_77 (
        .y(_node_42),
        .a(7'd17),
        .b(_value__q)
    );
    wire [3:0] _node_43;
    MUX_UNSIGNED #(.width(4)) u_mux_78 (
        .y(_node_43),
        .sel(_node_42),
        .a(_T_344_17),
        .b(_node_41)
    );
    wire _node_44;
    EQ_UNSIGNED #(.width(7)) u_eq_79 (
        .y(_node_44),
        .a(7'd18),
        .b(_value__q)
    );
    wire [3:0] _node_45;
    MUX_UNSIGNED #(.width(4)) u_mux_80 (
        .y(_node_45),
        .sel(_node_44),
        .a(_T_344_18),
        .b(_node_43)
    );
    wire _node_46;
    EQ_UNSIGNED #(.width(7)) u_eq_81 (
        .y(_node_46),
        .a(7'd19),
        .b(_value__q)
    );
    wire [3:0] _node_47;
    MUX_UNSIGNED #(.width(4)) u_mux_82 (
        .y(_node_47),
        .sel(_node_46),
        .a(_T_344_19),
        .b(_node_45)
    );
    wire _node_48;
    EQ_UNSIGNED #(.width(7)) u_eq_83 (
        .y(_node_48),
        .a(7'd20),
        .b(_value__q)
    );
    wire [3:0] _node_49;
    MUX_UNSIGNED #(.width(4)) u_mux_84 (
        .y(_node_49),
        .sel(_node_48),
        .a(_T_344_20),
        .b(_node_47)
    );
    wire _node_50;
    EQ_UNSIGNED #(.width(7)) u_eq_85 (
        .y(_node_50),
        .a(7'd21),
        .b(_value__q)
    );
    wire [3:0] _node_51;
    MUX_UNSIGNED #(.width(4)) u_mux_86 (
        .y(_node_51),
        .sel(_node_50),
        .a(_T_344_21),
        .b(_node_49)
    );
    wire _node_52;
    EQ_UNSIGNED #(.width(7)) u_eq_87 (
        .y(_node_52),
        .a(7'd22),
        .b(_value__q)
    );
    wire [3:0] _node_53;
    MUX_UNSIGNED #(.width(4)) u_mux_88 (
        .y(_node_53),
        .sel(_node_52),
        .a(_T_344_22),
        .b(_node_51)
    );
    wire _node_54;
    EQ_UNSIGNED #(.width(7)) u_eq_89 (
        .y(_node_54),
        .a(7'd23),
        .b(_value__q)
    );
    wire [3:0] _node_55;
    MUX_UNSIGNED #(.width(4)) u_mux_90 (
        .y(_node_55),
        .sel(_node_54),
        .a(_T_344_23),
        .b(_node_53)
    );
    wire _node_56;
    EQ_UNSIGNED #(.width(7)) u_eq_91 (
        .y(_node_56),
        .a(7'd24),
        .b(_value__q)
    );
    wire [3:0] _node_57;
    MUX_UNSIGNED #(.width(4)) u_mux_92 (
        .y(_node_57),
        .sel(_node_56),
        .a(_T_344_24),
        .b(_node_55)
    );
    wire _node_58;
    EQ_UNSIGNED #(.width(7)) u_eq_93 (
        .y(_node_58),
        .a(7'd25),
        .b(_value__q)
    );
    wire [3:0] _node_59;
    MUX_UNSIGNED #(.width(4)) u_mux_94 (
        .y(_node_59),
        .sel(_node_58),
        .a(_T_344_25),
        .b(_node_57)
    );
    wire _node_60;
    EQ_UNSIGNED #(.width(7)) u_eq_95 (
        .y(_node_60),
        .a(7'd26),
        .b(_value__q)
    );
    wire [3:0] _node_61;
    MUX_UNSIGNED #(.width(4)) u_mux_96 (
        .y(_node_61),
        .sel(_node_60),
        .a(_T_344_26),
        .b(_node_59)
    );
    wire _node_62;
    EQ_UNSIGNED #(.width(7)) u_eq_97 (
        .y(_node_62),
        .a(7'd27),
        .b(_value__q)
    );
    wire [3:0] _node_63;
    MUX_UNSIGNED #(.width(4)) u_mux_98 (
        .y(_node_63),
        .sel(_node_62),
        .a(_T_344_27),
        .b(_node_61)
    );
    wire _node_64;
    EQ_UNSIGNED #(.width(7)) u_eq_99 (
        .y(_node_64),
        .a(7'd28),
        .b(_value__q)
    );
    wire [3:0] _node_65;
    MUX_UNSIGNED #(.width(4)) u_mux_100 (
        .y(_node_65),
        .sel(_node_64),
        .a(_T_344_28),
        .b(_node_63)
    );
    wire _node_66;
    EQ_UNSIGNED #(.width(7)) u_eq_101 (
        .y(_node_66),
        .a(7'd29),
        .b(_value__q)
    );
    wire [3:0] _node_67;
    MUX_UNSIGNED #(.width(4)) u_mux_102 (
        .y(_node_67),
        .sel(_node_66),
        .a(_T_344_29),
        .b(_node_65)
    );
    wire _node_68;
    EQ_UNSIGNED #(.width(7)) u_eq_103 (
        .y(_node_68),
        .a(7'd30),
        .b(_value__q)
    );
    wire [3:0] _node_69;
    MUX_UNSIGNED #(.width(4)) u_mux_104 (
        .y(_node_69),
        .sel(_node_68),
        .a(_T_344_30),
        .b(_node_67)
    );
    wire _node_70;
    EQ_UNSIGNED #(.width(7)) u_eq_105 (
        .y(_node_70),
        .a(7'd31),
        .b(_value__q)
    );
    wire [3:0] _node_71;
    MUX_UNSIGNED #(.width(4)) u_mux_106 (
        .y(_node_71),
        .sel(_node_70),
        .a(_T_344_31),
        .b(_node_69)
    );
    wire _node_72;
    EQ_UNSIGNED #(.width(7)) u_eq_107 (
        .y(_node_72),
        .a(7'd32),
        .b(_value__q)
    );
    wire [3:0] _node_73;
    MUX_UNSIGNED #(.width(4)) u_mux_108 (
        .y(_node_73),
        .sel(_node_72),
        .a(_T_344_32),
        .b(_node_71)
    );
    wire _node_74;
    EQ_UNSIGNED #(.width(7)) u_eq_109 (
        .y(_node_74),
        .a(7'd33),
        .b(_value__q)
    );
    wire [3:0] _node_75;
    MUX_UNSIGNED #(.width(4)) u_mux_110 (
        .y(_node_75),
        .sel(_node_74),
        .a(_T_344_33),
        .b(_node_73)
    );
    wire _node_76;
    EQ_UNSIGNED #(.width(7)) u_eq_111 (
        .y(_node_76),
        .a(7'd34),
        .b(_value__q)
    );
    wire [3:0] _node_77;
    MUX_UNSIGNED #(.width(4)) u_mux_112 (
        .y(_node_77),
        .sel(_node_76),
        .a(_T_344_34),
        .b(_node_75)
    );
    wire _node_78;
    EQ_UNSIGNED #(.width(7)) u_eq_113 (
        .y(_node_78),
        .a(7'd35),
        .b(_value__q)
    );
    wire [3:0] _node_79;
    MUX_UNSIGNED #(.width(4)) u_mux_114 (
        .y(_node_79),
        .sel(_node_78),
        .a(_T_344_35),
        .b(_node_77)
    );
    wire _node_80;
    EQ_UNSIGNED #(.width(7)) u_eq_115 (
        .y(_node_80),
        .a(7'd36),
        .b(_value__q)
    );
    wire [3:0] _node_81;
    MUX_UNSIGNED #(.width(4)) u_mux_116 (
        .y(_node_81),
        .sel(_node_80),
        .a(_T_344_36),
        .b(_node_79)
    );
    wire _node_82;
    EQ_UNSIGNED #(.width(7)) u_eq_117 (
        .y(_node_82),
        .a(7'd37),
        .b(_value__q)
    );
    wire [3:0] _node_83;
    MUX_UNSIGNED #(.width(4)) u_mux_118 (
        .y(_node_83),
        .sel(_node_82),
        .a(_T_344_37),
        .b(_node_81)
    );
    wire _node_84;
    EQ_UNSIGNED #(.width(7)) u_eq_119 (
        .y(_node_84),
        .a(7'd38),
        .b(_value__q)
    );
    wire [3:0] _node_85;
    MUX_UNSIGNED #(.width(4)) u_mux_120 (
        .y(_node_85),
        .sel(_node_84),
        .a(_T_344_38),
        .b(_node_83)
    );
    wire _node_86;
    EQ_UNSIGNED #(.width(7)) u_eq_121 (
        .y(_node_86),
        .a(7'd39),
        .b(_value__q)
    );
    wire [3:0] _node_87;
    MUX_UNSIGNED #(.width(4)) u_mux_122 (
        .y(_node_87),
        .sel(_node_86),
        .a(_T_344_39),
        .b(_node_85)
    );
    wire _node_88;
    EQ_UNSIGNED #(.width(7)) u_eq_123 (
        .y(_node_88),
        .a(7'd40),
        .b(_value__q)
    );
    wire [3:0] _node_89;
    MUX_UNSIGNED #(.width(4)) u_mux_124 (
        .y(_node_89),
        .sel(_node_88),
        .a(_T_344_40),
        .b(_node_87)
    );
    wire _node_90;
    EQ_UNSIGNED #(.width(7)) u_eq_125 (
        .y(_node_90),
        .a(7'd41),
        .b(_value__q)
    );
    wire [3:0] _node_91;
    MUX_UNSIGNED #(.width(4)) u_mux_126 (
        .y(_node_91),
        .sel(_node_90),
        .a(_T_344_41),
        .b(_node_89)
    );
    wire _node_92;
    EQ_UNSIGNED #(.width(7)) u_eq_127 (
        .y(_node_92),
        .a(7'd42),
        .b(_value__q)
    );
    wire [3:0] _node_93;
    MUX_UNSIGNED #(.width(4)) u_mux_128 (
        .y(_node_93),
        .sel(_node_92),
        .a(_T_344_42),
        .b(_node_91)
    );
    wire _node_94;
    EQ_UNSIGNED #(.width(7)) u_eq_129 (
        .y(_node_94),
        .a(7'd43),
        .b(_value__q)
    );
    wire [3:0] _node_95;
    MUX_UNSIGNED #(.width(4)) u_mux_130 (
        .y(_node_95),
        .sel(_node_94),
        .a(_T_344_43),
        .b(_node_93)
    );
    wire _node_96;
    EQ_UNSIGNED #(.width(7)) u_eq_131 (
        .y(_node_96),
        .a(7'd44),
        .b(_value__q)
    );
    wire [3:0] _node_97;
    MUX_UNSIGNED #(.width(4)) u_mux_132 (
        .y(_node_97),
        .sel(_node_96),
        .a(_T_344_44),
        .b(_node_95)
    );
    wire _node_98;
    EQ_UNSIGNED #(.width(7)) u_eq_133 (
        .y(_node_98),
        .a(7'd45),
        .b(_value__q)
    );
    wire [3:0] _node_99;
    MUX_UNSIGNED #(.width(4)) u_mux_134 (
        .y(_node_99),
        .sel(_node_98),
        .a(_T_344_45),
        .b(_node_97)
    );
    wire _node_100;
    EQ_UNSIGNED #(.width(7)) u_eq_135 (
        .y(_node_100),
        .a(7'd46),
        .b(_value__q)
    );
    wire [3:0] _node_101;
    MUX_UNSIGNED #(.width(4)) u_mux_136 (
        .y(_node_101),
        .sel(_node_100),
        .a(_T_344_46),
        .b(_node_99)
    );
    wire _node_102;
    EQ_UNSIGNED #(.width(7)) u_eq_137 (
        .y(_node_102),
        .a(7'd47),
        .b(_value__q)
    );
    wire [3:0] _node_103;
    MUX_UNSIGNED #(.width(4)) u_mux_138 (
        .y(_node_103),
        .sel(_node_102),
        .a(_T_344_47),
        .b(_node_101)
    );
    wire _node_104;
    EQ_UNSIGNED #(.width(7)) u_eq_139 (
        .y(_node_104),
        .a(7'd48),
        .b(_value__q)
    );
    wire [3:0] _node_105;
    MUX_UNSIGNED #(.width(4)) u_mux_140 (
        .y(_node_105),
        .sel(_node_104),
        .a(_T_344_48),
        .b(_node_103)
    );
    wire _node_106;
    EQ_UNSIGNED #(.width(7)) u_eq_141 (
        .y(_node_106),
        .a(7'd49),
        .b(_value__q)
    );
    wire [3:0] _node_107;
    MUX_UNSIGNED #(.width(4)) u_mux_142 (
        .y(_node_107),
        .sel(_node_106),
        .a(_T_344_49),
        .b(_node_105)
    );
    wire _node_108;
    EQ_UNSIGNED #(.width(7)) u_eq_143 (
        .y(_node_108),
        .a(7'd50),
        .b(_value__q)
    );
    wire [3:0] _node_109;
    MUX_UNSIGNED #(.width(4)) u_mux_144 (
        .y(_node_109),
        .sel(_node_108),
        .a(_T_344_50),
        .b(_node_107)
    );
    wire _node_110;
    EQ_UNSIGNED #(.width(7)) u_eq_145 (
        .y(_node_110),
        .a(7'd51),
        .b(_value__q)
    );
    wire [3:0] _node_111;
    MUX_UNSIGNED #(.width(4)) u_mux_146 (
        .y(_node_111),
        .sel(_node_110),
        .a(_T_344_51),
        .b(_node_109)
    );
    wire _node_112;
    EQ_UNSIGNED #(.width(7)) u_eq_147 (
        .y(_node_112),
        .a(7'd52),
        .b(_value__q)
    );
    wire [3:0] _node_113;
    MUX_UNSIGNED #(.width(4)) u_mux_148 (
        .y(_node_113),
        .sel(_node_112),
        .a(_T_344_52),
        .b(_node_111)
    );
    wire _node_114;
    EQ_UNSIGNED #(.width(7)) u_eq_149 (
        .y(_node_114),
        .a(7'd53),
        .b(_value__q)
    );
    wire [3:0] _node_115;
    MUX_UNSIGNED #(.width(4)) u_mux_150 (
        .y(_node_115),
        .sel(_node_114),
        .a(_T_344_53),
        .b(_node_113)
    );
    wire _node_116;
    EQ_UNSIGNED #(.width(7)) u_eq_151 (
        .y(_node_116),
        .a(7'd54),
        .b(_value__q)
    );
    wire [3:0] _node_117;
    MUX_UNSIGNED #(.width(4)) u_mux_152 (
        .y(_node_117),
        .sel(_node_116),
        .a(_T_344_54),
        .b(_node_115)
    );
    wire _node_118;
    EQ_UNSIGNED #(.width(7)) u_eq_153 (
        .y(_node_118),
        .a(7'd55),
        .b(_value__q)
    );
    wire [3:0] _node_119;
    MUX_UNSIGNED #(.width(4)) u_mux_154 (
        .y(_node_119),
        .sel(_node_118),
        .a(_T_344_55),
        .b(_node_117)
    );
    wire _node_120;
    EQ_UNSIGNED #(.width(7)) u_eq_155 (
        .y(_node_120),
        .a(7'd56),
        .b(_value__q)
    );
    wire [3:0] _node_121;
    MUX_UNSIGNED #(.width(4)) u_mux_156 (
        .y(_node_121),
        .sel(_node_120),
        .a(_T_344_56),
        .b(_node_119)
    );
    wire _node_122;
    EQ_UNSIGNED #(.width(7)) u_eq_157 (
        .y(_node_122),
        .a(7'd57),
        .b(_value__q)
    );
    wire [3:0] _node_123;
    MUX_UNSIGNED #(.width(4)) u_mux_158 (
        .y(_node_123),
        .sel(_node_122),
        .a(_T_344_57),
        .b(_node_121)
    );
    wire _node_124;
    EQ_UNSIGNED #(.width(7)) u_eq_159 (
        .y(_node_124),
        .a(7'd58),
        .b(_value__q)
    );
    wire [3:0] _node_125;
    MUX_UNSIGNED #(.width(4)) u_mux_160 (
        .y(_node_125),
        .sel(_node_124),
        .a(_T_344_58),
        .b(_node_123)
    );
    wire _node_126;
    EQ_UNSIGNED #(.width(7)) u_eq_161 (
        .y(_node_126),
        .a(7'd59),
        .b(_value__q)
    );
    wire [3:0] _node_127;
    MUX_UNSIGNED #(.width(4)) u_mux_162 (
        .y(_node_127),
        .sel(_node_126),
        .a(_T_344_59),
        .b(_node_125)
    );
    wire _node_128;
    EQ_UNSIGNED #(.width(7)) u_eq_163 (
        .y(_node_128),
        .a(7'd60),
        .b(_value__q)
    );
    wire [3:0] _node_129;
    MUX_UNSIGNED #(.width(4)) u_mux_164 (
        .y(_node_129),
        .sel(_node_128),
        .a(_T_344_60),
        .b(_node_127)
    );
    wire _node_130;
    EQ_UNSIGNED #(.width(7)) u_eq_165 (
        .y(_node_130),
        .a(7'd61),
        .b(_value__q)
    );
    wire [3:0] _node_131;
    MUX_UNSIGNED #(.width(4)) u_mux_166 (
        .y(_node_131),
        .sel(_node_130),
        .a(_T_344_61),
        .b(_node_129)
    );
    wire _node_132;
    EQ_UNSIGNED #(.width(7)) u_eq_167 (
        .y(_node_132),
        .a(7'd62),
        .b(_value__q)
    );
    wire [3:0] _node_133;
    MUX_UNSIGNED #(.width(4)) u_mux_168 (
        .y(_node_133),
        .sel(_node_132),
        .a(_T_344_62),
        .b(_node_131)
    );
    wire _node_134;
    EQ_UNSIGNED #(.width(7)) u_eq_169 (
        .y(_node_134),
        .a(7'd63),
        .b(_value__q)
    );
    wire [3:0] _node_135;
    MUX_UNSIGNED #(.width(4)) u_mux_170 (
        .y(_node_135),
        .sel(_node_134),
        .a(_T_344_63),
        .b(_node_133)
    );
    wire _node_136;
    EQ_UNSIGNED #(.width(7)) u_eq_171 (
        .y(_node_136),
        .a(7'd64),
        .b(_value__q)
    );
    wire [3:0] _node_137;
    MUX_UNSIGNED #(.width(4)) u_mux_172 (
        .y(_node_137),
        .sel(_node_136),
        .a(_T_344_64),
        .b(_node_135)
    );
    wire _node_138;
    EQ_UNSIGNED #(.width(7)) u_eq_173 (
        .y(_node_138),
        .a(7'd65),
        .b(_value__q)
    );
    wire [3:0] _node_139;
    MUX_UNSIGNED #(.width(4)) u_mux_174 (
        .y(_node_139),
        .sel(_node_138),
        .a(_T_344_65),
        .b(_node_137)
    );
    wire _node_140;
    EQ_UNSIGNED #(.width(7)) u_eq_175 (
        .y(_node_140),
        .a(7'd66),
        .b(_value__q)
    );
    wire [3:0] _node_141;
    MUX_UNSIGNED #(.width(4)) u_mux_176 (
        .y(_node_141),
        .sel(_node_140),
        .a(_T_344_66),
        .b(_node_139)
    );
    wire _node_142;
    EQ_UNSIGNED #(.width(7)) u_eq_177 (
        .y(_node_142),
        .a(7'd67),
        .b(_value__q)
    );
    wire [3:0] _node_143;
    MUX_UNSIGNED #(.width(4)) u_mux_178 (
        .y(_node_143),
        .sel(_node_142),
        .a(_T_344_67),
        .b(_node_141)
    );
    wire _node_144;
    EQ_UNSIGNED #(.width(7)) u_eq_179 (
        .y(_node_144),
        .a(7'd68),
        .b(_value__q)
    );
    wire [3:0] _node_145;
    MUX_UNSIGNED #(.width(4)) u_mux_180 (
        .y(_node_145),
        .sel(_node_144),
        .a(_T_344_68),
        .b(_node_143)
    );
    wire _node_146;
    EQ_UNSIGNED #(.width(7)) u_eq_181 (
        .y(_node_146),
        .a(7'd69),
        .b(_value__q)
    );
    wire [3:0] _node_147;
    MUX_UNSIGNED #(.width(4)) u_mux_182 (
        .y(_node_147),
        .sel(_node_146),
        .a(_T_344_69),
        .b(_node_145)
    );
    wire _node_148;
    EQ_UNSIGNED #(.width(7)) u_eq_183 (
        .y(_node_148),
        .a(7'd70),
        .b(_value__q)
    );
    wire [3:0] _node_149;
    MUX_UNSIGNED #(.width(4)) u_mux_184 (
        .y(_node_149),
        .sel(_node_148),
        .a(_T_344_70),
        .b(_node_147)
    );
    wire _node_150;
    EQ_UNSIGNED #(.width(7)) u_eq_185 (
        .y(_node_150),
        .a(7'd71),
        .b(_value__q)
    );
    wire [3:0] _node_151;
    MUX_UNSIGNED #(.width(4)) u_mux_186 (
        .y(_node_151),
        .sel(_node_150),
        .a(_T_344_71),
        .b(_node_149)
    );
    wire _node_152;
    EQ_UNSIGNED #(.width(7)) u_eq_187 (
        .y(_node_152),
        .a(7'd72),
        .b(_value__q)
    );
    wire [3:0] _node_153;
    MUX_UNSIGNED #(.width(4)) u_mux_188 (
        .y(_node_153),
        .sel(_node_152),
        .a(_T_344_72),
        .b(_node_151)
    );
    wire _node_154;
    EQ_UNSIGNED #(.width(7)) u_eq_189 (
        .y(_node_154),
        .a(7'd73),
        .b(_value__q)
    );
    wire [3:0] _node_155;
    MUX_UNSIGNED #(.width(4)) u_mux_190 (
        .y(_node_155),
        .sel(_node_154),
        .a(_T_344_73),
        .b(_node_153)
    );
    wire _node_156;
    EQ_UNSIGNED #(.width(7)) u_eq_191 (
        .y(_node_156),
        .a(7'd74),
        .b(_value__q)
    );
    wire [3:0] _node_157;
    MUX_UNSIGNED #(.width(4)) u_mux_192 (
        .y(_node_157),
        .sel(_node_156),
        .a(_T_344_74),
        .b(_node_155)
    );
    wire _node_158;
    EQ_UNSIGNED #(.width(7)) u_eq_193 (
        .y(_node_158),
        .a(7'd75),
        .b(_value__q)
    );
    wire [3:0] _node_159;
    MUX_UNSIGNED #(.width(4)) u_mux_194 (
        .y(_node_159),
        .sel(_node_158),
        .a(_T_344_75),
        .b(_node_157)
    );
    wire _node_160;
    EQ_UNSIGNED #(.width(7)) u_eq_195 (
        .y(_node_160),
        .a(7'd76),
        .b(_value__q)
    );
    wire [3:0] _node_161;
    MUX_UNSIGNED #(.width(4)) u_mux_196 (
        .y(_node_161),
        .sel(_node_160),
        .a(_T_344_76),
        .b(_node_159)
    );
    wire _node_162;
    EQ_UNSIGNED #(.width(7)) u_eq_197 (
        .y(_node_162),
        .a(7'd77),
        .b(_value__q)
    );
    wire [3:0] _node_163;
    MUX_UNSIGNED #(.width(4)) u_mux_198 (
        .y(_node_163),
        .sel(_node_162),
        .a(_T_344_77),
        .b(_node_161)
    );
    wire _node_164;
    EQ_UNSIGNED #(.width(7)) u_eq_199 (
        .y(_node_164),
        .a(7'd78),
        .b(_value__q)
    );
    wire [3:0] _node_165;
    MUX_UNSIGNED #(.width(4)) u_mux_200 (
        .y(_node_165),
        .sel(_node_164),
        .a(_T_344_78),
        .b(_node_163)
    );
    wire _node_166;
    EQ_UNSIGNED #(.width(7)) u_eq_201 (
        .y(_node_166),
        .a(7'd79),
        .b(_value__q)
    );
    wire [3:0] _node_167;
    MUX_UNSIGNED #(.width(4)) u_mux_202 (
        .y(_node_167),
        .sel(_node_166),
        .a(_T_344_79),
        .b(_node_165)
    );
    wire _node_168;
    EQ_UNSIGNED #(.width(7)) u_eq_203 (
        .y(_node_168),
        .a(7'd80),
        .b(_value__q)
    );
    wire [3:0] _node_169;
    MUX_UNSIGNED #(.width(4)) u_mux_204 (
        .y(_node_169),
        .sel(_node_168),
        .a(_T_344_80),
        .b(_node_167)
    );
    wire _node_170;
    EQ_UNSIGNED #(.width(7)) u_eq_205 (
        .y(_node_170),
        .a(7'd81),
        .b(_value__q)
    );
    wire [3:0] _node_171;
    MUX_UNSIGNED #(.width(4)) u_mux_206 (
        .y(_node_171),
        .sel(_node_170),
        .a(_T_344_81),
        .b(_node_169)
    );
    wire _node_172;
    EQ_UNSIGNED #(.width(7)) u_eq_207 (
        .y(_node_172),
        .a(7'd82),
        .b(_value__q)
    );
    wire [3:0] _node_173;
    MUX_UNSIGNED #(.width(4)) u_mux_208 (
        .y(_node_173),
        .sel(_node_172),
        .a(_T_344_82),
        .b(_node_171)
    );
    wire _node_174;
    EQ_UNSIGNED #(.width(7)) u_eq_209 (
        .y(_node_174),
        .a(7'd83),
        .b(_value__q)
    );
    wire [3:0] _node_175;
    MUX_UNSIGNED #(.width(4)) u_mux_210 (
        .y(_node_175),
        .sel(_node_174),
        .a(_T_344_83),
        .b(_node_173)
    );
    wire _node_176;
    EQ_UNSIGNED #(.width(7)) u_eq_211 (
        .y(_node_176),
        .a(7'd84),
        .b(_value__q)
    );
    wire [3:0] _node_177;
    MUX_UNSIGNED #(.width(4)) u_mux_212 (
        .y(_node_177),
        .sel(_node_176),
        .a(_T_344_84),
        .b(_node_175)
    );
    wire _node_178;
    EQ_UNSIGNED #(.width(7)) u_eq_213 (
        .y(_node_178),
        .a(7'd85),
        .b(_value__q)
    );
    wire [3:0] _node_179;
    MUX_UNSIGNED #(.width(4)) u_mux_214 (
        .y(_node_179),
        .sel(_node_178),
        .a(_T_344_85),
        .b(_node_177)
    );
    wire _node_180;
    EQ_UNSIGNED #(.width(7)) u_eq_215 (
        .y(_node_180),
        .a(7'd86),
        .b(_value__q)
    );
    wire [3:0] _node_181;
    MUX_UNSIGNED #(.width(4)) u_mux_216 (
        .y(_node_181),
        .sel(_node_180),
        .a(_T_344_86),
        .b(_node_179)
    );
    wire _node_182;
    EQ_UNSIGNED #(.width(7)) u_eq_217 (
        .y(_node_182),
        .a(7'd87),
        .b(_value__q)
    );
    wire [3:0] _node_183;
    MUX_UNSIGNED #(.width(4)) u_mux_218 (
        .y(_node_183),
        .sel(_node_182),
        .a(_T_344_87),
        .b(_node_181)
    );
    wire _node_184;
    EQ_UNSIGNED #(.width(7)) u_eq_219 (
        .y(_node_184),
        .a(7'd88),
        .b(_value__q)
    );
    wire [3:0] _node_185;
    MUX_UNSIGNED #(.width(4)) u_mux_220 (
        .y(_node_185),
        .sel(_node_184),
        .a(_T_344_88),
        .b(_node_183)
    );
    wire _node_186;
    EQ_UNSIGNED #(.width(7)) u_eq_221 (
        .y(_node_186),
        .a(7'd89),
        .b(_value__q)
    );
    wire [3:0] _node_187;
    MUX_UNSIGNED #(.width(4)) u_mux_222 (
        .y(_node_187),
        .sel(_node_186),
        .a(_T_344_89),
        .b(_node_185)
    );
    wire _node_188;
    EQ_UNSIGNED #(.width(7)) u_eq_223 (
        .y(_node_188),
        .a(7'd90),
        .b(_value__q)
    );
    wire [3:0] _node_189;
    MUX_UNSIGNED #(.width(4)) u_mux_224 (
        .y(_node_189),
        .sel(_node_188),
        .a(_T_344_90),
        .b(_node_187)
    );
    wire _node_190;
    EQ_UNSIGNED #(.width(7)) u_eq_225 (
        .y(_node_190),
        .a(7'd91),
        .b(_value__q)
    );
    wire [3:0] _node_191;
    MUX_UNSIGNED #(.width(4)) u_mux_226 (
        .y(_node_191),
        .sel(_node_190),
        .a(_T_344_91),
        .b(_node_189)
    );
    wire _node_192;
    EQ_UNSIGNED #(.width(7)) u_eq_227 (
        .y(_node_192),
        .a(7'd92),
        .b(_value__q)
    );
    wire [3:0] _node_193;
    MUX_UNSIGNED #(.width(4)) u_mux_228 (
        .y(_node_193),
        .sel(_node_192),
        .a(_T_344_92),
        .b(_node_191)
    );
    wire _node_194;
    EQ_UNSIGNED #(.width(7)) u_eq_229 (
        .y(_node_194),
        .a(7'd93),
        .b(_value__q)
    );
    wire [3:0] _node_195;
    MUX_UNSIGNED #(.width(4)) u_mux_230 (
        .y(_node_195),
        .sel(_node_194),
        .a(_T_344_93),
        .b(_node_193)
    );
    wire _node_196;
    EQ_UNSIGNED #(.width(7)) u_eq_231 (
        .y(_node_196),
        .a(7'd94),
        .b(_value__q)
    );
    wire [3:0] _node_197;
    MUX_UNSIGNED #(.width(4)) u_mux_232 (
        .y(_node_197),
        .sel(_node_196),
        .a(_T_344_94),
        .b(_node_195)
    );
    wire _node_198;
    EQ_UNSIGNED #(.width(7)) u_eq_233 (
        .y(_node_198),
        .a(7'd95),
        .b(_value__q)
    );
    wire [3:0] _node_199;
    MUX_UNSIGNED #(.width(4)) u_mux_234 (
        .y(_node_199),
        .sel(_node_198),
        .a(_T_344_95),
        .b(_node_197)
    );
    wire _node_200;
    EQ_UNSIGNED #(.width(7)) u_eq_235 (
        .y(_node_200),
        .a(7'd96),
        .b(_value__q)
    );
    wire [3:0] _node_201;
    MUX_UNSIGNED #(.width(4)) u_mux_236 (
        .y(_node_201),
        .sel(_node_200),
        .a(_T_344_96),
        .b(_node_199)
    );
    wire _node_202;
    EQ_UNSIGNED #(.width(7)) u_eq_237 (
        .y(_node_202),
        .a(7'd97),
        .b(_value__q)
    );
    wire [3:0] _node_203;
    MUX_UNSIGNED #(.width(4)) u_mux_238 (
        .y(_node_203),
        .sel(_node_202),
        .a(_T_344_97),
        .b(_node_201)
    );
    wire _node_204;
    EQ_UNSIGNED #(.width(7)) u_eq_239 (
        .y(_node_204),
        .a(7'd98),
        .b(_value__q)
    );
    wire [3:0] _node_205;
    MUX_UNSIGNED #(.width(4)) u_mux_240 (
        .y(_node_205),
        .sel(_node_204),
        .a(_T_344_98),
        .b(_node_203)
    );
    wire _node_206;
    EQ_UNSIGNED #(.width(7)) u_eq_241 (
        .y(_node_206),
        .a(7'd99),
        .b(_value__q)
    );
    wire [3:0] _node_207;
    MUX_UNSIGNED #(.width(4)) u_mux_242 (
        .y(_node_207),
        .sel(_node_206),
        .a(_T_344_99),
        .b(_node_205)
    );
    wire _node_208;
    EQ_UNSIGNED #(.width(7)) u_eq_243 (
        .y(_node_208),
        .a(7'd100),
        .b(_value__q)
    );
    wire [3:0] _node_209;
    MUX_UNSIGNED #(.width(4)) u_mux_244 (
        .y(_node_209),
        .sel(_node_208),
        .a(_T_344_100),
        .b(_node_207)
    );
    wire _node_210;
    EQ_UNSIGNED #(.width(7)) u_eq_245 (
        .y(_node_210),
        .a(7'd0),
        .b(_value__q)
    );
    wire [3:0] _node_211;
    assign _node_211 = _T_551_0;
    wire _node_212;
    EQ_UNSIGNED #(.width(7)) u_eq_246 (
        .y(_node_212),
        .a(7'd1),
        .b(_value__q)
    );
    wire [3:0] _node_213;
    MUX_UNSIGNED #(.width(4)) u_mux_247 (
        .y(_node_213),
        .sel(_node_212),
        .a(_T_551_1),
        .b(_node_211)
    );
    wire _node_214;
    EQ_UNSIGNED #(.width(7)) u_eq_248 (
        .y(_node_214),
        .a(7'd2),
        .b(_value__q)
    );
    wire [3:0] _node_215;
    MUX_UNSIGNED #(.width(4)) u_mux_249 (
        .y(_node_215),
        .sel(_node_214),
        .a(_T_551_2),
        .b(_node_213)
    );
    wire _node_216;
    EQ_UNSIGNED #(.width(7)) u_eq_250 (
        .y(_node_216),
        .a(7'd3),
        .b(_value__q)
    );
    wire [3:0] _node_217;
    MUX_UNSIGNED #(.width(4)) u_mux_251 (
        .y(_node_217),
        .sel(_node_216),
        .a(_T_551_3),
        .b(_node_215)
    );
    wire _node_218;
    EQ_UNSIGNED #(.width(7)) u_eq_252 (
        .y(_node_218),
        .a(7'd4),
        .b(_value__q)
    );
    wire [3:0] _node_219;
    MUX_UNSIGNED #(.width(4)) u_mux_253 (
        .y(_node_219),
        .sel(_node_218),
        .a(_T_551_4),
        .b(_node_217)
    );
    wire _node_220;
    EQ_UNSIGNED #(.width(7)) u_eq_254 (
        .y(_node_220),
        .a(7'd5),
        .b(_value__q)
    );
    wire [3:0] _node_221;
    MUX_UNSIGNED #(.width(4)) u_mux_255 (
        .y(_node_221),
        .sel(_node_220),
        .a(_T_551_5),
        .b(_node_219)
    );
    wire _node_222;
    EQ_UNSIGNED #(.width(7)) u_eq_256 (
        .y(_node_222),
        .a(7'd6),
        .b(_value__q)
    );
    wire [3:0] _node_223;
    MUX_UNSIGNED #(.width(4)) u_mux_257 (
        .y(_node_223),
        .sel(_node_222),
        .a(_T_551_6),
        .b(_node_221)
    );
    wire _node_224;
    EQ_UNSIGNED #(.width(7)) u_eq_258 (
        .y(_node_224),
        .a(7'd7),
        .b(_value__q)
    );
    wire [3:0] _node_225;
    MUX_UNSIGNED #(.width(4)) u_mux_259 (
        .y(_node_225),
        .sel(_node_224),
        .a(_T_551_7),
        .b(_node_223)
    );
    wire _node_226;
    EQ_UNSIGNED #(.width(7)) u_eq_260 (
        .y(_node_226),
        .a(7'd8),
        .b(_value__q)
    );
    wire [3:0] _node_227;
    MUX_UNSIGNED #(.width(4)) u_mux_261 (
        .y(_node_227),
        .sel(_node_226),
        .a(_T_551_8),
        .b(_node_225)
    );
    wire _node_228;
    EQ_UNSIGNED #(.width(7)) u_eq_262 (
        .y(_node_228),
        .a(7'd9),
        .b(_value__q)
    );
    wire [3:0] _node_229;
    MUX_UNSIGNED #(.width(4)) u_mux_263 (
        .y(_node_229),
        .sel(_node_228),
        .a(_T_551_9),
        .b(_node_227)
    );
    wire _node_230;
    EQ_UNSIGNED #(.width(7)) u_eq_264 (
        .y(_node_230),
        .a(7'd10),
        .b(_value__q)
    );
    wire [3:0] _node_231;
    MUX_UNSIGNED #(.width(4)) u_mux_265 (
        .y(_node_231),
        .sel(_node_230),
        .a(_T_551_10),
        .b(_node_229)
    );
    wire _node_232;
    EQ_UNSIGNED #(.width(7)) u_eq_266 (
        .y(_node_232),
        .a(7'd11),
        .b(_value__q)
    );
    wire [3:0] _node_233;
    MUX_UNSIGNED #(.width(4)) u_mux_267 (
        .y(_node_233),
        .sel(_node_232),
        .a(_T_551_11),
        .b(_node_231)
    );
    wire _node_234;
    EQ_UNSIGNED #(.width(7)) u_eq_268 (
        .y(_node_234),
        .a(7'd12),
        .b(_value__q)
    );
    wire [3:0] _node_235;
    MUX_UNSIGNED #(.width(4)) u_mux_269 (
        .y(_node_235),
        .sel(_node_234),
        .a(_T_551_12),
        .b(_node_233)
    );
    wire _node_236;
    EQ_UNSIGNED #(.width(7)) u_eq_270 (
        .y(_node_236),
        .a(7'd13),
        .b(_value__q)
    );
    wire [3:0] _node_237;
    MUX_UNSIGNED #(.width(4)) u_mux_271 (
        .y(_node_237),
        .sel(_node_236),
        .a(_T_551_13),
        .b(_node_235)
    );
    wire _node_238;
    EQ_UNSIGNED #(.width(7)) u_eq_272 (
        .y(_node_238),
        .a(7'd14),
        .b(_value__q)
    );
    wire [3:0] _node_239;
    MUX_UNSIGNED #(.width(4)) u_mux_273 (
        .y(_node_239),
        .sel(_node_238),
        .a(_T_551_14),
        .b(_node_237)
    );
    wire _node_240;
    EQ_UNSIGNED #(.width(7)) u_eq_274 (
        .y(_node_240),
        .a(7'd15),
        .b(_value__q)
    );
    wire [3:0] _node_241;
    MUX_UNSIGNED #(.width(4)) u_mux_275 (
        .y(_node_241),
        .sel(_node_240),
        .a(_T_551_15),
        .b(_node_239)
    );
    wire _node_242;
    EQ_UNSIGNED #(.width(7)) u_eq_276 (
        .y(_node_242),
        .a(7'd16),
        .b(_value__q)
    );
    wire [3:0] _node_243;
    MUX_UNSIGNED #(.width(4)) u_mux_277 (
        .y(_node_243),
        .sel(_node_242),
        .a(_T_551_16),
        .b(_node_241)
    );
    wire _node_244;
    EQ_UNSIGNED #(.width(7)) u_eq_278 (
        .y(_node_244),
        .a(7'd17),
        .b(_value__q)
    );
    wire [3:0] _node_245;
    MUX_UNSIGNED #(.width(4)) u_mux_279 (
        .y(_node_245),
        .sel(_node_244),
        .a(_T_551_17),
        .b(_node_243)
    );
    wire _node_246;
    EQ_UNSIGNED #(.width(7)) u_eq_280 (
        .y(_node_246),
        .a(7'd18),
        .b(_value__q)
    );
    wire [3:0] _node_247;
    MUX_UNSIGNED #(.width(4)) u_mux_281 (
        .y(_node_247),
        .sel(_node_246),
        .a(_T_551_18),
        .b(_node_245)
    );
    wire _node_248;
    EQ_UNSIGNED #(.width(7)) u_eq_282 (
        .y(_node_248),
        .a(7'd19),
        .b(_value__q)
    );
    wire [3:0] _node_249;
    MUX_UNSIGNED #(.width(4)) u_mux_283 (
        .y(_node_249),
        .sel(_node_248),
        .a(_T_551_19),
        .b(_node_247)
    );
    wire _node_250;
    EQ_UNSIGNED #(.width(7)) u_eq_284 (
        .y(_node_250),
        .a(7'd20),
        .b(_value__q)
    );
    wire [3:0] _node_251;
    MUX_UNSIGNED #(.width(4)) u_mux_285 (
        .y(_node_251),
        .sel(_node_250),
        .a(_T_551_20),
        .b(_node_249)
    );
    wire _node_252;
    EQ_UNSIGNED #(.width(7)) u_eq_286 (
        .y(_node_252),
        .a(7'd21),
        .b(_value__q)
    );
    wire [3:0] _node_253;
    MUX_UNSIGNED #(.width(4)) u_mux_287 (
        .y(_node_253),
        .sel(_node_252),
        .a(_T_551_21),
        .b(_node_251)
    );
    wire _node_254;
    EQ_UNSIGNED #(.width(7)) u_eq_288 (
        .y(_node_254),
        .a(7'd22),
        .b(_value__q)
    );
    wire [3:0] _node_255;
    MUX_UNSIGNED #(.width(4)) u_mux_289 (
        .y(_node_255),
        .sel(_node_254),
        .a(_T_551_22),
        .b(_node_253)
    );
    wire _node_256;
    EQ_UNSIGNED #(.width(7)) u_eq_290 (
        .y(_node_256),
        .a(7'd23),
        .b(_value__q)
    );
    wire [3:0] _node_257;
    MUX_UNSIGNED #(.width(4)) u_mux_291 (
        .y(_node_257),
        .sel(_node_256),
        .a(_T_551_23),
        .b(_node_255)
    );
    wire _node_258;
    EQ_UNSIGNED #(.width(7)) u_eq_292 (
        .y(_node_258),
        .a(7'd24),
        .b(_value__q)
    );
    wire [3:0] _node_259;
    MUX_UNSIGNED #(.width(4)) u_mux_293 (
        .y(_node_259),
        .sel(_node_258),
        .a(_T_551_24),
        .b(_node_257)
    );
    wire _node_260;
    EQ_UNSIGNED #(.width(7)) u_eq_294 (
        .y(_node_260),
        .a(7'd25),
        .b(_value__q)
    );
    wire [3:0] _node_261;
    MUX_UNSIGNED #(.width(4)) u_mux_295 (
        .y(_node_261),
        .sel(_node_260),
        .a(_T_551_25),
        .b(_node_259)
    );
    wire _node_262;
    EQ_UNSIGNED #(.width(7)) u_eq_296 (
        .y(_node_262),
        .a(7'd26),
        .b(_value__q)
    );
    wire [3:0] _node_263;
    MUX_UNSIGNED #(.width(4)) u_mux_297 (
        .y(_node_263),
        .sel(_node_262),
        .a(_T_551_26),
        .b(_node_261)
    );
    wire _node_264;
    EQ_UNSIGNED #(.width(7)) u_eq_298 (
        .y(_node_264),
        .a(7'd27),
        .b(_value__q)
    );
    wire [3:0] _node_265;
    MUX_UNSIGNED #(.width(4)) u_mux_299 (
        .y(_node_265),
        .sel(_node_264),
        .a(_T_551_27),
        .b(_node_263)
    );
    wire _node_266;
    EQ_UNSIGNED #(.width(7)) u_eq_300 (
        .y(_node_266),
        .a(7'd28),
        .b(_value__q)
    );
    wire [3:0] _node_267;
    MUX_UNSIGNED #(.width(4)) u_mux_301 (
        .y(_node_267),
        .sel(_node_266),
        .a(_T_551_28),
        .b(_node_265)
    );
    wire _node_268;
    EQ_UNSIGNED #(.width(7)) u_eq_302 (
        .y(_node_268),
        .a(7'd29),
        .b(_value__q)
    );
    wire [3:0] _node_269;
    MUX_UNSIGNED #(.width(4)) u_mux_303 (
        .y(_node_269),
        .sel(_node_268),
        .a(_T_551_29),
        .b(_node_267)
    );
    wire _node_270;
    EQ_UNSIGNED #(.width(7)) u_eq_304 (
        .y(_node_270),
        .a(7'd30),
        .b(_value__q)
    );
    wire [3:0] _node_271;
    MUX_UNSIGNED #(.width(4)) u_mux_305 (
        .y(_node_271),
        .sel(_node_270),
        .a(_T_551_30),
        .b(_node_269)
    );
    wire _node_272;
    EQ_UNSIGNED #(.width(7)) u_eq_306 (
        .y(_node_272),
        .a(7'd31),
        .b(_value__q)
    );
    wire [3:0] _node_273;
    MUX_UNSIGNED #(.width(4)) u_mux_307 (
        .y(_node_273),
        .sel(_node_272),
        .a(_T_551_31),
        .b(_node_271)
    );
    wire _node_274;
    EQ_UNSIGNED #(.width(7)) u_eq_308 (
        .y(_node_274),
        .a(7'd32),
        .b(_value__q)
    );
    wire [3:0] _node_275;
    MUX_UNSIGNED #(.width(4)) u_mux_309 (
        .y(_node_275),
        .sel(_node_274),
        .a(_T_551_32),
        .b(_node_273)
    );
    wire _node_276;
    EQ_UNSIGNED #(.width(7)) u_eq_310 (
        .y(_node_276),
        .a(7'd33),
        .b(_value__q)
    );
    wire [3:0] _node_277;
    MUX_UNSIGNED #(.width(4)) u_mux_311 (
        .y(_node_277),
        .sel(_node_276),
        .a(_T_551_33),
        .b(_node_275)
    );
    wire _node_278;
    EQ_UNSIGNED #(.width(7)) u_eq_312 (
        .y(_node_278),
        .a(7'd34),
        .b(_value__q)
    );
    wire [3:0] _node_279;
    MUX_UNSIGNED #(.width(4)) u_mux_313 (
        .y(_node_279),
        .sel(_node_278),
        .a(_T_551_34),
        .b(_node_277)
    );
    wire _node_280;
    EQ_UNSIGNED #(.width(7)) u_eq_314 (
        .y(_node_280),
        .a(7'd35),
        .b(_value__q)
    );
    wire [3:0] _node_281;
    MUX_UNSIGNED #(.width(4)) u_mux_315 (
        .y(_node_281),
        .sel(_node_280),
        .a(_T_551_35),
        .b(_node_279)
    );
    wire _node_282;
    EQ_UNSIGNED #(.width(7)) u_eq_316 (
        .y(_node_282),
        .a(7'd36),
        .b(_value__q)
    );
    wire [3:0] _node_283;
    MUX_UNSIGNED #(.width(4)) u_mux_317 (
        .y(_node_283),
        .sel(_node_282),
        .a(_T_551_36),
        .b(_node_281)
    );
    wire _node_284;
    EQ_UNSIGNED #(.width(7)) u_eq_318 (
        .y(_node_284),
        .a(7'd37),
        .b(_value__q)
    );
    wire [3:0] _node_285;
    MUX_UNSIGNED #(.width(4)) u_mux_319 (
        .y(_node_285),
        .sel(_node_284),
        .a(_T_551_37),
        .b(_node_283)
    );
    wire _node_286;
    EQ_UNSIGNED #(.width(7)) u_eq_320 (
        .y(_node_286),
        .a(7'd38),
        .b(_value__q)
    );
    wire [3:0] _node_287;
    MUX_UNSIGNED #(.width(4)) u_mux_321 (
        .y(_node_287),
        .sel(_node_286),
        .a(_T_551_38),
        .b(_node_285)
    );
    wire _node_288;
    EQ_UNSIGNED #(.width(7)) u_eq_322 (
        .y(_node_288),
        .a(7'd39),
        .b(_value__q)
    );
    wire [3:0] _node_289;
    MUX_UNSIGNED #(.width(4)) u_mux_323 (
        .y(_node_289),
        .sel(_node_288),
        .a(_T_551_39),
        .b(_node_287)
    );
    wire _node_290;
    EQ_UNSIGNED #(.width(7)) u_eq_324 (
        .y(_node_290),
        .a(7'd40),
        .b(_value__q)
    );
    wire [3:0] _node_291;
    MUX_UNSIGNED #(.width(4)) u_mux_325 (
        .y(_node_291),
        .sel(_node_290),
        .a(_T_551_40),
        .b(_node_289)
    );
    wire _node_292;
    EQ_UNSIGNED #(.width(7)) u_eq_326 (
        .y(_node_292),
        .a(7'd41),
        .b(_value__q)
    );
    wire [3:0] _node_293;
    MUX_UNSIGNED #(.width(4)) u_mux_327 (
        .y(_node_293),
        .sel(_node_292),
        .a(_T_551_41),
        .b(_node_291)
    );
    wire _node_294;
    EQ_UNSIGNED #(.width(7)) u_eq_328 (
        .y(_node_294),
        .a(7'd42),
        .b(_value__q)
    );
    wire [3:0] _node_295;
    MUX_UNSIGNED #(.width(4)) u_mux_329 (
        .y(_node_295),
        .sel(_node_294),
        .a(_T_551_42),
        .b(_node_293)
    );
    wire _node_296;
    EQ_UNSIGNED #(.width(7)) u_eq_330 (
        .y(_node_296),
        .a(7'd43),
        .b(_value__q)
    );
    wire [3:0] _node_297;
    MUX_UNSIGNED #(.width(4)) u_mux_331 (
        .y(_node_297),
        .sel(_node_296),
        .a(_T_551_43),
        .b(_node_295)
    );
    wire _node_298;
    EQ_UNSIGNED #(.width(7)) u_eq_332 (
        .y(_node_298),
        .a(7'd44),
        .b(_value__q)
    );
    wire [3:0] _node_299;
    MUX_UNSIGNED #(.width(4)) u_mux_333 (
        .y(_node_299),
        .sel(_node_298),
        .a(_T_551_44),
        .b(_node_297)
    );
    wire _node_300;
    EQ_UNSIGNED #(.width(7)) u_eq_334 (
        .y(_node_300),
        .a(7'd45),
        .b(_value__q)
    );
    wire [3:0] _node_301;
    MUX_UNSIGNED #(.width(4)) u_mux_335 (
        .y(_node_301),
        .sel(_node_300),
        .a(_T_551_45),
        .b(_node_299)
    );
    wire _node_302;
    EQ_UNSIGNED #(.width(7)) u_eq_336 (
        .y(_node_302),
        .a(7'd46),
        .b(_value__q)
    );
    wire [3:0] _node_303;
    MUX_UNSIGNED #(.width(4)) u_mux_337 (
        .y(_node_303),
        .sel(_node_302),
        .a(_T_551_46),
        .b(_node_301)
    );
    wire _node_304;
    EQ_UNSIGNED #(.width(7)) u_eq_338 (
        .y(_node_304),
        .a(7'd47),
        .b(_value__q)
    );
    wire [3:0] _node_305;
    MUX_UNSIGNED #(.width(4)) u_mux_339 (
        .y(_node_305),
        .sel(_node_304),
        .a(_T_551_47),
        .b(_node_303)
    );
    wire _node_306;
    EQ_UNSIGNED #(.width(7)) u_eq_340 (
        .y(_node_306),
        .a(7'd48),
        .b(_value__q)
    );
    wire [3:0] _node_307;
    MUX_UNSIGNED #(.width(4)) u_mux_341 (
        .y(_node_307),
        .sel(_node_306),
        .a(_T_551_48),
        .b(_node_305)
    );
    wire _node_308;
    EQ_UNSIGNED #(.width(7)) u_eq_342 (
        .y(_node_308),
        .a(7'd49),
        .b(_value__q)
    );
    wire [3:0] _node_309;
    MUX_UNSIGNED #(.width(4)) u_mux_343 (
        .y(_node_309),
        .sel(_node_308),
        .a(_T_551_49),
        .b(_node_307)
    );
    wire _node_310;
    EQ_UNSIGNED #(.width(7)) u_eq_344 (
        .y(_node_310),
        .a(7'd50),
        .b(_value__q)
    );
    wire [3:0] _node_311;
    MUX_UNSIGNED #(.width(4)) u_mux_345 (
        .y(_node_311),
        .sel(_node_310),
        .a(_T_551_50),
        .b(_node_309)
    );
    wire _node_312;
    EQ_UNSIGNED #(.width(7)) u_eq_346 (
        .y(_node_312),
        .a(7'd51),
        .b(_value__q)
    );
    wire [3:0] _node_313;
    MUX_UNSIGNED #(.width(4)) u_mux_347 (
        .y(_node_313),
        .sel(_node_312),
        .a(_T_551_51),
        .b(_node_311)
    );
    wire _node_314;
    EQ_UNSIGNED #(.width(7)) u_eq_348 (
        .y(_node_314),
        .a(7'd52),
        .b(_value__q)
    );
    wire [3:0] _node_315;
    MUX_UNSIGNED #(.width(4)) u_mux_349 (
        .y(_node_315),
        .sel(_node_314),
        .a(_T_551_52),
        .b(_node_313)
    );
    wire _node_316;
    EQ_UNSIGNED #(.width(7)) u_eq_350 (
        .y(_node_316),
        .a(7'd53),
        .b(_value__q)
    );
    wire [3:0] _node_317;
    MUX_UNSIGNED #(.width(4)) u_mux_351 (
        .y(_node_317),
        .sel(_node_316),
        .a(_T_551_53),
        .b(_node_315)
    );
    wire _node_318;
    EQ_UNSIGNED #(.width(7)) u_eq_352 (
        .y(_node_318),
        .a(7'd54),
        .b(_value__q)
    );
    wire [3:0] _node_319;
    MUX_UNSIGNED #(.width(4)) u_mux_353 (
        .y(_node_319),
        .sel(_node_318),
        .a(_T_551_54),
        .b(_node_317)
    );
    wire _node_320;
    EQ_UNSIGNED #(.width(7)) u_eq_354 (
        .y(_node_320),
        .a(7'd55),
        .b(_value__q)
    );
    wire [3:0] _node_321;
    MUX_UNSIGNED #(.width(4)) u_mux_355 (
        .y(_node_321),
        .sel(_node_320),
        .a(_T_551_55),
        .b(_node_319)
    );
    wire _node_322;
    EQ_UNSIGNED #(.width(7)) u_eq_356 (
        .y(_node_322),
        .a(7'd56),
        .b(_value__q)
    );
    wire [3:0] _node_323;
    MUX_UNSIGNED #(.width(4)) u_mux_357 (
        .y(_node_323),
        .sel(_node_322),
        .a(_T_551_56),
        .b(_node_321)
    );
    wire _node_324;
    EQ_UNSIGNED #(.width(7)) u_eq_358 (
        .y(_node_324),
        .a(7'd57),
        .b(_value__q)
    );
    wire [3:0] _node_325;
    MUX_UNSIGNED #(.width(4)) u_mux_359 (
        .y(_node_325),
        .sel(_node_324),
        .a(_T_551_57),
        .b(_node_323)
    );
    wire _node_326;
    EQ_UNSIGNED #(.width(7)) u_eq_360 (
        .y(_node_326),
        .a(7'd58),
        .b(_value__q)
    );
    wire [3:0] _node_327;
    MUX_UNSIGNED #(.width(4)) u_mux_361 (
        .y(_node_327),
        .sel(_node_326),
        .a(_T_551_58),
        .b(_node_325)
    );
    wire _node_328;
    EQ_UNSIGNED #(.width(7)) u_eq_362 (
        .y(_node_328),
        .a(7'd59),
        .b(_value__q)
    );
    wire [3:0] _node_329;
    MUX_UNSIGNED #(.width(4)) u_mux_363 (
        .y(_node_329),
        .sel(_node_328),
        .a(_T_551_59),
        .b(_node_327)
    );
    wire _node_330;
    EQ_UNSIGNED #(.width(7)) u_eq_364 (
        .y(_node_330),
        .a(7'd60),
        .b(_value__q)
    );
    wire [3:0] _node_331;
    MUX_UNSIGNED #(.width(4)) u_mux_365 (
        .y(_node_331),
        .sel(_node_330),
        .a(_T_551_60),
        .b(_node_329)
    );
    wire _node_332;
    EQ_UNSIGNED #(.width(7)) u_eq_366 (
        .y(_node_332),
        .a(7'd61),
        .b(_value__q)
    );
    wire [3:0] _node_333;
    MUX_UNSIGNED #(.width(4)) u_mux_367 (
        .y(_node_333),
        .sel(_node_332),
        .a(_T_551_61),
        .b(_node_331)
    );
    wire _node_334;
    EQ_UNSIGNED #(.width(7)) u_eq_368 (
        .y(_node_334),
        .a(7'd62),
        .b(_value__q)
    );
    wire [3:0] _node_335;
    MUX_UNSIGNED #(.width(4)) u_mux_369 (
        .y(_node_335),
        .sel(_node_334),
        .a(_T_551_62),
        .b(_node_333)
    );
    wire _node_336;
    EQ_UNSIGNED #(.width(7)) u_eq_370 (
        .y(_node_336),
        .a(7'd63),
        .b(_value__q)
    );
    wire [3:0] _node_337;
    MUX_UNSIGNED #(.width(4)) u_mux_371 (
        .y(_node_337),
        .sel(_node_336),
        .a(_T_551_63),
        .b(_node_335)
    );
    wire _node_338;
    EQ_UNSIGNED #(.width(7)) u_eq_372 (
        .y(_node_338),
        .a(7'd64),
        .b(_value__q)
    );
    wire [3:0] _node_339;
    MUX_UNSIGNED #(.width(4)) u_mux_373 (
        .y(_node_339),
        .sel(_node_338),
        .a(_T_551_64),
        .b(_node_337)
    );
    wire _node_340;
    EQ_UNSIGNED #(.width(7)) u_eq_374 (
        .y(_node_340),
        .a(7'd65),
        .b(_value__q)
    );
    wire [3:0] _node_341;
    MUX_UNSIGNED #(.width(4)) u_mux_375 (
        .y(_node_341),
        .sel(_node_340),
        .a(_T_551_65),
        .b(_node_339)
    );
    wire _node_342;
    EQ_UNSIGNED #(.width(7)) u_eq_376 (
        .y(_node_342),
        .a(7'd66),
        .b(_value__q)
    );
    wire [3:0] _node_343;
    MUX_UNSIGNED #(.width(4)) u_mux_377 (
        .y(_node_343),
        .sel(_node_342),
        .a(_T_551_66),
        .b(_node_341)
    );
    wire _node_344;
    EQ_UNSIGNED #(.width(7)) u_eq_378 (
        .y(_node_344),
        .a(7'd67),
        .b(_value__q)
    );
    wire [3:0] _node_345;
    MUX_UNSIGNED #(.width(4)) u_mux_379 (
        .y(_node_345),
        .sel(_node_344),
        .a(_T_551_67),
        .b(_node_343)
    );
    wire _node_346;
    EQ_UNSIGNED #(.width(7)) u_eq_380 (
        .y(_node_346),
        .a(7'd68),
        .b(_value__q)
    );
    wire [3:0] _node_347;
    MUX_UNSIGNED #(.width(4)) u_mux_381 (
        .y(_node_347),
        .sel(_node_346),
        .a(_T_551_68),
        .b(_node_345)
    );
    wire _node_348;
    EQ_UNSIGNED #(.width(7)) u_eq_382 (
        .y(_node_348),
        .a(7'd69),
        .b(_value__q)
    );
    wire [3:0] _node_349;
    MUX_UNSIGNED #(.width(4)) u_mux_383 (
        .y(_node_349),
        .sel(_node_348),
        .a(_T_551_69),
        .b(_node_347)
    );
    wire _node_350;
    EQ_UNSIGNED #(.width(7)) u_eq_384 (
        .y(_node_350),
        .a(7'd70),
        .b(_value__q)
    );
    wire [3:0] _node_351;
    MUX_UNSIGNED #(.width(4)) u_mux_385 (
        .y(_node_351),
        .sel(_node_350),
        .a(_T_551_70),
        .b(_node_349)
    );
    wire _node_352;
    EQ_UNSIGNED #(.width(7)) u_eq_386 (
        .y(_node_352),
        .a(7'd71),
        .b(_value__q)
    );
    wire [3:0] _node_353;
    MUX_UNSIGNED #(.width(4)) u_mux_387 (
        .y(_node_353),
        .sel(_node_352),
        .a(_T_551_71),
        .b(_node_351)
    );
    wire _node_354;
    EQ_UNSIGNED #(.width(7)) u_eq_388 (
        .y(_node_354),
        .a(7'd72),
        .b(_value__q)
    );
    wire [3:0] _node_355;
    MUX_UNSIGNED #(.width(4)) u_mux_389 (
        .y(_node_355),
        .sel(_node_354),
        .a(_T_551_72),
        .b(_node_353)
    );
    wire _node_356;
    EQ_UNSIGNED #(.width(7)) u_eq_390 (
        .y(_node_356),
        .a(7'd73),
        .b(_value__q)
    );
    wire [3:0] _node_357;
    MUX_UNSIGNED #(.width(4)) u_mux_391 (
        .y(_node_357),
        .sel(_node_356),
        .a(_T_551_73),
        .b(_node_355)
    );
    wire _node_358;
    EQ_UNSIGNED #(.width(7)) u_eq_392 (
        .y(_node_358),
        .a(7'd74),
        .b(_value__q)
    );
    wire [3:0] _node_359;
    MUX_UNSIGNED #(.width(4)) u_mux_393 (
        .y(_node_359),
        .sel(_node_358),
        .a(_T_551_74),
        .b(_node_357)
    );
    wire _node_360;
    EQ_UNSIGNED #(.width(7)) u_eq_394 (
        .y(_node_360),
        .a(7'd75),
        .b(_value__q)
    );
    wire [3:0] _node_361;
    MUX_UNSIGNED #(.width(4)) u_mux_395 (
        .y(_node_361),
        .sel(_node_360),
        .a(_T_551_75),
        .b(_node_359)
    );
    wire _node_362;
    EQ_UNSIGNED #(.width(7)) u_eq_396 (
        .y(_node_362),
        .a(7'd76),
        .b(_value__q)
    );
    wire [3:0] _node_363;
    MUX_UNSIGNED #(.width(4)) u_mux_397 (
        .y(_node_363),
        .sel(_node_362),
        .a(_T_551_76),
        .b(_node_361)
    );
    wire _node_364;
    EQ_UNSIGNED #(.width(7)) u_eq_398 (
        .y(_node_364),
        .a(7'd77),
        .b(_value__q)
    );
    wire [3:0] _node_365;
    MUX_UNSIGNED #(.width(4)) u_mux_399 (
        .y(_node_365),
        .sel(_node_364),
        .a(_T_551_77),
        .b(_node_363)
    );
    wire _node_366;
    EQ_UNSIGNED #(.width(7)) u_eq_400 (
        .y(_node_366),
        .a(7'd78),
        .b(_value__q)
    );
    wire [3:0] _node_367;
    MUX_UNSIGNED #(.width(4)) u_mux_401 (
        .y(_node_367),
        .sel(_node_366),
        .a(_T_551_78),
        .b(_node_365)
    );
    wire _node_368;
    EQ_UNSIGNED #(.width(7)) u_eq_402 (
        .y(_node_368),
        .a(7'd79),
        .b(_value__q)
    );
    wire [3:0] _node_369;
    MUX_UNSIGNED #(.width(4)) u_mux_403 (
        .y(_node_369),
        .sel(_node_368),
        .a(_T_551_79),
        .b(_node_367)
    );
    wire _node_370;
    EQ_UNSIGNED #(.width(7)) u_eq_404 (
        .y(_node_370),
        .a(7'd80),
        .b(_value__q)
    );
    wire [3:0] _node_371;
    MUX_UNSIGNED #(.width(4)) u_mux_405 (
        .y(_node_371),
        .sel(_node_370),
        .a(_T_551_80),
        .b(_node_369)
    );
    wire _node_372;
    EQ_UNSIGNED #(.width(7)) u_eq_406 (
        .y(_node_372),
        .a(7'd81),
        .b(_value__q)
    );
    wire [3:0] _node_373;
    MUX_UNSIGNED #(.width(4)) u_mux_407 (
        .y(_node_373),
        .sel(_node_372),
        .a(_T_551_81),
        .b(_node_371)
    );
    wire _node_374;
    EQ_UNSIGNED #(.width(7)) u_eq_408 (
        .y(_node_374),
        .a(7'd82),
        .b(_value__q)
    );
    wire [3:0] _node_375;
    MUX_UNSIGNED #(.width(4)) u_mux_409 (
        .y(_node_375),
        .sel(_node_374),
        .a(_T_551_82),
        .b(_node_373)
    );
    wire _node_376;
    EQ_UNSIGNED #(.width(7)) u_eq_410 (
        .y(_node_376),
        .a(7'd83),
        .b(_value__q)
    );
    wire [3:0] _node_377;
    MUX_UNSIGNED #(.width(4)) u_mux_411 (
        .y(_node_377),
        .sel(_node_376),
        .a(_T_551_83),
        .b(_node_375)
    );
    wire _node_378;
    EQ_UNSIGNED #(.width(7)) u_eq_412 (
        .y(_node_378),
        .a(7'd84),
        .b(_value__q)
    );
    wire [3:0] _node_379;
    MUX_UNSIGNED #(.width(4)) u_mux_413 (
        .y(_node_379),
        .sel(_node_378),
        .a(_T_551_84),
        .b(_node_377)
    );
    wire _node_380;
    EQ_UNSIGNED #(.width(7)) u_eq_414 (
        .y(_node_380),
        .a(7'd85),
        .b(_value__q)
    );
    wire [3:0] _node_381;
    MUX_UNSIGNED #(.width(4)) u_mux_415 (
        .y(_node_381),
        .sel(_node_380),
        .a(_T_551_85),
        .b(_node_379)
    );
    wire _node_382;
    EQ_UNSIGNED #(.width(7)) u_eq_416 (
        .y(_node_382),
        .a(7'd86),
        .b(_value__q)
    );
    wire [3:0] _node_383;
    MUX_UNSIGNED #(.width(4)) u_mux_417 (
        .y(_node_383),
        .sel(_node_382),
        .a(_T_551_86),
        .b(_node_381)
    );
    wire _node_384;
    EQ_UNSIGNED #(.width(7)) u_eq_418 (
        .y(_node_384),
        .a(7'd87),
        .b(_value__q)
    );
    wire [3:0] _node_385;
    MUX_UNSIGNED #(.width(4)) u_mux_419 (
        .y(_node_385),
        .sel(_node_384),
        .a(_T_551_87),
        .b(_node_383)
    );
    wire _node_386;
    EQ_UNSIGNED #(.width(7)) u_eq_420 (
        .y(_node_386),
        .a(7'd88),
        .b(_value__q)
    );
    wire [3:0] _node_387;
    MUX_UNSIGNED #(.width(4)) u_mux_421 (
        .y(_node_387),
        .sel(_node_386),
        .a(_T_551_88),
        .b(_node_385)
    );
    wire _node_388;
    EQ_UNSIGNED #(.width(7)) u_eq_422 (
        .y(_node_388),
        .a(7'd89),
        .b(_value__q)
    );
    wire [3:0] _node_389;
    MUX_UNSIGNED #(.width(4)) u_mux_423 (
        .y(_node_389),
        .sel(_node_388),
        .a(_T_551_89),
        .b(_node_387)
    );
    wire _node_390;
    EQ_UNSIGNED #(.width(7)) u_eq_424 (
        .y(_node_390),
        .a(7'd90),
        .b(_value__q)
    );
    wire [3:0] _node_391;
    MUX_UNSIGNED #(.width(4)) u_mux_425 (
        .y(_node_391),
        .sel(_node_390),
        .a(_T_551_90),
        .b(_node_389)
    );
    wire _node_392;
    EQ_UNSIGNED #(.width(7)) u_eq_426 (
        .y(_node_392),
        .a(7'd91),
        .b(_value__q)
    );
    wire [3:0] _node_393;
    MUX_UNSIGNED #(.width(4)) u_mux_427 (
        .y(_node_393),
        .sel(_node_392),
        .a(_T_551_91),
        .b(_node_391)
    );
    wire _node_394;
    EQ_UNSIGNED #(.width(7)) u_eq_428 (
        .y(_node_394),
        .a(7'd92),
        .b(_value__q)
    );
    wire [3:0] _node_395;
    MUX_UNSIGNED #(.width(4)) u_mux_429 (
        .y(_node_395),
        .sel(_node_394),
        .a(_T_551_92),
        .b(_node_393)
    );
    wire _node_396;
    EQ_UNSIGNED #(.width(7)) u_eq_430 (
        .y(_node_396),
        .a(7'd93),
        .b(_value__q)
    );
    wire [3:0] _node_397;
    MUX_UNSIGNED #(.width(4)) u_mux_431 (
        .y(_node_397),
        .sel(_node_396),
        .a(_T_551_93),
        .b(_node_395)
    );
    wire _node_398;
    EQ_UNSIGNED #(.width(7)) u_eq_432 (
        .y(_node_398),
        .a(7'd94),
        .b(_value__q)
    );
    wire [3:0] _node_399;
    MUX_UNSIGNED #(.width(4)) u_mux_433 (
        .y(_node_399),
        .sel(_node_398),
        .a(_T_551_94),
        .b(_node_397)
    );
    wire _node_400;
    EQ_UNSIGNED #(.width(7)) u_eq_434 (
        .y(_node_400),
        .a(7'd95),
        .b(_value__q)
    );
    wire [3:0] _node_401;
    MUX_UNSIGNED #(.width(4)) u_mux_435 (
        .y(_node_401),
        .sel(_node_400),
        .a(_T_551_95),
        .b(_node_399)
    );
    wire _node_402;
    EQ_UNSIGNED #(.width(7)) u_eq_436 (
        .y(_node_402),
        .a(7'd96),
        .b(_value__q)
    );
    wire [3:0] _node_403;
    MUX_UNSIGNED #(.width(4)) u_mux_437 (
        .y(_node_403),
        .sel(_node_402),
        .a(_T_551_96),
        .b(_node_401)
    );
    wire _node_404;
    EQ_UNSIGNED #(.width(7)) u_eq_438 (
        .y(_node_404),
        .a(7'd97),
        .b(_value__q)
    );
    wire [3:0] _node_405;
    MUX_UNSIGNED #(.width(4)) u_mux_439 (
        .y(_node_405),
        .sel(_node_404),
        .a(_T_551_97),
        .b(_node_403)
    );
    wire _node_406;
    EQ_UNSIGNED #(.width(7)) u_eq_440 (
        .y(_node_406),
        .a(7'd98),
        .b(_value__q)
    );
    wire [3:0] _node_407;
    MUX_UNSIGNED #(.width(4)) u_mux_441 (
        .y(_node_407),
        .sel(_node_406),
        .a(_T_551_98),
        .b(_node_405)
    );
    wire _node_408;
    EQ_UNSIGNED #(.width(7)) u_eq_442 (
        .y(_node_408),
        .a(7'd99),
        .b(_value__q)
    );
    wire [3:0] _node_409;
    MUX_UNSIGNED #(.width(4)) u_mux_443 (
        .y(_node_409),
        .sel(_node_408),
        .a(_T_551_99),
        .b(_node_407)
    );
    wire _node_410;
    EQ_UNSIGNED #(.width(7)) u_eq_444 (
        .y(_node_410),
        .a(7'd100),
        .b(_value__q)
    );
    wire [3:0] _node_411;
    MUX_UNSIGNED #(.width(4)) u_mux_445 (
        .y(_node_411),
        .sel(_node_410),
        .a(_T_551_100),
        .b(_node_409)
    );
    wire [6:0] _T_658;
    BITS #(.width(9), .high(6), .low(0)) bits_446 (
        .y(_T_658),
        .in(__T_4__q)
    );
    wire _node_412;
    EQ_UNSIGNED #(.width(7)) u_eq_447 (
        .y(_node_412),
        .a(7'd0),
        .b(_T_658)
    );
    wire _node_413;
    assign _node_413 = _T_135_0;
    wire _node_414;
    EQ_UNSIGNED #(.width(7)) u_eq_448 (
        .y(_node_414),
        .a(7'd1),
        .b(_T_658)
    );
    wire _node_415;
    MUX_UNSIGNED #(.width(1)) u_mux_449 (
        .y(_node_415),
        .sel(_node_414),
        .a(_T_135_1),
        .b(_node_413)
    );
    wire _node_416;
    EQ_UNSIGNED #(.width(7)) u_eq_450 (
        .y(_node_416),
        .a(7'd2),
        .b(_T_658)
    );
    wire _node_417;
    MUX_UNSIGNED #(.width(1)) u_mux_451 (
        .y(_node_417),
        .sel(_node_416),
        .a(_T_135_2),
        .b(_node_415)
    );
    wire _node_418;
    EQ_UNSIGNED #(.width(7)) u_eq_452 (
        .y(_node_418),
        .a(7'd3),
        .b(_T_658)
    );
    wire _node_419;
    MUX_UNSIGNED #(.width(1)) u_mux_453 (
        .y(_node_419),
        .sel(_node_418),
        .a(_T_135_3),
        .b(_node_417)
    );
    wire _node_420;
    EQ_UNSIGNED #(.width(7)) u_eq_454 (
        .y(_node_420),
        .a(7'd4),
        .b(_T_658)
    );
    wire _node_421;
    MUX_UNSIGNED #(.width(1)) u_mux_455 (
        .y(_node_421),
        .sel(_node_420),
        .a(_T_135_4),
        .b(_node_419)
    );
    wire _node_422;
    EQ_UNSIGNED #(.width(7)) u_eq_456 (
        .y(_node_422),
        .a(7'd5),
        .b(_T_658)
    );
    wire _node_423;
    MUX_UNSIGNED #(.width(1)) u_mux_457 (
        .y(_node_423),
        .sel(_node_422),
        .a(_T_135_5),
        .b(_node_421)
    );
    wire _node_424;
    EQ_UNSIGNED #(.width(7)) u_eq_458 (
        .y(_node_424),
        .a(7'd6),
        .b(_T_658)
    );
    wire _node_425;
    MUX_UNSIGNED #(.width(1)) u_mux_459 (
        .y(_node_425),
        .sel(_node_424),
        .a(_T_135_6),
        .b(_node_423)
    );
    wire _node_426;
    EQ_UNSIGNED #(.width(7)) u_eq_460 (
        .y(_node_426),
        .a(7'd7),
        .b(_T_658)
    );
    wire _node_427;
    MUX_UNSIGNED #(.width(1)) u_mux_461 (
        .y(_node_427),
        .sel(_node_426),
        .a(_T_135_7),
        .b(_node_425)
    );
    wire _node_428;
    EQ_UNSIGNED #(.width(7)) u_eq_462 (
        .y(_node_428),
        .a(7'd8),
        .b(_T_658)
    );
    wire _node_429;
    MUX_UNSIGNED #(.width(1)) u_mux_463 (
        .y(_node_429),
        .sel(_node_428),
        .a(_T_135_8),
        .b(_node_427)
    );
    wire _node_430;
    EQ_UNSIGNED #(.width(7)) u_eq_464 (
        .y(_node_430),
        .a(7'd9),
        .b(_T_658)
    );
    wire _node_431;
    MUX_UNSIGNED #(.width(1)) u_mux_465 (
        .y(_node_431),
        .sel(_node_430),
        .a(_T_135_9),
        .b(_node_429)
    );
    wire _node_432;
    EQ_UNSIGNED #(.width(7)) u_eq_466 (
        .y(_node_432),
        .a(7'd10),
        .b(_T_658)
    );
    wire _node_433;
    MUX_UNSIGNED #(.width(1)) u_mux_467 (
        .y(_node_433),
        .sel(_node_432),
        .a(_T_135_10),
        .b(_node_431)
    );
    wire _node_434;
    EQ_UNSIGNED #(.width(7)) u_eq_468 (
        .y(_node_434),
        .a(7'd11),
        .b(_T_658)
    );
    wire _node_435;
    MUX_UNSIGNED #(.width(1)) u_mux_469 (
        .y(_node_435),
        .sel(_node_434),
        .a(_T_135_11),
        .b(_node_433)
    );
    wire _node_436;
    EQ_UNSIGNED #(.width(7)) u_eq_470 (
        .y(_node_436),
        .a(7'd12),
        .b(_T_658)
    );
    wire _node_437;
    MUX_UNSIGNED #(.width(1)) u_mux_471 (
        .y(_node_437),
        .sel(_node_436),
        .a(_T_135_12),
        .b(_node_435)
    );
    wire _node_438;
    EQ_UNSIGNED #(.width(7)) u_eq_472 (
        .y(_node_438),
        .a(7'd13),
        .b(_T_658)
    );
    wire _node_439;
    MUX_UNSIGNED #(.width(1)) u_mux_473 (
        .y(_node_439),
        .sel(_node_438),
        .a(_T_135_13),
        .b(_node_437)
    );
    wire _node_440;
    EQ_UNSIGNED #(.width(7)) u_eq_474 (
        .y(_node_440),
        .a(7'd14),
        .b(_T_658)
    );
    wire _node_441;
    MUX_UNSIGNED #(.width(1)) u_mux_475 (
        .y(_node_441),
        .sel(_node_440),
        .a(_T_135_14),
        .b(_node_439)
    );
    wire _node_442;
    EQ_UNSIGNED #(.width(7)) u_eq_476 (
        .y(_node_442),
        .a(7'd15),
        .b(_T_658)
    );
    wire _node_443;
    MUX_UNSIGNED #(.width(1)) u_mux_477 (
        .y(_node_443),
        .sel(_node_442),
        .a(_T_135_15),
        .b(_node_441)
    );
    wire _node_444;
    EQ_UNSIGNED #(.width(7)) u_eq_478 (
        .y(_node_444),
        .a(7'd16),
        .b(_T_658)
    );
    wire _node_445;
    MUX_UNSIGNED #(.width(1)) u_mux_479 (
        .y(_node_445),
        .sel(_node_444),
        .a(_T_135_16),
        .b(_node_443)
    );
    wire _node_446;
    EQ_UNSIGNED #(.width(7)) u_eq_480 (
        .y(_node_446),
        .a(7'd17),
        .b(_T_658)
    );
    wire _node_447;
    MUX_UNSIGNED #(.width(1)) u_mux_481 (
        .y(_node_447),
        .sel(_node_446),
        .a(_T_135_17),
        .b(_node_445)
    );
    wire _node_448;
    EQ_UNSIGNED #(.width(7)) u_eq_482 (
        .y(_node_448),
        .a(7'd18),
        .b(_T_658)
    );
    wire _node_449;
    MUX_UNSIGNED #(.width(1)) u_mux_483 (
        .y(_node_449),
        .sel(_node_448),
        .a(_T_135_18),
        .b(_node_447)
    );
    wire _node_450;
    EQ_UNSIGNED #(.width(7)) u_eq_484 (
        .y(_node_450),
        .a(7'd19),
        .b(_T_658)
    );
    wire _node_451;
    MUX_UNSIGNED #(.width(1)) u_mux_485 (
        .y(_node_451),
        .sel(_node_450),
        .a(_T_135_19),
        .b(_node_449)
    );
    wire _node_452;
    EQ_UNSIGNED #(.width(7)) u_eq_486 (
        .y(_node_452),
        .a(7'd20),
        .b(_T_658)
    );
    wire _node_453;
    MUX_UNSIGNED #(.width(1)) u_mux_487 (
        .y(_node_453),
        .sel(_node_452),
        .a(_T_135_20),
        .b(_node_451)
    );
    wire _node_454;
    EQ_UNSIGNED #(.width(7)) u_eq_488 (
        .y(_node_454),
        .a(7'd21),
        .b(_T_658)
    );
    wire _node_455;
    MUX_UNSIGNED #(.width(1)) u_mux_489 (
        .y(_node_455),
        .sel(_node_454),
        .a(_T_135_21),
        .b(_node_453)
    );
    wire _node_456;
    EQ_UNSIGNED #(.width(7)) u_eq_490 (
        .y(_node_456),
        .a(7'd22),
        .b(_T_658)
    );
    wire _node_457;
    MUX_UNSIGNED #(.width(1)) u_mux_491 (
        .y(_node_457),
        .sel(_node_456),
        .a(_T_135_22),
        .b(_node_455)
    );
    wire _node_458;
    EQ_UNSIGNED #(.width(7)) u_eq_492 (
        .y(_node_458),
        .a(7'd23),
        .b(_T_658)
    );
    wire _node_459;
    MUX_UNSIGNED #(.width(1)) u_mux_493 (
        .y(_node_459),
        .sel(_node_458),
        .a(_T_135_23),
        .b(_node_457)
    );
    wire _node_460;
    EQ_UNSIGNED #(.width(7)) u_eq_494 (
        .y(_node_460),
        .a(7'd24),
        .b(_T_658)
    );
    wire _node_461;
    MUX_UNSIGNED #(.width(1)) u_mux_495 (
        .y(_node_461),
        .sel(_node_460),
        .a(_T_135_24),
        .b(_node_459)
    );
    wire _node_462;
    EQ_UNSIGNED #(.width(7)) u_eq_496 (
        .y(_node_462),
        .a(7'd25),
        .b(_T_658)
    );
    wire _node_463;
    MUX_UNSIGNED #(.width(1)) u_mux_497 (
        .y(_node_463),
        .sel(_node_462),
        .a(_T_135_25),
        .b(_node_461)
    );
    wire _node_464;
    EQ_UNSIGNED #(.width(7)) u_eq_498 (
        .y(_node_464),
        .a(7'd26),
        .b(_T_658)
    );
    wire _node_465;
    MUX_UNSIGNED #(.width(1)) u_mux_499 (
        .y(_node_465),
        .sel(_node_464),
        .a(_T_135_26),
        .b(_node_463)
    );
    wire _node_466;
    EQ_UNSIGNED #(.width(7)) u_eq_500 (
        .y(_node_466),
        .a(7'd27),
        .b(_T_658)
    );
    wire _node_467;
    MUX_UNSIGNED #(.width(1)) u_mux_501 (
        .y(_node_467),
        .sel(_node_466),
        .a(_T_135_27),
        .b(_node_465)
    );
    wire _node_468;
    EQ_UNSIGNED #(.width(7)) u_eq_502 (
        .y(_node_468),
        .a(7'd28),
        .b(_T_658)
    );
    wire _node_469;
    MUX_UNSIGNED #(.width(1)) u_mux_503 (
        .y(_node_469),
        .sel(_node_468),
        .a(_T_135_28),
        .b(_node_467)
    );
    wire _node_470;
    EQ_UNSIGNED #(.width(7)) u_eq_504 (
        .y(_node_470),
        .a(7'd29),
        .b(_T_658)
    );
    wire _node_471;
    MUX_UNSIGNED #(.width(1)) u_mux_505 (
        .y(_node_471),
        .sel(_node_470),
        .a(_T_135_29),
        .b(_node_469)
    );
    wire _node_472;
    EQ_UNSIGNED #(.width(7)) u_eq_506 (
        .y(_node_472),
        .a(7'd30),
        .b(_T_658)
    );
    wire _node_473;
    MUX_UNSIGNED #(.width(1)) u_mux_507 (
        .y(_node_473),
        .sel(_node_472),
        .a(_T_135_30),
        .b(_node_471)
    );
    wire _node_474;
    EQ_UNSIGNED #(.width(7)) u_eq_508 (
        .y(_node_474),
        .a(7'd31),
        .b(_T_658)
    );
    wire _node_475;
    MUX_UNSIGNED #(.width(1)) u_mux_509 (
        .y(_node_475),
        .sel(_node_474),
        .a(_T_135_31),
        .b(_node_473)
    );
    wire _node_476;
    EQ_UNSIGNED #(.width(7)) u_eq_510 (
        .y(_node_476),
        .a(7'd32),
        .b(_T_658)
    );
    wire _node_477;
    MUX_UNSIGNED #(.width(1)) u_mux_511 (
        .y(_node_477),
        .sel(_node_476),
        .a(_T_135_32),
        .b(_node_475)
    );
    wire _node_478;
    EQ_UNSIGNED #(.width(7)) u_eq_512 (
        .y(_node_478),
        .a(7'd33),
        .b(_T_658)
    );
    wire _node_479;
    MUX_UNSIGNED #(.width(1)) u_mux_513 (
        .y(_node_479),
        .sel(_node_478),
        .a(_T_135_33),
        .b(_node_477)
    );
    wire _node_480;
    EQ_UNSIGNED #(.width(7)) u_eq_514 (
        .y(_node_480),
        .a(7'd34),
        .b(_T_658)
    );
    wire _node_481;
    MUX_UNSIGNED #(.width(1)) u_mux_515 (
        .y(_node_481),
        .sel(_node_480),
        .a(_T_135_34),
        .b(_node_479)
    );
    wire _node_482;
    EQ_UNSIGNED #(.width(7)) u_eq_516 (
        .y(_node_482),
        .a(7'd35),
        .b(_T_658)
    );
    wire _node_483;
    MUX_UNSIGNED #(.width(1)) u_mux_517 (
        .y(_node_483),
        .sel(_node_482),
        .a(_T_135_35),
        .b(_node_481)
    );
    wire _node_484;
    EQ_UNSIGNED #(.width(7)) u_eq_518 (
        .y(_node_484),
        .a(7'd36),
        .b(_T_658)
    );
    wire _node_485;
    MUX_UNSIGNED #(.width(1)) u_mux_519 (
        .y(_node_485),
        .sel(_node_484),
        .a(_T_135_36),
        .b(_node_483)
    );
    wire _node_486;
    EQ_UNSIGNED #(.width(7)) u_eq_520 (
        .y(_node_486),
        .a(7'd37),
        .b(_T_658)
    );
    wire _node_487;
    MUX_UNSIGNED #(.width(1)) u_mux_521 (
        .y(_node_487),
        .sel(_node_486),
        .a(_T_135_37),
        .b(_node_485)
    );
    wire _node_488;
    EQ_UNSIGNED #(.width(7)) u_eq_522 (
        .y(_node_488),
        .a(7'd38),
        .b(_T_658)
    );
    wire _node_489;
    MUX_UNSIGNED #(.width(1)) u_mux_523 (
        .y(_node_489),
        .sel(_node_488),
        .a(_T_135_38),
        .b(_node_487)
    );
    wire _node_490;
    EQ_UNSIGNED #(.width(7)) u_eq_524 (
        .y(_node_490),
        .a(7'd39),
        .b(_T_658)
    );
    wire _node_491;
    MUX_UNSIGNED #(.width(1)) u_mux_525 (
        .y(_node_491),
        .sel(_node_490),
        .a(_T_135_39),
        .b(_node_489)
    );
    wire _node_492;
    EQ_UNSIGNED #(.width(7)) u_eq_526 (
        .y(_node_492),
        .a(7'd40),
        .b(_T_658)
    );
    wire _node_493;
    MUX_UNSIGNED #(.width(1)) u_mux_527 (
        .y(_node_493),
        .sel(_node_492),
        .a(_T_135_40),
        .b(_node_491)
    );
    wire _node_494;
    EQ_UNSIGNED #(.width(7)) u_eq_528 (
        .y(_node_494),
        .a(7'd41),
        .b(_T_658)
    );
    wire _node_495;
    MUX_UNSIGNED #(.width(1)) u_mux_529 (
        .y(_node_495),
        .sel(_node_494),
        .a(_T_135_41),
        .b(_node_493)
    );
    wire _node_496;
    EQ_UNSIGNED #(.width(7)) u_eq_530 (
        .y(_node_496),
        .a(7'd42),
        .b(_T_658)
    );
    wire _node_497;
    MUX_UNSIGNED #(.width(1)) u_mux_531 (
        .y(_node_497),
        .sel(_node_496),
        .a(_T_135_42),
        .b(_node_495)
    );
    wire _node_498;
    EQ_UNSIGNED #(.width(7)) u_eq_532 (
        .y(_node_498),
        .a(7'd43),
        .b(_T_658)
    );
    wire _node_499;
    MUX_UNSIGNED #(.width(1)) u_mux_533 (
        .y(_node_499),
        .sel(_node_498),
        .a(_T_135_43),
        .b(_node_497)
    );
    wire _node_500;
    EQ_UNSIGNED #(.width(7)) u_eq_534 (
        .y(_node_500),
        .a(7'd44),
        .b(_T_658)
    );
    wire _node_501;
    MUX_UNSIGNED #(.width(1)) u_mux_535 (
        .y(_node_501),
        .sel(_node_500),
        .a(_T_135_44),
        .b(_node_499)
    );
    wire _node_502;
    EQ_UNSIGNED #(.width(7)) u_eq_536 (
        .y(_node_502),
        .a(7'd45),
        .b(_T_658)
    );
    wire _node_503;
    MUX_UNSIGNED #(.width(1)) u_mux_537 (
        .y(_node_503),
        .sel(_node_502),
        .a(_T_135_45),
        .b(_node_501)
    );
    wire _node_504;
    EQ_UNSIGNED #(.width(7)) u_eq_538 (
        .y(_node_504),
        .a(7'd46),
        .b(_T_658)
    );
    wire _node_505;
    MUX_UNSIGNED #(.width(1)) u_mux_539 (
        .y(_node_505),
        .sel(_node_504),
        .a(_T_135_46),
        .b(_node_503)
    );
    wire _node_506;
    EQ_UNSIGNED #(.width(7)) u_eq_540 (
        .y(_node_506),
        .a(7'd47),
        .b(_T_658)
    );
    wire _node_507;
    MUX_UNSIGNED #(.width(1)) u_mux_541 (
        .y(_node_507),
        .sel(_node_506),
        .a(_T_135_47),
        .b(_node_505)
    );
    wire _node_508;
    EQ_UNSIGNED #(.width(7)) u_eq_542 (
        .y(_node_508),
        .a(7'd48),
        .b(_T_658)
    );
    wire _node_509;
    MUX_UNSIGNED #(.width(1)) u_mux_543 (
        .y(_node_509),
        .sel(_node_508),
        .a(_T_135_48),
        .b(_node_507)
    );
    wire _node_510;
    EQ_UNSIGNED #(.width(7)) u_eq_544 (
        .y(_node_510),
        .a(7'd49),
        .b(_T_658)
    );
    wire _node_511;
    MUX_UNSIGNED #(.width(1)) u_mux_545 (
        .y(_node_511),
        .sel(_node_510),
        .a(_T_135_49),
        .b(_node_509)
    );
    wire _node_512;
    EQ_UNSIGNED #(.width(7)) u_eq_546 (
        .y(_node_512),
        .a(7'd50),
        .b(_T_658)
    );
    wire _node_513;
    MUX_UNSIGNED #(.width(1)) u_mux_547 (
        .y(_node_513),
        .sel(_node_512),
        .a(_T_135_50),
        .b(_node_511)
    );
    wire _node_514;
    EQ_UNSIGNED #(.width(7)) u_eq_548 (
        .y(_node_514),
        .a(7'd51),
        .b(_T_658)
    );
    wire _node_515;
    MUX_UNSIGNED #(.width(1)) u_mux_549 (
        .y(_node_515),
        .sel(_node_514),
        .a(_T_135_51),
        .b(_node_513)
    );
    wire _node_516;
    EQ_UNSIGNED #(.width(7)) u_eq_550 (
        .y(_node_516),
        .a(7'd52),
        .b(_T_658)
    );
    wire _node_517;
    MUX_UNSIGNED #(.width(1)) u_mux_551 (
        .y(_node_517),
        .sel(_node_516),
        .a(_T_135_52),
        .b(_node_515)
    );
    wire _node_518;
    EQ_UNSIGNED #(.width(7)) u_eq_552 (
        .y(_node_518),
        .a(7'd53),
        .b(_T_658)
    );
    wire _node_519;
    MUX_UNSIGNED #(.width(1)) u_mux_553 (
        .y(_node_519),
        .sel(_node_518),
        .a(_T_135_53),
        .b(_node_517)
    );
    wire _node_520;
    EQ_UNSIGNED #(.width(7)) u_eq_554 (
        .y(_node_520),
        .a(7'd54),
        .b(_T_658)
    );
    wire _node_521;
    MUX_UNSIGNED #(.width(1)) u_mux_555 (
        .y(_node_521),
        .sel(_node_520),
        .a(_T_135_54),
        .b(_node_519)
    );
    wire _node_522;
    EQ_UNSIGNED #(.width(7)) u_eq_556 (
        .y(_node_522),
        .a(7'd55),
        .b(_T_658)
    );
    wire _node_523;
    MUX_UNSIGNED #(.width(1)) u_mux_557 (
        .y(_node_523),
        .sel(_node_522),
        .a(_T_135_55),
        .b(_node_521)
    );
    wire _node_524;
    EQ_UNSIGNED #(.width(7)) u_eq_558 (
        .y(_node_524),
        .a(7'd56),
        .b(_T_658)
    );
    wire _node_525;
    MUX_UNSIGNED #(.width(1)) u_mux_559 (
        .y(_node_525),
        .sel(_node_524),
        .a(_T_135_56),
        .b(_node_523)
    );
    wire _node_526;
    EQ_UNSIGNED #(.width(7)) u_eq_560 (
        .y(_node_526),
        .a(7'd57),
        .b(_T_658)
    );
    wire _node_527;
    MUX_UNSIGNED #(.width(1)) u_mux_561 (
        .y(_node_527),
        .sel(_node_526),
        .a(_T_135_57),
        .b(_node_525)
    );
    wire _node_528;
    EQ_UNSIGNED #(.width(7)) u_eq_562 (
        .y(_node_528),
        .a(7'd58),
        .b(_T_658)
    );
    wire _node_529;
    MUX_UNSIGNED #(.width(1)) u_mux_563 (
        .y(_node_529),
        .sel(_node_528),
        .a(_T_135_58),
        .b(_node_527)
    );
    wire _node_530;
    EQ_UNSIGNED #(.width(7)) u_eq_564 (
        .y(_node_530),
        .a(7'd59),
        .b(_T_658)
    );
    wire _node_531;
    MUX_UNSIGNED #(.width(1)) u_mux_565 (
        .y(_node_531),
        .sel(_node_530),
        .a(_T_135_59),
        .b(_node_529)
    );
    wire _node_532;
    EQ_UNSIGNED #(.width(7)) u_eq_566 (
        .y(_node_532),
        .a(7'd60),
        .b(_T_658)
    );
    wire _node_533;
    MUX_UNSIGNED #(.width(1)) u_mux_567 (
        .y(_node_533),
        .sel(_node_532),
        .a(_T_135_60),
        .b(_node_531)
    );
    wire _node_534;
    EQ_UNSIGNED #(.width(7)) u_eq_568 (
        .y(_node_534),
        .a(7'd61),
        .b(_T_658)
    );
    wire _node_535;
    MUX_UNSIGNED #(.width(1)) u_mux_569 (
        .y(_node_535),
        .sel(_node_534),
        .a(_T_135_61),
        .b(_node_533)
    );
    wire _node_536;
    EQ_UNSIGNED #(.width(7)) u_eq_570 (
        .y(_node_536),
        .a(7'd62),
        .b(_T_658)
    );
    wire _node_537;
    MUX_UNSIGNED #(.width(1)) u_mux_571 (
        .y(_node_537),
        .sel(_node_536),
        .a(_T_135_62),
        .b(_node_535)
    );
    wire _node_538;
    EQ_UNSIGNED #(.width(7)) u_eq_572 (
        .y(_node_538),
        .a(7'd63),
        .b(_T_658)
    );
    wire _node_539;
    MUX_UNSIGNED #(.width(1)) u_mux_573 (
        .y(_node_539),
        .sel(_node_538),
        .a(_T_135_63),
        .b(_node_537)
    );
    wire _node_540;
    EQ_UNSIGNED #(.width(7)) u_eq_574 (
        .y(_node_540),
        .a(7'd64),
        .b(_T_658)
    );
    wire _node_541;
    MUX_UNSIGNED #(.width(1)) u_mux_575 (
        .y(_node_541),
        .sel(_node_540),
        .a(_T_135_64),
        .b(_node_539)
    );
    wire _node_542;
    EQ_UNSIGNED #(.width(7)) u_eq_576 (
        .y(_node_542),
        .a(7'd65),
        .b(_T_658)
    );
    wire _node_543;
    MUX_UNSIGNED #(.width(1)) u_mux_577 (
        .y(_node_543),
        .sel(_node_542),
        .a(_T_135_65),
        .b(_node_541)
    );
    wire _node_544;
    EQ_UNSIGNED #(.width(7)) u_eq_578 (
        .y(_node_544),
        .a(7'd66),
        .b(_T_658)
    );
    wire _node_545;
    MUX_UNSIGNED #(.width(1)) u_mux_579 (
        .y(_node_545),
        .sel(_node_544),
        .a(_T_135_66),
        .b(_node_543)
    );
    wire _node_546;
    EQ_UNSIGNED #(.width(7)) u_eq_580 (
        .y(_node_546),
        .a(7'd67),
        .b(_T_658)
    );
    wire _node_547;
    MUX_UNSIGNED #(.width(1)) u_mux_581 (
        .y(_node_547),
        .sel(_node_546),
        .a(_T_135_67),
        .b(_node_545)
    );
    wire _node_548;
    EQ_UNSIGNED #(.width(7)) u_eq_582 (
        .y(_node_548),
        .a(7'd68),
        .b(_T_658)
    );
    wire _node_549;
    MUX_UNSIGNED #(.width(1)) u_mux_583 (
        .y(_node_549),
        .sel(_node_548),
        .a(_T_135_68),
        .b(_node_547)
    );
    wire _node_550;
    EQ_UNSIGNED #(.width(7)) u_eq_584 (
        .y(_node_550),
        .a(7'd69),
        .b(_T_658)
    );
    wire _node_551;
    MUX_UNSIGNED #(.width(1)) u_mux_585 (
        .y(_node_551),
        .sel(_node_550),
        .a(_T_135_69),
        .b(_node_549)
    );
    wire _node_552;
    EQ_UNSIGNED #(.width(7)) u_eq_586 (
        .y(_node_552),
        .a(7'd70),
        .b(_T_658)
    );
    wire _node_553;
    MUX_UNSIGNED #(.width(1)) u_mux_587 (
        .y(_node_553),
        .sel(_node_552),
        .a(_T_135_70),
        .b(_node_551)
    );
    wire _node_554;
    EQ_UNSIGNED #(.width(7)) u_eq_588 (
        .y(_node_554),
        .a(7'd71),
        .b(_T_658)
    );
    wire _node_555;
    MUX_UNSIGNED #(.width(1)) u_mux_589 (
        .y(_node_555),
        .sel(_node_554),
        .a(_T_135_71),
        .b(_node_553)
    );
    wire _node_556;
    EQ_UNSIGNED #(.width(7)) u_eq_590 (
        .y(_node_556),
        .a(7'd72),
        .b(_T_658)
    );
    wire _node_557;
    MUX_UNSIGNED #(.width(1)) u_mux_591 (
        .y(_node_557),
        .sel(_node_556),
        .a(_T_135_72),
        .b(_node_555)
    );
    wire _node_558;
    EQ_UNSIGNED #(.width(7)) u_eq_592 (
        .y(_node_558),
        .a(7'd73),
        .b(_T_658)
    );
    wire _node_559;
    MUX_UNSIGNED #(.width(1)) u_mux_593 (
        .y(_node_559),
        .sel(_node_558),
        .a(_T_135_73),
        .b(_node_557)
    );
    wire _node_560;
    EQ_UNSIGNED #(.width(7)) u_eq_594 (
        .y(_node_560),
        .a(7'd74),
        .b(_T_658)
    );
    wire _node_561;
    MUX_UNSIGNED #(.width(1)) u_mux_595 (
        .y(_node_561),
        .sel(_node_560),
        .a(_T_135_74),
        .b(_node_559)
    );
    wire _node_562;
    EQ_UNSIGNED #(.width(7)) u_eq_596 (
        .y(_node_562),
        .a(7'd75),
        .b(_T_658)
    );
    wire _node_563;
    MUX_UNSIGNED #(.width(1)) u_mux_597 (
        .y(_node_563),
        .sel(_node_562),
        .a(_T_135_75),
        .b(_node_561)
    );
    wire _node_564;
    EQ_UNSIGNED #(.width(7)) u_eq_598 (
        .y(_node_564),
        .a(7'd76),
        .b(_T_658)
    );
    wire _node_565;
    MUX_UNSIGNED #(.width(1)) u_mux_599 (
        .y(_node_565),
        .sel(_node_564),
        .a(_T_135_76),
        .b(_node_563)
    );
    wire _node_566;
    EQ_UNSIGNED #(.width(7)) u_eq_600 (
        .y(_node_566),
        .a(7'd77),
        .b(_T_658)
    );
    wire _node_567;
    MUX_UNSIGNED #(.width(1)) u_mux_601 (
        .y(_node_567),
        .sel(_node_566),
        .a(_T_135_77),
        .b(_node_565)
    );
    wire _node_568;
    EQ_UNSIGNED #(.width(7)) u_eq_602 (
        .y(_node_568),
        .a(7'd78),
        .b(_T_658)
    );
    wire _node_569;
    MUX_UNSIGNED #(.width(1)) u_mux_603 (
        .y(_node_569),
        .sel(_node_568),
        .a(_T_135_78),
        .b(_node_567)
    );
    wire _node_570;
    EQ_UNSIGNED #(.width(7)) u_eq_604 (
        .y(_node_570),
        .a(7'd79),
        .b(_T_658)
    );
    wire _node_571;
    MUX_UNSIGNED #(.width(1)) u_mux_605 (
        .y(_node_571),
        .sel(_node_570),
        .a(_T_135_79),
        .b(_node_569)
    );
    wire _node_572;
    EQ_UNSIGNED #(.width(7)) u_eq_606 (
        .y(_node_572),
        .a(7'd80),
        .b(_T_658)
    );
    wire _node_573;
    MUX_UNSIGNED #(.width(1)) u_mux_607 (
        .y(_node_573),
        .sel(_node_572),
        .a(_T_135_80),
        .b(_node_571)
    );
    wire _node_574;
    EQ_UNSIGNED #(.width(7)) u_eq_608 (
        .y(_node_574),
        .a(7'd81),
        .b(_T_658)
    );
    wire _node_575;
    MUX_UNSIGNED #(.width(1)) u_mux_609 (
        .y(_node_575),
        .sel(_node_574),
        .a(_T_135_81),
        .b(_node_573)
    );
    wire _node_576;
    EQ_UNSIGNED #(.width(7)) u_eq_610 (
        .y(_node_576),
        .a(7'd82),
        .b(_T_658)
    );
    wire _node_577;
    MUX_UNSIGNED #(.width(1)) u_mux_611 (
        .y(_node_577),
        .sel(_node_576),
        .a(_T_135_82),
        .b(_node_575)
    );
    wire _node_578;
    EQ_UNSIGNED #(.width(7)) u_eq_612 (
        .y(_node_578),
        .a(7'd83),
        .b(_T_658)
    );
    wire _node_579;
    MUX_UNSIGNED #(.width(1)) u_mux_613 (
        .y(_node_579),
        .sel(_node_578),
        .a(_T_135_83),
        .b(_node_577)
    );
    wire _node_580;
    EQ_UNSIGNED #(.width(7)) u_eq_614 (
        .y(_node_580),
        .a(7'd84),
        .b(_T_658)
    );
    wire _node_581;
    MUX_UNSIGNED #(.width(1)) u_mux_615 (
        .y(_node_581),
        .sel(_node_580),
        .a(_T_135_84),
        .b(_node_579)
    );
    wire _node_582;
    EQ_UNSIGNED #(.width(7)) u_eq_616 (
        .y(_node_582),
        .a(7'd85),
        .b(_T_658)
    );
    wire _node_583;
    MUX_UNSIGNED #(.width(1)) u_mux_617 (
        .y(_node_583),
        .sel(_node_582),
        .a(_T_135_85),
        .b(_node_581)
    );
    wire _node_584;
    EQ_UNSIGNED #(.width(7)) u_eq_618 (
        .y(_node_584),
        .a(7'd86),
        .b(_T_658)
    );
    wire _node_585;
    MUX_UNSIGNED #(.width(1)) u_mux_619 (
        .y(_node_585),
        .sel(_node_584),
        .a(_T_135_86),
        .b(_node_583)
    );
    wire _node_586;
    EQ_UNSIGNED #(.width(7)) u_eq_620 (
        .y(_node_586),
        .a(7'd87),
        .b(_T_658)
    );
    wire _node_587;
    MUX_UNSIGNED #(.width(1)) u_mux_621 (
        .y(_node_587),
        .sel(_node_586),
        .a(_T_135_87),
        .b(_node_585)
    );
    wire _node_588;
    EQ_UNSIGNED #(.width(7)) u_eq_622 (
        .y(_node_588),
        .a(7'd88),
        .b(_T_658)
    );
    wire _node_589;
    MUX_UNSIGNED #(.width(1)) u_mux_623 (
        .y(_node_589),
        .sel(_node_588),
        .a(_T_135_88),
        .b(_node_587)
    );
    wire _node_590;
    EQ_UNSIGNED #(.width(7)) u_eq_624 (
        .y(_node_590),
        .a(7'd89),
        .b(_T_658)
    );
    wire _node_591;
    MUX_UNSIGNED #(.width(1)) u_mux_625 (
        .y(_node_591),
        .sel(_node_590),
        .a(_T_135_89),
        .b(_node_589)
    );
    wire _node_592;
    EQ_UNSIGNED #(.width(7)) u_eq_626 (
        .y(_node_592),
        .a(7'd90),
        .b(_T_658)
    );
    wire _node_593;
    MUX_UNSIGNED #(.width(1)) u_mux_627 (
        .y(_node_593),
        .sel(_node_592),
        .a(_T_135_90),
        .b(_node_591)
    );
    wire _node_594;
    EQ_UNSIGNED #(.width(7)) u_eq_628 (
        .y(_node_594),
        .a(7'd91),
        .b(_T_658)
    );
    wire _node_595;
    MUX_UNSIGNED #(.width(1)) u_mux_629 (
        .y(_node_595),
        .sel(_node_594),
        .a(_T_135_91),
        .b(_node_593)
    );
    wire _node_596;
    EQ_UNSIGNED #(.width(7)) u_eq_630 (
        .y(_node_596),
        .a(7'd92),
        .b(_T_658)
    );
    wire _node_597;
    MUX_UNSIGNED #(.width(1)) u_mux_631 (
        .y(_node_597),
        .sel(_node_596),
        .a(_T_135_92),
        .b(_node_595)
    );
    wire _node_598;
    EQ_UNSIGNED #(.width(7)) u_eq_632 (
        .y(_node_598),
        .a(7'd93),
        .b(_T_658)
    );
    wire _node_599;
    MUX_UNSIGNED #(.width(1)) u_mux_633 (
        .y(_node_599),
        .sel(_node_598),
        .a(_T_135_93),
        .b(_node_597)
    );
    wire _node_600;
    EQ_UNSIGNED #(.width(7)) u_eq_634 (
        .y(_node_600),
        .a(7'd94),
        .b(_T_658)
    );
    wire _node_601;
    MUX_UNSIGNED #(.width(1)) u_mux_635 (
        .y(_node_601),
        .sel(_node_600),
        .a(_T_135_94),
        .b(_node_599)
    );
    wire _node_602;
    EQ_UNSIGNED #(.width(7)) u_eq_636 (
        .y(_node_602),
        .a(7'd95),
        .b(_T_658)
    );
    wire _node_603;
    MUX_UNSIGNED #(.width(1)) u_mux_637 (
        .y(_node_603),
        .sel(_node_602),
        .a(_T_135_95),
        .b(_node_601)
    );
    wire _node_604;
    EQ_UNSIGNED #(.width(7)) u_eq_638 (
        .y(_node_604),
        .a(7'd96),
        .b(_T_658)
    );
    wire _node_605;
    MUX_UNSIGNED #(.width(1)) u_mux_639 (
        .y(_node_605),
        .sel(_node_604),
        .a(_T_135_96),
        .b(_node_603)
    );
    wire _node_606;
    EQ_UNSIGNED #(.width(7)) u_eq_640 (
        .y(_node_606),
        .a(7'd97),
        .b(_T_658)
    );
    wire _node_607;
    MUX_UNSIGNED #(.width(1)) u_mux_641 (
        .y(_node_607),
        .sel(_node_606),
        .a(_T_135_97),
        .b(_node_605)
    );
    wire _node_608;
    EQ_UNSIGNED #(.width(7)) u_eq_642 (
        .y(_node_608),
        .a(7'd98),
        .b(_T_658)
    );
    wire _node_609;
    MUX_UNSIGNED #(.width(1)) u_mux_643 (
        .y(_node_609),
        .sel(_node_608),
        .a(_T_135_98),
        .b(_node_607)
    );
    wire _node_610;
    EQ_UNSIGNED #(.width(7)) u_eq_644 (
        .y(_node_610),
        .a(7'd99),
        .b(_T_658)
    );
    wire _node_611;
    MUX_UNSIGNED #(.width(1)) u_mux_645 (
        .y(_node_611),
        .sel(_node_610),
        .a(_T_135_99),
        .b(_node_609)
    );
    wire _node_612;
    EQ_UNSIGNED #(.width(7)) u_eq_646 (
        .y(_node_612),
        .a(7'd100),
        .b(_T_658)
    );
    wire _node_613;
    MUX_UNSIGNED #(.width(1)) u_mux_647 (
        .y(_node_613),
        .sel(_node_612),
        .a(_T_135_100),
        .b(_node_611)
    );
    wire _T_659;
    BITWISEAND #(.width(1)) bitwiseand_648 (
        .y(_T_659),
        .a(_c__io_in_valid),
        .b(_c__io_in_ready)
    );
    wire _T_661;
    EQ_UNSIGNED #(.width(7)) u_eq_649 (
        .y(_T_661),
        .a(_value__q),
        .b(7'h63)
    );
    wire [7:0] _T_663;
    wire [6:0] _WTEMP_11;
    PAD_UNSIGNED #(.width(1), .n(7)) u_pad_650 (
        .y(_WTEMP_11),
        .in(1'h1)
    );
    ADD_UNSIGNED #(.width(7)) u_add_651 (
        .y(_T_663),
        .a(_value__q),
        .b(_WTEMP_11)
    );
    wire [6:0] _T_664;
    TAIL #(.width(8), .n(1)) tail_652 (
        .y(_T_664),
        .in(_T_663)
    );
    wire _T_667;
    EQ_UNSIGNED #(.width(1)) u_eq_653 (
        .y(_T_667),
        .a(__T_7__q),
        .b(1'h0)
    );
    wire _T_669;
    wire [8:0] _WTEMP_12;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_654 (
        .y(_WTEMP_12),
        .in(7'h63)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_655 (
        .y(_T_669),
        .a(__T_4__q),
        .b(_WTEMP_12)
    );
    wire [9:0] _T_672;
    wire [8:0] _WTEMP_13;
    PAD_UNSIGNED #(.width(1), .n(9)) u_pad_656 (
        .y(_WTEMP_13),
        .in(1'h1)
    );
    ADD_UNSIGNED #(.width(9)) u_add_657 (
        .y(_T_672),
        .a(__T_4__q),
        .b(_WTEMP_13)
    );
    wire [8:0] _T_673;
    TAIL #(.width(10), .n(1)) tail_658 (
        .y(_T_673),
        .in(_T_672)
    );
    wire _node_614;
    MUX_UNSIGNED #(.width(1)) u_mux_659 (
        .y(_node_614),
        .sel(_T_669),
        .a(1'h1),
        .b(__T_7__q)
    );
    wire [8:0] _node_615;
    MUX_UNSIGNED #(.width(9)) u_mux_660 (
        .y(_node_615),
        .sel(_T_667),
        .a(_T_673),
        .b(__T_4__q)
    );
    wire _node_616;
    MUX_UNSIGNED #(.width(1)) u_mux_661 (
        .y(_node_616),
        .sel(_T_667),
        .a(_node_614),
        .b(__T_7__q)
    );
    wire [6:0] _node_617;
    wire [6:0] _WTEMP_14;
    PAD_UNSIGNED #(.width(1), .n(7)) u_pad_662 (
        .y(_WTEMP_14),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(7)) u_mux_663 (
        .y(_node_617),
        .sel(_T_661),
        .a(_WTEMP_14),
        .b(_T_664)
    );
    wire _T_777_0;
    wire _T_777_1;
    wire _T_777_2;
    wire _T_777_3;
    wire _T_777_4;
    wire _T_777_5;
    wire _T_777_6;
    wire _T_777_7;
    wire _T_777_8;
    wire _T_777_9;
    wire _T_777_10;
    wire _T_777_11;
    wire _T_777_12;
    wire _T_777_13;
    wire _T_777_14;
    wire _T_777_15;
    wire _T_777_16;
    wire _T_777_17;
    wire _T_777_18;
    wire _T_777_19;
    wire _T_777_20;
    wire _T_777_21;
    wire _T_777_22;
    wire _T_777_23;
    wire _T_777_24;
    wire _T_777_25;
    wire _T_777_26;
    wire _T_777_27;
    wire _T_777_28;
    wire _T_777_29;
    wire _T_777_30;
    wire _T_777_31;
    wire _T_777_32;
    wire _T_777_33;
    wire _T_777_34;
    wire _T_777_35;
    wire _T_777_36;
    wire _T_777_37;
    wire _T_777_38;
    wire _T_777_39;
    wire _T_777_40;
    wire _T_777_41;
    wire _T_777_42;
    wire _T_777_43;
    wire _T_777_44;
    wire _T_777_45;
    wire _T_777_46;
    wire _T_777_47;
    wire _T_777_48;
    wire _T_777_49;
    wire _T_777_50;
    wire _T_777_51;
    wire _T_777_52;
    wire _T_777_53;
    wire _T_777_54;
    wire _T_777_55;
    wire _T_777_56;
    wire _T_777_57;
    wire _T_777_58;
    wire _T_777_59;
    wire _T_777_60;
    wire _T_777_61;
    wire _T_777_62;
    wire _T_777_63;
    wire _T_777_64;
    wire _T_777_65;
    wire _T_777_66;
    wire _T_777_67;
    wire _T_777_68;
    wire _T_777_69;
    wire _T_777_70;
    wire _T_777_71;
    wire _T_777_72;
    wire _T_777_73;
    wire _T_777_74;
    wire _T_777_75;
    wire _T_777_76;
    wire _T_777_77;
    wire _T_777_78;
    wire _T_777_79;
    wire _T_777_80;
    wire _T_777_81;
    wire _T_777_82;
    wire _T_777_83;
    wire _T_777_84;
    wire _T_777_85;
    wire _T_777_86;
    wire _T_777_87;
    wire _T_777_88;
    wire _T_777_89;
    wire _T_777_90;
    wire _T_777_91;
    wire _T_777_92;
    wire _T_777_93;
    wire _T_777_94;
    wire _T_777_95;
    wire _T_777_96;
    wire _T_777_97;
    wire _T_777_98;
    wire _T_777_99;
    wire _T_777_100;
    wire [6:0] _value_1__q;
    wire [6:0] _value_1__d;
    DFF_POSCLK #(.width(7)) value_1 (
        .q(_value_1__q),
        .d(_value_1__d),
        .clk(clock)
    );
    wire [6:0] _WTEMP_15;
    MUX_UNSIGNED #(.width(7)) u_mux_664 (
        .y(_value_1__d),
        .sel(reset),
        .a(7'h0),
        .b(_WTEMP_15)
    );
    wire [3:0] _T_986_0;
    wire [3:0] _T_986_1;
    wire [3:0] _T_986_2;
    wire [3:0] _T_986_3;
    wire [3:0] _T_986_4;
    wire [3:0] _T_986_5;
    wire [3:0] _T_986_6;
    wire [3:0] _T_986_7;
    wire [3:0] _T_986_8;
    wire [3:0] _T_986_9;
    wire [3:0] _T_986_10;
    wire [3:0] _T_986_11;
    wire [3:0] _T_986_12;
    wire [3:0] _T_986_13;
    wire [3:0] _T_986_14;
    wire [3:0] _T_986_15;
    wire [3:0] _T_986_16;
    wire [3:0] _T_986_17;
    wire [3:0] _T_986_18;
    wire [3:0] _T_986_19;
    wire [3:0] _T_986_20;
    wire [3:0] _T_986_21;
    wire [3:0] _T_986_22;
    wire [3:0] _T_986_23;
    wire [3:0] _T_986_24;
    wire [3:0] _T_986_25;
    wire [3:0] _T_986_26;
    wire [3:0] _T_986_27;
    wire [3:0] _T_986_28;
    wire [3:0] _T_986_29;
    wire [3:0] _T_986_30;
    wire [3:0] _T_986_31;
    wire [3:0] _T_986_32;
    wire [3:0] _T_986_33;
    wire [3:0] _T_986_34;
    wire [3:0] _T_986_35;
    wire [3:0] _T_986_36;
    wire [3:0] _T_986_37;
    wire [3:0] _T_986_38;
    wire [3:0] _T_986_39;
    wire [3:0] _T_986_40;
    wire [3:0] _T_986_41;
    wire [3:0] _T_986_42;
    wire [3:0] _T_986_43;
    wire [3:0] _T_986_44;
    wire [3:0] _T_986_45;
    wire [3:0] _T_986_46;
    wire [3:0] _T_986_47;
    wire [3:0] _T_986_48;
    wire [3:0] _T_986_49;
    wire [3:0] _T_986_50;
    wire [3:0] _T_986_51;
    wire [3:0] _T_986_52;
    wire [3:0] _T_986_53;
    wire [3:0] _T_986_54;
    wire [3:0] _T_986_55;
    wire [3:0] _T_986_56;
    wire [3:0] _T_986_57;
    wire [3:0] _T_986_58;
    wire [3:0] _T_986_59;
    wire [3:0] _T_986_60;
    wire [3:0] _T_986_61;
    wire [3:0] _T_986_62;
    wire [3:0] _T_986_63;
    wire [3:0] _T_986_64;
    wire [3:0] _T_986_65;
    wire [3:0] _T_986_66;
    wire [3:0] _T_986_67;
    wire [3:0] _T_986_68;
    wire [3:0] _T_986_69;
    wire [3:0] _T_986_70;
    wire [3:0] _T_986_71;
    wire [3:0] _T_986_72;
    wire [3:0] _T_986_73;
    wire [3:0] _T_986_74;
    wire [3:0] _T_986_75;
    wire [3:0] _T_986_76;
    wire [3:0] _T_986_77;
    wire [3:0] _T_986_78;
    wire [3:0] _T_986_79;
    wire [3:0] _T_986_80;
    wire [3:0] _T_986_81;
    wire [3:0] _T_986_82;
    wire [3:0] _T_986_83;
    wire [3:0] _T_986_84;
    wire [3:0] _T_986_85;
    wire [3:0] _T_986_86;
    wire [3:0] _T_986_87;
    wire [3:0] _T_986_88;
    wire [3:0] _T_986_89;
    wire [3:0] _T_986_90;
    wire [3:0] _T_986_91;
    wire [3:0] _T_986_92;
    wire [3:0] _T_986_93;
    wire [3:0] _T_986_94;
    wire [3:0] _T_986_95;
    wire [3:0] _T_986_96;
    wire [3:0] _T_986_97;
    wire [3:0] _T_986_98;
    wire [3:0] _T_986_99;
    wire [3:0] _T_986_100;
    wire [6:0] _T_1091;
    BITS #(.width(9), .high(6), .low(0)) bits_665 (
        .y(_T_1091),
        .in(__T_10__q)
    );
    wire _T_1094;
    EQ_UNSIGNED #(.width(1)) u_eq_666 (
        .y(_T_1094),
        .a(reset),
        .b(1'h0)
    );
    wire _node_618;
    EQ_UNSIGNED #(.width(7)) u_eq_667 (
        .y(_node_618),
        .a(7'd0),
        .b(_value_1__q)
    );
    wire [3:0] _node_619;
    assign _node_619 = _T_986_0;
    wire _node_620;
    EQ_UNSIGNED #(.width(7)) u_eq_668 (
        .y(_node_620),
        .a(7'd1),
        .b(_value_1__q)
    );
    wire [3:0] _node_621;
    MUX_UNSIGNED #(.width(4)) u_mux_669 (
        .y(_node_621),
        .sel(_node_620),
        .a(_T_986_1),
        .b(_node_619)
    );
    wire _node_622;
    EQ_UNSIGNED #(.width(7)) u_eq_670 (
        .y(_node_622),
        .a(7'd2),
        .b(_value_1__q)
    );
    wire [3:0] _node_623;
    MUX_UNSIGNED #(.width(4)) u_mux_671 (
        .y(_node_623),
        .sel(_node_622),
        .a(_T_986_2),
        .b(_node_621)
    );
    wire _node_624;
    EQ_UNSIGNED #(.width(7)) u_eq_672 (
        .y(_node_624),
        .a(7'd3),
        .b(_value_1__q)
    );
    wire [3:0] _node_625;
    MUX_UNSIGNED #(.width(4)) u_mux_673 (
        .y(_node_625),
        .sel(_node_624),
        .a(_T_986_3),
        .b(_node_623)
    );
    wire _node_626;
    EQ_UNSIGNED #(.width(7)) u_eq_674 (
        .y(_node_626),
        .a(7'd4),
        .b(_value_1__q)
    );
    wire [3:0] _node_627;
    MUX_UNSIGNED #(.width(4)) u_mux_675 (
        .y(_node_627),
        .sel(_node_626),
        .a(_T_986_4),
        .b(_node_625)
    );
    wire _node_628;
    EQ_UNSIGNED #(.width(7)) u_eq_676 (
        .y(_node_628),
        .a(7'd5),
        .b(_value_1__q)
    );
    wire [3:0] _node_629;
    MUX_UNSIGNED #(.width(4)) u_mux_677 (
        .y(_node_629),
        .sel(_node_628),
        .a(_T_986_5),
        .b(_node_627)
    );
    wire _node_630;
    EQ_UNSIGNED #(.width(7)) u_eq_678 (
        .y(_node_630),
        .a(7'd6),
        .b(_value_1__q)
    );
    wire [3:0] _node_631;
    MUX_UNSIGNED #(.width(4)) u_mux_679 (
        .y(_node_631),
        .sel(_node_630),
        .a(_T_986_6),
        .b(_node_629)
    );
    wire _node_632;
    EQ_UNSIGNED #(.width(7)) u_eq_680 (
        .y(_node_632),
        .a(7'd7),
        .b(_value_1__q)
    );
    wire [3:0] _node_633;
    MUX_UNSIGNED #(.width(4)) u_mux_681 (
        .y(_node_633),
        .sel(_node_632),
        .a(_T_986_7),
        .b(_node_631)
    );
    wire _node_634;
    EQ_UNSIGNED #(.width(7)) u_eq_682 (
        .y(_node_634),
        .a(7'd8),
        .b(_value_1__q)
    );
    wire [3:0] _node_635;
    MUX_UNSIGNED #(.width(4)) u_mux_683 (
        .y(_node_635),
        .sel(_node_634),
        .a(_T_986_8),
        .b(_node_633)
    );
    wire _node_636;
    EQ_UNSIGNED #(.width(7)) u_eq_684 (
        .y(_node_636),
        .a(7'd9),
        .b(_value_1__q)
    );
    wire [3:0] _node_637;
    MUX_UNSIGNED #(.width(4)) u_mux_685 (
        .y(_node_637),
        .sel(_node_636),
        .a(_T_986_9),
        .b(_node_635)
    );
    wire _node_638;
    EQ_UNSIGNED #(.width(7)) u_eq_686 (
        .y(_node_638),
        .a(7'd10),
        .b(_value_1__q)
    );
    wire [3:0] _node_639;
    MUX_UNSIGNED #(.width(4)) u_mux_687 (
        .y(_node_639),
        .sel(_node_638),
        .a(_T_986_10),
        .b(_node_637)
    );
    wire _node_640;
    EQ_UNSIGNED #(.width(7)) u_eq_688 (
        .y(_node_640),
        .a(7'd11),
        .b(_value_1__q)
    );
    wire [3:0] _node_641;
    MUX_UNSIGNED #(.width(4)) u_mux_689 (
        .y(_node_641),
        .sel(_node_640),
        .a(_T_986_11),
        .b(_node_639)
    );
    wire _node_642;
    EQ_UNSIGNED #(.width(7)) u_eq_690 (
        .y(_node_642),
        .a(7'd12),
        .b(_value_1__q)
    );
    wire [3:0] _node_643;
    MUX_UNSIGNED #(.width(4)) u_mux_691 (
        .y(_node_643),
        .sel(_node_642),
        .a(_T_986_12),
        .b(_node_641)
    );
    wire _node_644;
    EQ_UNSIGNED #(.width(7)) u_eq_692 (
        .y(_node_644),
        .a(7'd13),
        .b(_value_1__q)
    );
    wire [3:0] _node_645;
    MUX_UNSIGNED #(.width(4)) u_mux_693 (
        .y(_node_645),
        .sel(_node_644),
        .a(_T_986_13),
        .b(_node_643)
    );
    wire _node_646;
    EQ_UNSIGNED #(.width(7)) u_eq_694 (
        .y(_node_646),
        .a(7'd14),
        .b(_value_1__q)
    );
    wire [3:0] _node_647;
    MUX_UNSIGNED #(.width(4)) u_mux_695 (
        .y(_node_647),
        .sel(_node_646),
        .a(_T_986_14),
        .b(_node_645)
    );
    wire _node_648;
    EQ_UNSIGNED #(.width(7)) u_eq_696 (
        .y(_node_648),
        .a(7'd15),
        .b(_value_1__q)
    );
    wire [3:0] _node_649;
    MUX_UNSIGNED #(.width(4)) u_mux_697 (
        .y(_node_649),
        .sel(_node_648),
        .a(_T_986_15),
        .b(_node_647)
    );
    wire _node_650;
    EQ_UNSIGNED #(.width(7)) u_eq_698 (
        .y(_node_650),
        .a(7'd16),
        .b(_value_1__q)
    );
    wire [3:0] _node_651;
    MUX_UNSIGNED #(.width(4)) u_mux_699 (
        .y(_node_651),
        .sel(_node_650),
        .a(_T_986_16),
        .b(_node_649)
    );
    wire _node_652;
    EQ_UNSIGNED #(.width(7)) u_eq_700 (
        .y(_node_652),
        .a(7'd17),
        .b(_value_1__q)
    );
    wire [3:0] _node_653;
    MUX_UNSIGNED #(.width(4)) u_mux_701 (
        .y(_node_653),
        .sel(_node_652),
        .a(_T_986_17),
        .b(_node_651)
    );
    wire _node_654;
    EQ_UNSIGNED #(.width(7)) u_eq_702 (
        .y(_node_654),
        .a(7'd18),
        .b(_value_1__q)
    );
    wire [3:0] _node_655;
    MUX_UNSIGNED #(.width(4)) u_mux_703 (
        .y(_node_655),
        .sel(_node_654),
        .a(_T_986_18),
        .b(_node_653)
    );
    wire _node_656;
    EQ_UNSIGNED #(.width(7)) u_eq_704 (
        .y(_node_656),
        .a(7'd19),
        .b(_value_1__q)
    );
    wire [3:0] _node_657;
    MUX_UNSIGNED #(.width(4)) u_mux_705 (
        .y(_node_657),
        .sel(_node_656),
        .a(_T_986_19),
        .b(_node_655)
    );
    wire _node_658;
    EQ_UNSIGNED #(.width(7)) u_eq_706 (
        .y(_node_658),
        .a(7'd20),
        .b(_value_1__q)
    );
    wire [3:0] _node_659;
    MUX_UNSIGNED #(.width(4)) u_mux_707 (
        .y(_node_659),
        .sel(_node_658),
        .a(_T_986_20),
        .b(_node_657)
    );
    wire _node_660;
    EQ_UNSIGNED #(.width(7)) u_eq_708 (
        .y(_node_660),
        .a(7'd21),
        .b(_value_1__q)
    );
    wire [3:0] _node_661;
    MUX_UNSIGNED #(.width(4)) u_mux_709 (
        .y(_node_661),
        .sel(_node_660),
        .a(_T_986_21),
        .b(_node_659)
    );
    wire _node_662;
    EQ_UNSIGNED #(.width(7)) u_eq_710 (
        .y(_node_662),
        .a(7'd22),
        .b(_value_1__q)
    );
    wire [3:0] _node_663;
    MUX_UNSIGNED #(.width(4)) u_mux_711 (
        .y(_node_663),
        .sel(_node_662),
        .a(_T_986_22),
        .b(_node_661)
    );
    wire _node_664;
    EQ_UNSIGNED #(.width(7)) u_eq_712 (
        .y(_node_664),
        .a(7'd23),
        .b(_value_1__q)
    );
    wire [3:0] _node_665;
    MUX_UNSIGNED #(.width(4)) u_mux_713 (
        .y(_node_665),
        .sel(_node_664),
        .a(_T_986_23),
        .b(_node_663)
    );
    wire _node_666;
    EQ_UNSIGNED #(.width(7)) u_eq_714 (
        .y(_node_666),
        .a(7'd24),
        .b(_value_1__q)
    );
    wire [3:0] _node_667;
    MUX_UNSIGNED #(.width(4)) u_mux_715 (
        .y(_node_667),
        .sel(_node_666),
        .a(_T_986_24),
        .b(_node_665)
    );
    wire _node_668;
    EQ_UNSIGNED #(.width(7)) u_eq_716 (
        .y(_node_668),
        .a(7'd25),
        .b(_value_1__q)
    );
    wire [3:0] _node_669;
    MUX_UNSIGNED #(.width(4)) u_mux_717 (
        .y(_node_669),
        .sel(_node_668),
        .a(_T_986_25),
        .b(_node_667)
    );
    wire _node_670;
    EQ_UNSIGNED #(.width(7)) u_eq_718 (
        .y(_node_670),
        .a(7'd26),
        .b(_value_1__q)
    );
    wire [3:0] _node_671;
    MUX_UNSIGNED #(.width(4)) u_mux_719 (
        .y(_node_671),
        .sel(_node_670),
        .a(_T_986_26),
        .b(_node_669)
    );
    wire _node_672;
    EQ_UNSIGNED #(.width(7)) u_eq_720 (
        .y(_node_672),
        .a(7'd27),
        .b(_value_1__q)
    );
    wire [3:0] _node_673;
    MUX_UNSIGNED #(.width(4)) u_mux_721 (
        .y(_node_673),
        .sel(_node_672),
        .a(_T_986_27),
        .b(_node_671)
    );
    wire _node_674;
    EQ_UNSIGNED #(.width(7)) u_eq_722 (
        .y(_node_674),
        .a(7'd28),
        .b(_value_1__q)
    );
    wire [3:0] _node_675;
    MUX_UNSIGNED #(.width(4)) u_mux_723 (
        .y(_node_675),
        .sel(_node_674),
        .a(_T_986_28),
        .b(_node_673)
    );
    wire _node_676;
    EQ_UNSIGNED #(.width(7)) u_eq_724 (
        .y(_node_676),
        .a(7'd29),
        .b(_value_1__q)
    );
    wire [3:0] _node_677;
    MUX_UNSIGNED #(.width(4)) u_mux_725 (
        .y(_node_677),
        .sel(_node_676),
        .a(_T_986_29),
        .b(_node_675)
    );
    wire _node_678;
    EQ_UNSIGNED #(.width(7)) u_eq_726 (
        .y(_node_678),
        .a(7'd30),
        .b(_value_1__q)
    );
    wire [3:0] _node_679;
    MUX_UNSIGNED #(.width(4)) u_mux_727 (
        .y(_node_679),
        .sel(_node_678),
        .a(_T_986_30),
        .b(_node_677)
    );
    wire _node_680;
    EQ_UNSIGNED #(.width(7)) u_eq_728 (
        .y(_node_680),
        .a(7'd31),
        .b(_value_1__q)
    );
    wire [3:0] _node_681;
    MUX_UNSIGNED #(.width(4)) u_mux_729 (
        .y(_node_681),
        .sel(_node_680),
        .a(_T_986_31),
        .b(_node_679)
    );
    wire _node_682;
    EQ_UNSIGNED #(.width(7)) u_eq_730 (
        .y(_node_682),
        .a(7'd32),
        .b(_value_1__q)
    );
    wire [3:0] _node_683;
    MUX_UNSIGNED #(.width(4)) u_mux_731 (
        .y(_node_683),
        .sel(_node_682),
        .a(_T_986_32),
        .b(_node_681)
    );
    wire _node_684;
    EQ_UNSIGNED #(.width(7)) u_eq_732 (
        .y(_node_684),
        .a(7'd33),
        .b(_value_1__q)
    );
    wire [3:0] _node_685;
    MUX_UNSIGNED #(.width(4)) u_mux_733 (
        .y(_node_685),
        .sel(_node_684),
        .a(_T_986_33),
        .b(_node_683)
    );
    wire _node_686;
    EQ_UNSIGNED #(.width(7)) u_eq_734 (
        .y(_node_686),
        .a(7'd34),
        .b(_value_1__q)
    );
    wire [3:0] _node_687;
    MUX_UNSIGNED #(.width(4)) u_mux_735 (
        .y(_node_687),
        .sel(_node_686),
        .a(_T_986_34),
        .b(_node_685)
    );
    wire _node_688;
    EQ_UNSIGNED #(.width(7)) u_eq_736 (
        .y(_node_688),
        .a(7'd35),
        .b(_value_1__q)
    );
    wire [3:0] _node_689;
    MUX_UNSIGNED #(.width(4)) u_mux_737 (
        .y(_node_689),
        .sel(_node_688),
        .a(_T_986_35),
        .b(_node_687)
    );
    wire _node_690;
    EQ_UNSIGNED #(.width(7)) u_eq_738 (
        .y(_node_690),
        .a(7'd36),
        .b(_value_1__q)
    );
    wire [3:0] _node_691;
    MUX_UNSIGNED #(.width(4)) u_mux_739 (
        .y(_node_691),
        .sel(_node_690),
        .a(_T_986_36),
        .b(_node_689)
    );
    wire _node_692;
    EQ_UNSIGNED #(.width(7)) u_eq_740 (
        .y(_node_692),
        .a(7'd37),
        .b(_value_1__q)
    );
    wire [3:0] _node_693;
    MUX_UNSIGNED #(.width(4)) u_mux_741 (
        .y(_node_693),
        .sel(_node_692),
        .a(_T_986_37),
        .b(_node_691)
    );
    wire _node_694;
    EQ_UNSIGNED #(.width(7)) u_eq_742 (
        .y(_node_694),
        .a(7'd38),
        .b(_value_1__q)
    );
    wire [3:0] _node_695;
    MUX_UNSIGNED #(.width(4)) u_mux_743 (
        .y(_node_695),
        .sel(_node_694),
        .a(_T_986_38),
        .b(_node_693)
    );
    wire _node_696;
    EQ_UNSIGNED #(.width(7)) u_eq_744 (
        .y(_node_696),
        .a(7'd39),
        .b(_value_1__q)
    );
    wire [3:0] _node_697;
    MUX_UNSIGNED #(.width(4)) u_mux_745 (
        .y(_node_697),
        .sel(_node_696),
        .a(_T_986_39),
        .b(_node_695)
    );
    wire _node_698;
    EQ_UNSIGNED #(.width(7)) u_eq_746 (
        .y(_node_698),
        .a(7'd40),
        .b(_value_1__q)
    );
    wire [3:0] _node_699;
    MUX_UNSIGNED #(.width(4)) u_mux_747 (
        .y(_node_699),
        .sel(_node_698),
        .a(_T_986_40),
        .b(_node_697)
    );
    wire _node_700;
    EQ_UNSIGNED #(.width(7)) u_eq_748 (
        .y(_node_700),
        .a(7'd41),
        .b(_value_1__q)
    );
    wire [3:0] _node_701;
    MUX_UNSIGNED #(.width(4)) u_mux_749 (
        .y(_node_701),
        .sel(_node_700),
        .a(_T_986_41),
        .b(_node_699)
    );
    wire _node_702;
    EQ_UNSIGNED #(.width(7)) u_eq_750 (
        .y(_node_702),
        .a(7'd42),
        .b(_value_1__q)
    );
    wire [3:0] _node_703;
    MUX_UNSIGNED #(.width(4)) u_mux_751 (
        .y(_node_703),
        .sel(_node_702),
        .a(_T_986_42),
        .b(_node_701)
    );
    wire _node_704;
    EQ_UNSIGNED #(.width(7)) u_eq_752 (
        .y(_node_704),
        .a(7'd43),
        .b(_value_1__q)
    );
    wire [3:0] _node_705;
    MUX_UNSIGNED #(.width(4)) u_mux_753 (
        .y(_node_705),
        .sel(_node_704),
        .a(_T_986_43),
        .b(_node_703)
    );
    wire _node_706;
    EQ_UNSIGNED #(.width(7)) u_eq_754 (
        .y(_node_706),
        .a(7'd44),
        .b(_value_1__q)
    );
    wire [3:0] _node_707;
    MUX_UNSIGNED #(.width(4)) u_mux_755 (
        .y(_node_707),
        .sel(_node_706),
        .a(_T_986_44),
        .b(_node_705)
    );
    wire _node_708;
    EQ_UNSIGNED #(.width(7)) u_eq_756 (
        .y(_node_708),
        .a(7'd45),
        .b(_value_1__q)
    );
    wire [3:0] _node_709;
    MUX_UNSIGNED #(.width(4)) u_mux_757 (
        .y(_node_709),
        .sel(_node_708),
        .a(_T_986_45),
        .b(_node_707)
    );
    wire _node_710;
    EQ_UNSIGNED #(.width(7)) u_eq_758 (
        .y(_node_710),
        .a(7'd46),
        .b(_value_1__q)
    );
    wire [3:0] _node_711;
    MUX_UNSIGNED #(.width(4)) u_mux_759 (
        .y(_node_711),
        .sel(_node_710),
        .a(_T_986_46),
        .b(_node_709)
    );
    wire _node_712;
    EQ_UNSIGNED #(.width(7)) u_eq_760 (
        .y(_node_712),
        .a(7'd47),
        .b(_value_1__q)
    );
    wire [3:0] _node_713;
    MUX_UNSIGNED #(.width(4)) u_mux_761 (
        .y(_node_713),
        .sel(_node_712),
        .a(_T_986_47),
        .b(_node_711)
    );
    wire _node_714;
    EQ_UNSIGNED #(.width(7)) u_eq_762 (
        .y(_node_714),
        .a(7'd48),
        .b(_value_1__q)
    );
    wire [3:0] _node_715;
    MUX_UNSIGNED #(.width(4)) u_mux_763 (
        .y(_node_715),
        .sel(_node_714),
        .a(_T_986_48),
        .b(_node_713)
    );
    wire _node_716;
    EQ_UNSIGNED #(.width(7)) u_eq_764 (
        .y(_node_716),
        .a(7'd49),
        .b(_value_1__q)
    );
    wire [3:0] _node_717;
    MUX_UNSIGNED #(.width(4)) u_mux_765 (
        .y(_node_717),
        .sel(_node_716),
        .a(_T_986_49),
        .b(_node_715)
    );
    wire _node_718;
    EQ_UNSIGNED #(.width(7)) u_eq_766 (
        .y(_node_718),
        .a(7'd50),
        .b(_value_1__q)
    );
    wire [3:0] _node_719;
    MUX_UNSIGNED #(.width(4)) u_mux_767 (
        .y(_node_719),
        .sel(_node_718),
        .a(_T_986_50),
        .b(_node_717)
    );
    wire _node_720;
    EQ_UNSIGNED #(.width(7)) u_eq_768 (
        .y(_node_720),
        .a(7'd51),
        .b(_value_1__q)
    );
    wire [3:0] _node_721;
    MUX_UNSIGNED #(.width(4)) u_mux_769 (
        .y(_node_721),
        .sel(_node_720),
        .a(_T_986_51),
        .b(_node_719)
    );
    wire _node_722;
    EQ_UNSIGNED #(.width(7)) u_eq_770 (
        .y(_node_722),
        .a(7'd52),
        .b(_value_1__q)
    );
    wire [3:0] _node_723;
    MUX_UNSIGNED #(.width(4)) u_mux_771 (
        .y(_node_723),
        .sel(_node_722),
        .a(_T_986_52),
        .b(_node_721)
    );
    wire _node_724;
    EQ_UNSIGNED #(.width(7)) u_eq_772 (
        .y(_node_724),
        .a(7'd53),
        .b(_value_1__q)
    );
    wire [3:0] _node_725;
    MUX_UNSIGNED #(.width(4)) u_mux_773 (
        .y(_node_725),
        .sel(_node_724),
        .a(_T_986_53),
        .b(_node_723)
    );
    wire _node_726;
    EQ_UNSIGNED #(.width(7)) u_eq_774 (
        .y(_node_726),
        .a(7'd54),
        .b(_value_1__q)
    );
    wire [3:0] _node_727;
    MUX_UNSIGNED #(.width(4)) u_mux_775 (
        .y(_node_727),
        .sel(_node_726),
        .a(_T_986_54),
        .b(_node_725)
    );
    wire _node_728;
    EQ_UNSIGNED #(.width(7)) u_eq_776 (
        .y(_node_728),
        .a(7'd55),
        .b(_value_1__q)
    );
    wire [3:0] _node_729;
    MUX_UNSIGNED #(.width(4)) u_mux_777 (
        .y(_node_729),
        .sel(_node_728),
        .a(_T_986_55),
        .b(_node_727)
    );
    wire _node_730;
    EQ_UNSIGNED #(.width(7)) u_eq_778 (
        .y(_node_730),
        .a(7'd56),
        .b(_value_1__q)
    );
    wire [3:0] _node_731;
    MUX_UNSIGNED #(.width(4)) u_mux_779 (
        .y(_node_731),
        .sel(_node_730),
        .a(_T_986_56),
        .b(_node_729)
    );
    wire _node_732;
    EQ_UNSIGNED #(.width(7)) u_eq_780 (
        .y(_node_732),
        .a(7'd57),
        .b(_value_1__q)
    );
    wire [3:0] _node_733;
    MUX_UNSIGNED #(.width(4)) u_mux_781 (
        .y(_node_733),
        .sel(_node_732),
        .a(_T_986_57),
        .b(_node_731)
    );
    wire _node_734;
    EQ_UNSIGNED #(.width(7)) u_eq_782 (
        .y(_node_734),
        .a(7'd58),
        .b(_value_1__q)
    );
    wire [3:0] _node_735;
    MUX_UNSIGNED #(.width(4)) u_mux_783 (
        .y(_node_735),
        .sel(_node_734),
        .a(_T_986_58),
        .b(_node_733)
    );
    wire _node_736;
    EQ_UNSIGNED #(.width(7)) u_eq_784 (
        .y(_node_736),
        .a(7'd59),
        .b(_value_1__q)
    );
    wire [3:0] _node_737;
    MUX_UNSIGNED #(.width(4)) u_mux_785 (
        .y(_node_737),
        .sel(_node_736),
        .a(_T_986_59),
        .b(_node_735)
    );
    wire _node_738;
    EQ_UNSIGNED #(.width(7)) u_eq_786 (
        .y(_node_738),
        .a(7'd60),
        .b(_value_1__q)
    );
    wire [3:0] _node_739;
    MUX_UNSIGNED #(.width(4)) u_mux_787 (
        .y(_node_739),
        .sel(_node_738),
        .a(_T_986_60),
        .b(_node_737)
    );
    wire _node_740;
    EQ_UNSIGNED #(.width(7)) u_eq_788 (
        .y(_node_740),
        .a(7'd61),
        .b(_value_1__q)
    );
    wire [3:0] _node_741;
    MUX_UNSIGNED #(.width(4)) u_mux_789 (
        .y(_node_741),
        .sel(_node_740),
        .a(_T_986_61),
        .b(_node_739)
    );
    wire _node_742;
    EQ_UNSIGNED #(.width(7)) u_eq_790 (
        .y(_node_742),
        .a(7'd62),
        .b(_value_1__q)
    );
    wire [3:0] _node_743;
    MUX_UNSIGNED #(.width(4)) u_mux_791 (
        .y(_node_743),
        .sel(_node_742),
        .a(_T_986_62),
        .b(_node_741)
    );
    wire _node_744;
    EQ_UNSIGNED #(.width(7)) u_eq_792 (
        .y(_node_744),
        .a(7'd63),
        .b(_value_1__q)
    );
    wire [3:0] _node_745;
    MUX_UNSIGNED #(.width(4)) u_mux_793 (
        .y(_node_745),
        .sel(_node_744),
        .a(_T_986_63),
        .b(_node_743)
    );
    wire _node_746;
    EQ_UNSIGNED #(.width(7)) u_eq_794 (
        .y(_node_746),
        .a(7'd64),
        .b(_value_1__q)
    );
    wire [3:0] _node_747;
    MUX_UNSIGNED #(.width(4)) u_mux_795 (
        .y(_node_747),
        .sel(_node_746),
        .a(_T_986_64),
        .b(_node_745)
    );
    wire _node_748;
    EQ_UNSIGNED #(.width(7)) u_eq_796 (
        .y(_node_748),
        .a(7'd65),
        .b(_value_1__q)
    );
    wire [3:0] _node_749;
    MUX_UNSIGNED #(.width(4)) u_mux_797 (
        .y(_node_749),
        .sel(_node_748),
        .a(_T_986_65),
        .b(_node_747)
    );
    wire _node_750;
    EQ_UNSIGNED #(.width(7)) u_eq_798 (
        .y(_node_750),
        .a(7'd66),
        .b(_value_1__q)
    );
    wire [3:0] _node_751;
    MUX_UNSIGNED #(.width(4)) u_mux_799 (
        .y(_node_751),
        .sel(_node_750),
        .a(_T_986_66),
        .b(_node_749)
    );
    wire _node_752;
    EQ_UNSIGNED #(.width(7)) u_eq_800 (
        .y(_node_752),
        .a(7'd67),
        .b(_value_1__q)
    );
    wire [3:0] _node_753;
    MUX_UNSIGNED #(.width(4)) u_mux_801 (
        .y(_node_753),
        .sel(_node_752),
        .a(_T_986_67),
        .b(_node_751)
    );
    wire _node_754;
    EQ_UNSIGNED #(.width(7)) u_eq_802 (
        .y(_node_754),
        .a(7'd68),
        .b(_value_1__q)
    );
    wire [3:0] _node_755;
    MUX_UNSIGNED #(.width(4)) u_mux_803 (
        .y(_node_755),
        .sel(_node_754),
        .a(_T_986_68),
        .b(_node_753)
    );
    wire _node_756;
    EQ_UNSIGNED #(.width(7)) u_eq_804 (
        .y(_node_756),
        .a(7'd69),
        .b(_value_1__q)
    );
    wire [3:0] _node_757;
    MUX_UNSIGNED #(.width(4)) u_mux_805 (
        .y(_node_757),
        .sel(_node_756),
        .a(_T_986_69),
        .b(_node_755)
    );
    wire _node_758;
    EQ_UNSIGNED #(.width(7)) u_eq_806 (
        .y(_node_758),
        .a(7'd70),
        .b(_value_1__q)
    );
    wire [3:0] _node_759;
    MUX_UNSIGNED #(.width(4)) u_mux_807 (
        .y(_node_759),
        .sel(_node_758),
        .a(_T_986_70),
        .b(_node_757)
    );
    wire _node_760;
    EQ_UNSIGNED #(.width(7)) u_eq_808 (
        .y(_node_760),
        .a(7'd71),
        .b(_value_1__q)
    );
    wire [3:0] _node_761;
    MUX_UNSIGNED #(.width(4)) u_mux_809 (
        .y(_node_761),
        .sel(_node_760),
        .a(_T_986_71),
        .b(_node_759)
    );
    wire _node_762;
    EQ_UNSIGNED #(.width(7)) u_eq_810 (
        .y(_node_762),
        .a(7'd72),
        .b(_value_1__q)
    );
    wire [3:0] _node_763;
    MUX_UNSIGNED #(.width(4)) u_mux_811 (
        .y(_node_763),
        .sel(_node_762),
        .a(_T_986_72),
        .b(_node_761)
    );
    wire _node_764;
    EQ_UNSIGNED #(.width(7)) u_eq_812 (
        .y(_node_764),
        .a(7'd73),
        .b(_value_1__q)
    );
    wire [3:0] _node_765;
    MUX_UNSIGNED #(.width(4)) u_mux_813 (
        .y(_node_765),
        .sel(_node_764),
        .a(_T_986_73),
        .b(_node_763)
    );
    wire _node_766;
    EQ_UNSIGNED #(.width(7)) u_eq_814 (
        .y(_node_766),
        .a(7'd74),
        .b(_value_1__q)
    );
    wire [3:0] _node_767;
    MUX_UNSIGNED #(.width(4)) u_mux_815 (
        .y(_node_767),
        .sel(_node_766),
        .a(_T_986_74),
        .b(_node_765)
    );
    wire _node_768;
    EQ_UNSIGNED #(.width(7)) u_eq_816 (
        .y(_node_768),
        .a(7'd75),
        .b(_value_1__q)
    );
    wire [3:0] _node_769;
    MUX_UNSIGNED #(.width(4)) u_mux_817 (
        .y(_node_769),
        .sel(_node_768),
        .a(_T_986_75),
        .b(_node_767)
    );
    wire _node_770;
    EQ_UNSIGNED #(.width(7)) u_eq_818 (
        .y(_node_770),
        .a(7'd76),
        .b(_value_1__q)
    );
    wire [3:0] _node_771;
    MUX_UNSIGNED #(.width(4)) u_mux_819 (
        .y(_node_771),
        .sel(_node_770),
        .a(_T_986_76),
        .b(_node_769)
    );
    wire _node_772;
    EQ_UNSIGNED #(.width(7)) u_eq_820 (
        .y(_node_772),
        .a(7'd77),
        .b(_value_1__q)
    );
    wire [3:0] _node_773;
    MUX_UNSIGNED #(.width(4)) u_mux_821 (
        .y(_node_773),
        .sel(_node_772),
        .a(_T_986_77),
        .b(_node_771)
    );
    wire _node_774;
    EQ_UNSIGNED #(.width(7)) u_eq_822 (
        .y(_node_774),
        .a(7'd78),
        .b(_value_1__q)
    );
    wire [3:0] _node_775;
    MUX_UNSIGNED #(.width(4)) u_mux_823 (
        .y(_node_775),
        .sel(_node_774),
        .a(_T_986_78),
        .b(_node_773)
    );
    wire _node_776;
    EQ_UNSIGNED #(.width(7)) u_eq_824 (
        .y(_node_776),
        .a(7'd79),
        .b(_value_1__q)
    );
    wire [3:0] _node_777;
    MUX_UNSIGNED #(.width(4)) u_mux_825 (
        .y(_node_777),
        .sel(_node_776),
        .a(_T_986_79),
        .b(_node_775)
    );
    wire _node_778;
    EQ_UNSIGNED #(.width(7)) u_eq_826 (
        .y(_node_778),
        .a(7'd80),
        .b(_value_1__q)
    );
    wire [3:0] _node_779;
    MUX_UNSIGNED #(.width(4)) u_mux_827 (
        .y(_node_779),
        .sel(_node_778),
        .a(_T_986_80),
        .b(_node_777)
    );
    wire _node_780;
    EQ_UNSIGNED #(.width(7)) u_eq_828 (
        .y(_node_780),
        .a(7'd81),
        .b(_value_1__q)
    );
    wire [3:0] _node_781;
    MUX_UNSIGNED #(.width(4)) u_mux_829 (
        .y(_node_781),
        .sel(_node_780),
        .a(_T_986_81),
        .b(_node_779)
    );
    wire _node_782;
    EQ_UNSIGNED #(.width(7)) u_eq_830 (
        .y(_node_782),
        .a(7'd82),
        .b(_value_1__q)
    );
    wire [3:0] _node_783;
    MUX_UNSIGNED #(.width(4)) u_mux_831 (
        .y(_node_783),
        .sel(_node_782),
        .a(_T_986_82),
        .b(_node_781)
    );
    wire _node_784;
    EQ_UNSIGNED #(.width(7)) u_eq_832 (
        .y(_node_784),
        .a(7'd83),
        .b(_value_1__q)
    );
    wire [3:0] _node_785;
    MUX_UNSIGNED #(.width(4)) u_mux_833 (
        .y(_node_785),
        .sel(_node_784),
        .a(_T_986_83),
        .b(_node_783)
    );
    wire _node_786;
    EQ_UNSIGNED #(.width(7)) u_eq_834 (
        .y(_node_786),
        .a(7'd84),
        .b(_value_1__q)
    );
    wire [3:0] _node_787;
    MUX_UNSIGNED #(.width(4)) u_mux_835 (
        .y(_node_787),
        .sel(_node_786),
        .a(_T_986_84),
        .b(_node_785)
    );
    wire _node_788;
    EQ_UNSIGNED #(.width(7)) u_eq_836 (
        .y(_node_788),
        .a(7'd85),
        .b(_value_1__q)
    );
    wire [3:0] _node_789;
    MUX_UNSIGNED #(.width(4)) u_mux_837 (
        .y(_node_789),
        .sel(_node_788),
        .a(_T_986_85),
        .b(_node_787)
    );
    wire _node_790;
    EQ_UNSIGNED #(.width(7)) u_eq_838 (
        .y(_node_790),
        .a(7'd86),
        .b(_value_1__q)
    );
    wire [3:0] _node_791;
    MUX_UNSIGNED #(.width(4)) u_mux_839 (
        .y(_node_791),
        .sel(_node_790),
        .a(_T_986_86),
        .b(_node_789)
    );
    wire _node_792;
    EQ_UNSIGNED #(.width(7)) u_eq_840 (
        .y(_node_792),
        .a(7'd87),
        .b(_value_1__q)
    );
    wire [3:0] _node_793;
    MUX_UNSIGNED #(.width(4)) u_mux_841 (
        .y(_node_793),
        .sel(_node_792),
        .a(_T_986_87),
        .b(_node_791)
    );
    wire _node_794;
    EQ_UNSIGNED #(.width(7)) u_eq_842 (
        .y(_node_794),
        .a(7'd88),
        .b(_value_1__q)
    );
    wire [3:0] _node_795;
    MUX_UNSIGNED #(.width(4)) u_mux_843 (
        .y(_node_795),
        .sel(_node_794),
        .a(_T_986_88),
        .b(_node_793)
    );
    wire _node_796;
    EQ_UNSIGNED #(.width(7)) u_eq_844 (
        .y(_node_796),
        .a(7'd89),
        .b(_value_1__q)
    );
    wire [3:0] _node_797;
    MUX_UNSIGNED #(.width(4)) u_mux_845 (
        .y(_node_797),
        .sel(_node_796),
        .a(_T_986_89),
        .b(_node_795)
    );
    wire _node_798;
    EQ_UNSIGNED #(.width(7)) u_eq_846 (
        .y(_node_798),
        .a(7'd90),
        .b(_value_1__q)
    );
    wire [3:0] _node_799;
    MUX_UNSIGNED #(.width(4)) u_mux_847 (
        .y(_node_799),
        .sel(_node_798),
        .a(_T_986_90),
        .b(_node_797)
    );
    wire _node_800;
    EQ_UNSIGNED #(.width(7)) u_eq_848 (
        .y(_node_800),
        .a(7'd91),
        .b(_value_1__q)
    );
    wire [3:0] _node_801;
    MUX_UNSIGNED #(.width(4)) u_mux_849 (
        .y(_node_801),
        .sel(_node_800),
        .a(_T_986_91),
        .b(_node_799)
    );
    wire _node_802;
    EQ_UNSIGNED #(.width(7)) u_eq_850 (
        .y(_node_802),
        .a(7'd92),
        .b(_value_1__q)
    );
    wire [3:0] _node_803;
    MUX_UNSIGNED #(.width(4)) u_mux_851 (
        .y(_node_803),
        .sel(_node_802),
        .a(_T_986_92),
        .b(_node_801)
    );
    wire _node_804;
    EQ_UNSIGNED #(.width(7)) u_eq_852 (
        .y(_node_804),
        .a(7'd93),
        .b(_value_1__q)
    );
    wire [3:0] _node_805;
    MUX_UNSIGNED #(.width(4)) u_mux_853 (
        .y(_node_805),
        .sel(_node_804),
        .a(_T_986_93),
        .b(_node_803)
    );
    wire _node_806;
    EQ_UNSIGNED #(.width(7)) u_eq_854 (
        .y(_node_806),
        .a(7'd94),
        .b(_value_1__q)
    );
    wire [3:0] _node_807;
    MUX_UNSIGNED #(.width(4)) u_mux_855 (
        .y(_node_807),
        .sel(_node_806),
        .a(_T_986_94),
        .b(_node_805)
    );
    wire _node_808;
    EQ_UNSIGNED #(.width(7)) u_eq_856 (
        .y(_node_808),
        .a(7'd95),
        .b(_value_1__q)
    );
    wire [3:0] _node_809;
    MUX_UNSIGNED #(.width(4)) u_mux_857 (
        .y(_node_809),
        .sel(_node_808),
        .a(_T_986_95),
        .b(_node_807)
    );
    wire _node_810;
    EQ_UNSIGNED #(.width(7)) u_eq_858 (
        .y(_node_810),
        .a(7'd96),
        .b(_value_1__q)
    );
    wire [3:0] _node_811;
    MUX_UNSIGNED #(.width(4)) u_mux_859 (
        .y(_node_811),
        .sel(_node_810),
        .a(_T_986_96),
        .b(_node_809)
    );
    wire _node_812;
    EQ_UNSIGNED #(.width(7)) u_eq_860 (
        .y(_node_812),
        .a(7'd97),
        .b(_value_1__q)
    );
    wire [3:0] _node_813;
    MUX_UNSIGNED #(.width(4)) u_mux_861 (
        .y(_node_813),
        .sel(_node_812),
        .a(_T_986_97),
        .b(_node_811)
    );
    wire _node_814;
    EQ_UNSIGNED #(.width(7)) u_eq_862 (
        .y(_node_814),
        .a(7'd98),
        .b(_value_1__q)
    );
    wire [3:0] _node_815;
    MUX_UNSIGNED #(.width(4)) u_mux_863 (
        .y(_node_815),
        .sel(_node_814),
        .a(_T_986_98),
        .b(_node_813)
    );
    wire _node_816;
    EQ_UNSIGNED #(.width(7)) u_eq_864 (
        .y(_node_816),
        .a(7'd99),
        .b(_value_1__q)
    );
    wire [3:0] _node_817;
    MUX_UNSIGNED #(.width(4)) u_mux_865 (
        .y(_node_817),
        .sel(_node_816),
        .a(_T_986_99),
        .b(_node_815)
    );
    wire _node_818;
    EQ_UNSIGNED #(.width(7)) u_eq_866 (
        .y(_node_818),
        .a(7'd100),
        .b(_value_1__q)
    );
    wire [3:0] _node_819;
    MUX_UNSIGNED #(.width(4)) u_mux_867 (
        .y(_node_819),
        .sel(_node_818),
        .a(_T_986_100),
        .b(_node_817)
    );
    wire _T_1096;
    wire [15:0] _WTEMP_16;
    PAD_UNSIGNED #(.width(4), .n(16)) u_pad_868 (
        .y(_WTEMP_16),
        .in(_node_819)
    );
    NEQ_UNSIGNED #(.width(16)) u_neq_869 (
        .y(_T_1096),
        .a(_c__io_out_bits),
        .b(_WTEMP_16)
    );
    wire _T_1099;
    EQ_UNSIGNED #(.width(1)) u_eq_870 (
        .y(_T_1099),
        .a(reset),
        .b(1'h0)
    );
    wire _T_1101;
    BITWISEOR #(.width(1)) bitwiseor_871 (
        .y(_T_1101),
        .a(1'h0),
        .b(reset)
    );
    wire _T_1103;
    EQ_UNSIGNED #(.width(1)) u_eq_872 (
        .y(_T_1103),
        .a(_T_1101),
        .b(1'h0)
    );
    wire _T_1105;
    EQ_UNSIGNED #(.width(7)) u_eq_873 (
        .y(_T_1105),
        .a(_value_1__q),
        .b(7'h63)
    );
    wire [7:0] _T_1107;
    wire [6:0] _WTEMP_17;
    PAD_UNSIGNED #(.width(1), .n(7)) u_pad_874 (
        .y(_WTEMP_17),
        .in(1'h1)
    );
    ADD_UNSIGNED #(.width(7)) u_add_875 (
        .y(_T_1107),
        .a(_value_1__q),
        .b(_WTEMP_17)
    );
    wire [6:0] _T_1108;
    TAIL #(.width(8), .n(1)) tail_876 (
        .y(_T_1108),
        .in(_T_1107)
    );
    wire _T_1111;
    EQ_UNSIGNED #(.width(1)) u_eq_877 (
        .y(_T_1111),
        .a(__T_13__q),
        .b(1'h0)
    );
    wire _T_1113;
    wire [8:0] _WTEMP_18;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_878 (
        .y(_WTEMP_18),
        .in(7'h63)
    );
    EQ_UNSIGNED #(.width(9)) u_eq_879 (
        .y(_T_1113),
        .a(__T_10__q),
        .b(_WTEMP_18)
    );
    wire [9:0] _T_1116;
    wire [8:0] _WTEMP_19;
    PAD_UNSIGNED #(.width(1), .n(9)) u_pad_880 (
        .y(_WTEMP_19),
        .in(1'h1)
    );
    ADD_UNSIGNED #(.width(9)) u_add_881 (
        .y(_T_1116),
        .a(__T_10__q),
        .b(_WTEMP_19)
    );
    wire [8:0] _T_1117;
    TAIL #(.width(10), .n(1)) tail_882 (
        .y(_T_1117),
        .in(_T_1116)
    );
    wire _node_820;
    MUX_UNSIGNED #(.width(1)) u_mux_883 (
        .y(_node_820),
        .sel(_T_1113),
        .a(1'h1),
        .b(__T_13__q)
    );
    wire [8:0] _node_821;
    MUX_UNSIGNED #(.width(9)) u_mux_884 (
        .y(_node_821),
        .sel(_T_1111),
        .a(_T_1117),
        .b(__T_10__q)
    );
    wire _node_822;
    MUX_UNSIGNED #(.width(1)) u_mux_885 (
        .y(_node_822),
        .sel(_T_1111),
        .a(_node_820),
        .b(__T_13__q)
    );
    wire [6:0] _node_823;
    wire [6:0] _WTEMP_20;
    PAD_UNSIGNED #(.width(1), .n(7)) u_pad_886 (
        .y(_WTEMP_20),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(7)) u_mux_887 (
        .y(_node_823),
        .sel(_T_1105),
        .a(_WTEMP_20),
        .b(_T_1108)
    );
    wire _node_824;
    EQ_UNSIGNED #(.width(7)) u_eq_888 (
        .y(_node_824),
        .a(7'd0),
        .b(_T_1091)
    );
    wire _node_825;
    assign _node_825 = _T_777_0;
    wire _node_826;
    EQ_UNSIGNED #(.width(7)) u_eq_889 (
        .y(_node_826),
        .a(7'd1),
        .b(_T_1091)
    );
    wire _node_827;
    MUX_UNSIGNED #(.width(1)) u_mux_890 (
        .y(_node_827),
        .sel(_node_826),
        .a(_T_777_1),
        .b(_node_825)
    );
    wire _node_828;
    EQ_UNSIGNED #(.width(7)) u_eq_891 (
        .y(_node_828),
        .a(7'd2),
        .b(_T_1091)
    );
    wire _node_829;
    MUX_UNSIGNED #(.width(1)) u_mux_892 (
        .y(_node_829),
        .sel(_node_828),
        .a(_T_777_2),
        .b(_node_827)
    );
    wire _node_830;
    EQ_UNSIGNED #(.width(7)) u_eq_893 (
        .y(_node_830),
        .a(7'd3),
        .b(_T_1091)
    );
    wire _node_831;
    MUX_UNSIGNED #(.width(1)) u_mux_894 (
        .y(_node_831),
        .sel(_node_830),
        .a(_T_777_3),
        .b(_node_829)
    );
    wire _node_832;
    EQ_UNSIGNED #(.width(7)) u_eq_895 (
        .y(_node_832),
        .a(7'd4),
        .b(_T_1091)
    );
    wire _node_833;
    MUX_UNSIGNED #(.width(1)) u_mux_896 (
        .y(_node_833),
        .sel(_node_832),
        .a(_T_777_4),
        .b(_node_831)
    );
    wire _node_834;
    EQ_UNSIGNED #(.width(7)) u_eq_897 (
        .y(_node_834),
        .a(7'd5),
        .b(_T_1091)
    );
    wire _node_835;
    MUX_UNSIGNED #(.width(1)) u_mux_898 (
        .y(_node_835),
        .sel(_node_834),
        .a(_T_777_5),
        .b(_node_833)
    );
    wire _node_836;
    EQ_UNSIGNED #(.width(7)) u_eq_899 (
        .y(_node_836),
        .a(7'd6),
        .b(_T_1091)
    );
    wire _node_837;
    MUX_UNSIGNED #(.width(1)) u_mux_900 (
        .y(_node_837),
        .sel(_node_836),
        .a(_T_777_6),
        .b(_node_835)
    );
    wire _node_838;
    EQ_UNSIGNED #(.width(7)) u_eq_901 (
        .y(_node_838),
        .a(7'd7),
        .b(_T_1091)
    );
    wire _node_839;
    MUX_UNSIGNED #(.width(1)) u_mux_902 (
        .y(_node_839),
        .sel(_node_838),
        .a(_T_777_7),
        .b(_node_837)
    );
    wire _node_840;
    EQ_UNSIGNED #(.width(7)) u_eq_903 (
        .y(_node_840),
        .a(7'd8),
        .b(_T_1091)
    );
    wire _node_841;
    MUX_UNSIGNED #(.width(1)) u_mux_904 (
        .y(_node_841),
        .sel(_node_840),
        .a(_T_777_8),
        .b(_node_839)
    );
    wire _node_842;
    EQ_UNSIGNED #(.width(7)) u_eq_905 (
        .y(_node_842),
        .a(7'd9),
        .b(_T_1091)
    );
    wire _node_843;
    MUX_UNSIGNED #(.width(1)) u_mux_906 (
        .y(_node_843),
        .sel(_node_842),
        .a(_T_777_9),
        .b(_node_841)
    );
    wire _node_844;
    EQ_UNSIGNED #(.width(7)) u_eq_907 (
        .y(_node_844),
        .a(7'd10),
        .b(_T_1091)
    );
    wire _node_845;
    MUX_UNSIGNED #(.width(1)) u_mux_908 (
        .y(_node_845),
        .sel(_node_844),
        .a(_T_777_10),
        .b(_node_843)
    );
    wire _node_846;
    EQ_UNSIGNED #(.width(7)) u_eq_909 (
        .y(_node_846),
        .a(7'd11),
        .b(_T_1091)
    );
    wire _node_847;
    MUX_UNSIGNED #(.width(1)) u_mux_910 (
        .y(_node_847),
        .sel(_node_846),
        .a(_T_777_11),
        .b(_node_845)
    );
    wire _node_848;
    EQ_UNSIGNED #(.width(7)) u_eq_911 (
        .y(_node_848),
        .a(7'd12),
        .b(_T_1091)
    );
    wire _node_849;
    MUX_UNSIGNED #(.width(1)) u_mux_912 (
        .y(_node_849),
        .sel(_node_848),
        .a(_T_777_12),
        .b(_node_847)
    );
    wire _node_850;
    EQ_UNSIGNED #(.width(7)) u_eq_913 (
        .y(_node_850),
        .a(7'd13),
        .b(_T_1091)
    );
    wire _node_851;
    MUX_UNSIGNED #(.width(1)) u_mux_914 (
        .y(_node_851),
        .sel(_node_850),
        .a(_T_777_13),
        .b(_node_849)
    );
    wire _node_852;
    EQ_UNSIGNED #(.width(7)) u_eq_915 (
        .y(_node_852),
        .a(7'd14),
        .b(_T_1091)
    );
    wire _node_853;
    MUX_UNSIGNED #(.width(1)) u_mux_916 (
        .y(_node_853),
        .sel(_node_852),
        .a(_T_777_14),
        .b(_node_851)
    );
    wire _node_854;
    EQ_UNSIGNED #(.width(7)) u_eq_917 (
        .y(_node_854),
        .a(7'd15),
        .b(_T_1091)
    );
    wire _node_855;
    MUX_UNSIGNED #(.width(1)) u_mux_918 (
        .y(_node_855),
        .sel(_node_854),
        .a(_T_777_15),
        .b(_node_853)
    );
    wire _node_856;
    EQ_UNSIGNED #(.width(7)) u_eq_919 (
        .y(_node_856),
        .a(7'd16),
        .b(_T_1091)
    );
    wire _node_857;
    MUX_UNSIGNED #(.width(1)) u_mux_920 (
        .y(_node_857),
        .sel(_node_856),
        .a(_T_777_16),
        .b(_node_855)
    );
    wire _node_858;
    EQ_UNSIGNED #(.width(7)) u_eq_921 (
        .y(_node_858),
        .a(7'd17),
        .b(_T_1091)
    );
    wire _node_859;
    MUX_UNSIGNED #(.width(1)) u_mux_922 (
        .y(_node_859),
        .sel(_node_858),
        .a(_T_777_17),
        .b(_node_857)
    );
    wire _node_860;
    EQ_UNSIGNED #(.width(7)) u_eq_923 (
        .y(_node_860),
        .a(7'd18),
        .b(_T_1091)
    );
    wire _node_861;
    MUX_UNSIGNED #(.width(1)) u_mux_924 (
        .y(_node_861),
        .sel(_node_860),
        .a(_T_777_18),
        .b(_node_859)
    );
    wire _node_862;
    EQ_UNSIGNED #(.width(7)) u_eq_925 (
        .y(_node_862),
        .a(7'd19),
        .b(_T_1091)
    );
    wire _node_863;
    MUX_UNSIGNED #(.width(1)) u_mux_926 (
        .y(_node_863),
        .sel(_node_862),
        .a(_T_777_19),
        .b(_node_861)
    );
    wire _node_864;
    EQ_UNSIGNED #(.width(7)) u_eq_927 (
        .y(_node_864),
        .a(7'd20),
        .b(_T_1091)
    );
    wire _node_865;
    MUX_UNSIGNED #(.width(1)) u_mux_928 (
        .y(_node_865),
        .sel(_node_864),
        .a(_T_777_20),
        .b(_node_863)
    );
    wire _node_866;
    EQ_UNSIGNED #(.width(7)) u_eq_929 (
        .y(_node_866),
        .a(7'd21),
        .b(_T_1091)
    );
    wire _node_867;
    MUX_UNSIGNED #(.width(1)) u_mux_930 (
        .y(_node_867),
        .sel(_node_866),
        .a(_T_777_21),
        .b(_node_865)
    );
    wire _node_868;
    EQ_UNSIGNED #(.width(7)) u_eq_931 (
        .y(_node_868),
        .a(7'd22),
        .b(_T_1091)
    );
    wire _node_869;
    MUX_UNSIGNED #(.width(1)) u_mux_932 (
        .y(_node_869),
        .sel(_node_868),
        .a(_T_777_22),
        .b(_node_867)
    );
    wire _node_870;
    EQ_UNSIGNED #(.width(7)) u_eq_933 (
        .y(_node_870),
        .a(7'd23),
        .b(_T_1091)
    );
    wire _node_871;
    MUX_UNSIGNED #(.width(1)) u_mux_934 (
        .y(_node_871),
        .sel(_node_870),
        .a(_T_777_23),
        .b(_node_869)
    );
    wire _node_872;
    EQ_UNSIGNED #(.width(7)) u_eq_935 (
        .y(_node_872),
        .a(7'd24),
        .b(_T_1091)
    );
    wire _node_873;
    MUX_UNSIGNED #(.width(1)) u_mux_936 (
        .y(_node_873),
        .sel(_node_872),
        .a(_T_777_24),
        .b(_node_871)
    );
    wire _node_874;
    EQ_UNSIGNED #(.width(7)) u_eq_937 (
        .y(_node_874),
        .a(7'd25),
        .b(_T_1091)
    );
    wire _node_875;
    MUX_UNSIGNED #(.width(1)) u_mux_938 (
        .y(_node_875),
        .sel(_node_874),
        .a(_T_777_25),
        .b(_node_873)
    );
    wire _node_876;
    EQ_UNSIGNED #(.width(7)) u_eq_939 (
        .y(_node_876),
        .a(7'd26),
        .b(_T_1091)
    );
    wire _node_877;
    MUX_UNSIGNED #(.width(1)) u_mux_940 (
        .y(_node_877),
        .sel(_node_876),
        .a(_T_777_26),
        .b(_node_875)
    );
    wire _node_878;
    EQ_UNSIGNED #(.width(7)) u_eq_941 (
        .y(_node_878),
        .a(7'd27),
        .b(_T_1091)
    );
    wire _node_879;
    MUX_UNSIGNED #(.width(1)) u_mux_942 (
        .y(_node_879),
        .sel(_node_878),
        .a(_T_777_27),
        .b(_node_877)
    );
    wire _node_880;
    EQ_UNSIGNED #(.width(7)) u_eq_943 (
        .y(_node_880),
        .a(7'd28),
        .b(_T_1091)
    );
    wire _node_881;
    MUX_UNSIGNED #(.width(1)) u_mux_944 (
        .y(_node_881),
        .sel(_node_880),
        .a(_T_777_28),
        .b(_node_879)
    );
    wire _node_882;
    EQ_UNSIGNED #(.width(7)) u_eq_945 (
        .y(_node_882),
        .a(7'd29),
        .b(_T_1091)
    );
    wire _node_883;
    MUX_UNSIGNED #(.width(1)) u_mux_946 (
        .y(_node_883),
        .sel(_node_882),
        .a(_T_777_29),
        .b(_node_881)
    );
    wire _node_884;
    EQ_UNSIGNED #(.width(7)) u_eq_947 (
        .y(_node_884),
        .a(7'd30),
        .b(_T_1091)
    );
    wire _node_885;
    MUX_UNSIGNED #(.width(1)) u_mux_948 (
        .y(_node_885),
        .sel(_node_884),
        .a(_T_777_30),
        .b(_node_883)
    );
    wire _node_886;
    EQ_UNSIGNED #(.width(7)) u_eq_949 (
        .y(_node_886),
        .a(7'd31),
        .b(_T_1091)
    );
    wire _node_887;
    MUX_UNSIGNED #(.width(1)) u_mux_950 (
        .y(_node_887),
        .sel(_node_886),
        .a(_T_777_31),
        .b(_node_885)
    );
    wire _node_888;
    EQ_UNSIGNED #(.width(7)) u_eq_951 (
        .y(_node_888),
        .a(7'd32),
        .b(_T_1091)
    );
    wire _node_889;
    MUX_UNSIGNED #(.width(1)) u_mux_952 (
        .y(_node_889),
        .sel(_node_888),
        .a(_T_777_32),
        .b(_node_887)
    );
    wire _node_890;
    EQ_UNSIGNED #(.width(7)) u_eq_953 (
        .y(_node_890),
        .a(7'd33),
        .b(_T_1091)
    );
    wire _node_891;
    MUX_UNSIGNED #(.width(1)) u_mux_954 (
        .y(_node_891),
        .sel(_node_890),
        .a(_T_777_33),
        .b(_node_889)
    );
    wire _node_892;
    EQ_UNSIGNED #(.width(7)) u_eq_955 (
        .y(_node_892),
        .a(7'd34),
        .b(_T_1091)
    );
    wire _node_893;
    MUX_UNSIGNED #(.width(1)) u_mux_956 (
        .y(_node_893),
        .sel(_node_892),
        .a(_T_777_34),
        .b(_node_891)
    );
    wire _node_894;
    EQ_UNSIGNED #(.width(7)) u_eq_957 (
        .y(_node_894),
        .a(7'd35),
        .b(_T_1091)
    );
    wire _node_895;
    MUX_UNSIGNED #(.width(1)) u_mux_958 (
        .y(_node_895),
        .sel(_node_894),
        .a(_T_777_35),
        .b(_node_893)
    );
    wire _node_896;
    EQ_UNSIGNED #(.width(7)) u_eq_959 (
        .y(_node_896),
        .a(7'd36),
        .b(_T_1091)
    );
    wire _node_897;
    MUX_UNSIGNED #(.width(1)) u_mux_960 (
        .y(_node_897),
        .sel(_node_896),
        .a(_T_777_36),
        .b(_node_895)
    );
    wire _node_898;
    EQ_UNSIGNED #(.width(7)) u_eq_961 (
        .y(_node_898),
        .a(7'd37),
        .b(_T_1091)
    );
    wire _node_899;
    MUX_UNSIGNED #(.width(1)) u_mux_962 (
        .y(_node_899),
        .sel(_node_898),
        .a(_T_777_37),
        .b(_node_897)
    );
    wire _node_900;
    EQ_UNSIGNED #(.width(7)) u_eq_963 (
        .y(_node_900),
        .a(7'd38),
        .b(_T_1091)
    );
    wire _node_901;
    MUX_UNSIGNED #(.width(1)) u_mux_964 (
        .y(_node_901),
        .sel(_node_900),
        .a(_T_777_38),
        .b(_node_899)
    );
    wire _node_902;
    EQ_UNSIGNED #(.width(7)) u_eq_965 (
        .y(_node_902),
        .a(7'd39),
        .b(_T_1091)
    );
    wire _node_903;
    MUX_UNSIGNED #(.width(1)) u_mux_966 (
        .y(_node_903),
        .sel(_node_902),
        .a(_T_777_39),
        .b(_node_901)
    );
    wire _node_904;
    EQ_UNSIGNED #(.width(7)) u_eq_967 (
        .y(_node_904),
        .a(7'd40),
        .b(_T_1091)
    );
    wire _node_905;
    MUX_UNSIGNED #(.width(1)) u_mux_968 (
        .y(_node_905),
        .sel(_node_904),
        .a(_T_777_40),
        .b(_node_903)
    );
    wire _node_906;
    EQ_UNSIGNED #(.width(7)) u_eq_969 (
        .y(_node_906),
        .a(7'd41),
        .b(_T_1091)
    );
    wire _node_907;
    MUX_UNSIGNED #(.width(1)) u_mux_970 (
        .y(_node_907),
        .sel(_node_906),
        .a(_T_777_41),
        .b(_node_905)
    );
    wire _node_908;
    EQ_UNSIGNED #(.width(7)) u_eq_971 (
        .y(_node_908),
        .a(7'd42),
        .b(_T_1091)
    );
    wire _node_909;
    MUX_UNSIGNED #(.width(1)) u_mux_972 (
        .y(_node_909),
        .sel(_node_908),
        .a(_T_777_42),
        .b(_node_907)
    );
    wire _node_910;
    EQ_UNSIGNED #(.width(7)) u_eq_973 (
        .y(_node_910),
        .a(7'd43),
        .b(_T_1091)
    );
    wire _node_911;
    MUX_UNSIGNED #(.width(1)) u_mux_974 (
        .y(_node_911),
        .sel(_node_910),
        .a(_T_777_43),
        .b(_node_909)
    );
    wire _node_912;
    EQ_UNSIGNED #(.width(7)) u_eq_975 (
        .y(_node_912),
        .a(7'd44),
        .b(_T_1091)
    );
    wire _node_913;
    MUX_UNSIGNED #(.width(1)) u_mux_976 (
        .y(_node_913),
        .sel(_node_912),
        .a(_T_777_44),
        .b(_node_911)
    );
    wire _node_914;
    EQ_UNSIGNED #(.width(7)) u_eq_977 (
        .y(_node_914),
        .a(7'd45),
        .b(_T_1091)
    );
    wire _node_915;
    MUX_UNSIGNED #(.width(1)) u_mux_978 (
        .y(_node_915),
        .sel(_node_914),
        .a(_T_777_45),
        .b(_node_913)
    );
    wire _node_916;
    EQ_UNSIGNED #(.width(7)) u_eq_979 (
        .y(_node_916),
        .a(7'd46),
        .b(_T_1091)
    );
    wire _node_917;
    MUX_UNSIGNED #(.width(1)) u_mux_980 (
        .y(_node_917),
        .sel(_node_916),
        .a(_T_777_46),
        .b(_node_915)
    );
    wire _node_918;
    EQ_UNSIGNED #(.width(7)) u_eq_981 (
        .y(_node_918),
        .a(7'd47),
        .b(_T_1091)
    );
    wire _node_919;
    MUX_UNSIGNED #(.width(1)) u_mux_982 (
        .y(_node_919),
        .sel(_node_918),
        .a(_T_777_47),
        .b(_node_917)
    );
    wire _node_920;
    EQ_UNSIGNED #(.width(7)) u_eq_983 (
        .y(_node_920),
        .a(7'd48),
        .b(_T_1091)
    );
    wire _node_921;
    MUX_UNSIGNED #(.width(1)) u_mux_984 (
        .y(_node_921),
        .sel(_node_920),
        .a(_T_777_48),
        .b(_node_919)
    );
    wire _node_922;
    EQ_UNSIGNED #(.width(7)) u_eq_985 (
        .y(_node_922),
        .a(7'd49),
        .b(_T_1091)
    );
    wire _node_923;
    MUX_UNSIGNED #(.width(1)) u_mux_986 (
        .y(_node_923),
        .sel(_node_922),
        .a(_T_777_49),
        .b(_node_921)
    );
    wire _node_924;
    EQ_UNSIGNED #(.width(7)) u_eq_987 (
        .y(_node_924),
        .a(7'd50),
        .b(_T_1091)
    );
    wire _node_925;
    MUX_UNSIGNED #(.width(1)) u_mux_988 (
        .y(_node_925),
        .sel(_node_924),
        .a(_T_777_50),
        .b(_node_923)
    );
    wire _node_926;
    EQ_UNSIGNED #(.width(7)) u_eq_989 (
        .y(_node_926),
        .a(7'd51),
        .b(_T_1091)
    );
    wire _node_927;
    MUX_UNSIGNED #(.width(1)) u_mux_990 (
        .y(_node_927),
        .sel(_node_926),
        .a(_T_777_51),
        .b(_node_925)
    );
    wire _node_928;
    EQ_UNSIGNED #(.width(7)) u_eq_991 (
        .y(_node_928),
        .a(7'd52),
        .b(_T_1091)
    );
    wire _node_929;
    MUX_UNSIGNED #(.width(1)) u_mux_992 (
        .y(_node_929),
        .sel(_node_928),
        .a(_T_777_52),
        .b(_node_927)
    );
    wire _node_930;
    EQ_UNSIGNED #(.width(7)) u_eq_993 (
        .y(_node_930),
        .a(7'd53),
        .b(_T_1091)
    );
    wire _node_931;
    MUX_UNSIGNED #(.width(1)) u_mux_994 (
        .y(_node_931),
        .sel(_node_930),
        .a(_T_777_53),
        .b(_node_929)
    );
    wire _node_932;
    EQ_UNSIGNED #(.width(7)) u_eq_995 (
        .y(_node_932),
        .a(7'd54),
        .b(_T_1091)
    );
    wire _node_933;
    MUX_UNSIGNED #(.width(1)) u_mux_996 (
        .y(_node_933),
        .sel(_node_932),
        .a(_T_777_54),
        .b(_node_931)
    );
    wire _node_934;
    EQ_UNSIGNED #(.width(7)) u_eq_997 (
        .y(_node_934),
        .a(7'd55),
        .b(_T_1091)
    );
    wire _node_935;
    MUX_UNSIGNED #(.width(1)) u_mux_998 (
        .y(_node_935),
        .sel(_node_934),
        .a(_T_777_55),
        .b(_node_933)
    );
    wire _node_936;
    EQ_UNSIGNED #(.width(7)) u_eq_999 (
        .y(_node_936),
        .a(7'd56),
        .b(_T_1091)
    );
    wire _node_937;
    MUX_UNSIGNED #(.width(1)) u_mux_1000 (
        .y(_node_937),
        .sel(_node_936),
        .a(_T_777_56),
        .b(_node_935)
    );
    wire _node_938;
    EQ_UNSIGNED #(.width(7)) u_eq_1001 (
        .y(_node_938),
        .a(7'd57),
        .b(_T_1091)
    );
    wire _node_939;
    MUX_UNSIGNED #(.width(1)) u_mux_1002 (
        .y(_node_939),
        .sel(_node_938),
        .a(_T_777_57),
        .b(_node_937)
    );
    wire _node_940;
    EQ_UNSIGNED #(.width(7)) u_eq_1003 (
        .y(_node_940),
        .a(7'd58),
        .b(_T_1091)
    );
    wire _node_941;
    MUX_UNSIGNED #(.width(1)) u_mux_1004 (
        .y(_node_941),
        .sel(_node_940),
        .a(_T_777_58),
        .b(_node_939)
    );
    wire _node_942;
    EQ_UNSIGNED #(.width(7)) u_eq_1005 (
        .y(_node_942),
        .a(7'd59),
        .b(_T_1091)
    );
    wire _node_943;
    MUX_UNSIGNED #(.width(1)) u_mux_1006 (
        .y(_node_943),
        .sel(_node_942),
        .a(_T_777_59),
        .b(_node_941)
    );
    wire _node_944;
    EQ_UNSIGNED #(.width(7)) u_eq_1007 (
        .y(_node_944),
        .a(7'd60),
        .b(_T_1091)
    );
    wire _node_945;
    MUX_UNSIGNED #(.width(1)) u_mux_1008 (
        .y(_node_945),
        .sel(_node_944),
        .a(_T_777_60),
        .b(_node_943)
    );
    wire _node_946;
    EQ_UNSIGNED #(.width(7)) u_eq_1009 (
        .y(_node_946),
        .a(7'd61),
        .b(_T_1091)
    );
    wire _node_947;
    MUX_UNSIGNED #(.width(1)) u_mux_1010 (
        .y(_node_947),
        .sel(_node_946),
        .a(_T_777_61),
        .b(_node_945)
    );
    wire _node_948;
    EQ_UNSIGNED #(.width(7)) u_eq_1011 (
        .y(_node_948),
        .a(7'd62),
        .b(_T_1091)
    );
    wire _node_949;
    MUX_UNSIGNED #(.width(1)) u_mux_1012 (
        .y(_node_949),
        .sel(_node_948),
        .a(_T_777_62),
        .b(_node_947)
    );
    wire _node_950;
    EQ_UNSIGNED #(.width(7)) u_eq_1013 (
        .y(_node_950),
        .a(7'd63),
        .b(_T_1091)
    );
    wire _node_951;
    MUX_UNSIGNED #(.width(1)) u_mux_1014 (
        .y(_node_951),
        .sel(_node_950),
        .a(_T_777_63),
        .b(_node_949)
    );
    wire _node_952;
    EQ_UNSIGNED #(.width(7)) u_eq_1015 (
        .y(_node_952),
        .a(7'd64),
        .b(_T_1091)
    );
    wire _node_953;
    MUX_UNSIGNED #(.width(1)) u_mux_1016 (
        .y(_node_953),
        .sel(_node_952),
        .a(_T_777_64),
        .b(_node_951)
    );
    wire _node_954;
    EQ_UNSIGNED #(.width(7)) u_eq_1017 (
        .y(_node_954),
        .a(7'd65),
        .b(_T_1091)
    );
    wire _node_955;
    MUX_UNSIGNED #(.width(1)) u_mux_1018 (
        .y(_node_955),
        .sel(_node_954),
        .a(_T_777_65),
        .b(_node_953)
    );
    wire _node_956;
    EQ_UNSIGNED #(.width(7)) u_eq_1019 (
        .y(_node_956),
        .a(7'd66),
        .b(_T_1091)
    );
    wire _node_957;
    MUX_UNSIGNED #(.width(1)) u_mux_1020 (
        .y(_node_957),
        .sel(_node_956),
        .a(_T_777_66),
        .b(_node_955)
    );
    wire _node_958;
    EQ_UNSIGNED #(.width(7)) u_eq_1021 (
        .y(_node_958),
        .a(7'd67),
        .b(_T_1091)
    );
    wire _node_959;
    MUX_UNSIGNED #(.width(1)) u_mux_1022 (
        .y(_node_959),
        .sel(_node_958),
        .a(_T_777_67),
        .b(_node_957)
    );
    wire _node_960;
    EQ_UNSIGNED #(.width(7)) u_eq_1023 (
        .y(_node_960),
        .a(7'd68),
        .b(_T_1091)
    );
    wire _node_961;
    MUX_UNSIGNED #(.width(1)) u_mux_1024 (
        .y(_node_961),
        .sel(_node_960),
        .a(_T_777_68),
        .b(_node_959)
    );
    wire _node_962;
    EQ_UNSIGNED #(.width(7)) u_eq_1025 (
        .y(_node_962),
        .a(7'd69),
        .b(_T_1091)
    );
    wire _node_963;
    MUX_UNSIGNED #(.width(1)) u_mux_1026 (
        .y(_node_963),
        .sel(_node_962),
        .a(_T_777_69),
        .b(_node_961)
    );
    wire _node_964;
    EQ_UNSIGNED #(.width(7)) u_eq_1027 (
        .y(_node_964),
        .a(7'd70),
        .b(_T_1091)
    );
    wire _node_965;
    MUX_UNSIGNED #(.width(1)) u_mux_1028 (
        .y(_node_965),
        .sel(_node_964),
        .a(_T_777_70),
        .b(_node_963)
    );
    wire _node_966;
    EQ_UNSIGNED #(.width(7)) u_eq_1029 (
        .y(_node_966),
        .a(7'd71),
        .b(_T_1091)
    );
    wire _node_967;
    MUX_UNSIGNED #(.width(1)) u_mux_1030 (
        .y(_node_967),
        .sel(_node_966),
        .a(_T_777_71),
        .b(_node_965)
    );
    wire _node_968;
    EQ_UNSIGNED #(.width(7)) u_eq_1031 (
        .y(_node_968),
        .a(7'd72),
        .b(_T_1091)
    );
    wire _node_969;
    MUX_UNSIGNED #(.width(1)) u_mux_1032 (
        .y(_node_969),
        .sel(_node_968),
        .a(_T_777_72),
        .b(_node_967)
    );
    wire _node_970;
    EQ_UNSIGNED #(.width(7)) u_eq_1033 (
        .y(_node_970),
        .a(7'd73),
        .b(_T_1091)
    );
    wire _node_971;
    MUX_UNSIGNED #(.width(1)) u_mux_1034 (
        .y(_node_971),
        .sel(_node_970),
        .a(_T_777_73),
        .b(_node_969)
    );
    wire _node_972;
    EQ_UNSIGNED #(.width(7)) u_eq_1035 (
        .y(_node_972),
        .a(7'd74),
        .b(_T_1091)
    );
    wire _node_973;
    MUX_UNSIGNED #(.width(1)) u_mux_1036 (
        .y(_node_973),
        .sel(_node_972),
        .a(_T_777_74),
        .b(_node_971)
    );
    wire _node_974;
    EQ_UNSIGNED #(.width(7)) u_eq_1037 (
        .y(_node_974),
        .a(7'd75),
        .b(_T_1091)
    );
    wire _node_975;
    MUX_UNSIGNED #(.width(1)) u_mux_1038 (
        .y(_node_975),
        .sel(_node_974),
        .a(_T_777_75),
        .b(_node_973)
    );
    wire _node_976;
    EQ_UNSIGNED #(.width(7)) u_eq_1039 (
        .y(_node_976),
        .a(7'd76),
        .b(_T_1091)
    );
    wire _node_977;
    MUX_UNSIGNED #(.width(1)) u_mux_1040 (
        .y(_node_977),
        .sel(_node_976),
        .a(_T_777_76),
        .b(_node_975)
    );
    wire _node_978;
    EQ_UNSIGNED #(.width(7)) u_eq_1041 (
        .y(_node_978),
        .a(7'd77),
        .b(_T_1091)
    );
    wire _node_979;
    MUX_UNSIGNED #(.width(1)) u_mux_1042 (
        .y(_node_979),
        .sel(_node_978),
        .a(_T_777_77),
        .b(_node_977)
    );
    wire _node_980;
    EQ_UNSIGNED #(.width(7)) u_eq_1043 (
        .y(_node_980),
        .a(7'd78),
        .b(_T_1091)
    );
    wire _node_981;
    MUX_UNSIGNED #(.width(1)) u_mux_1044 (
        .y(_node_981),
        .sel(_node_980),
        .a(_T_777_78),
        .b(_node_979)
    );
    wire _node_982;
    EQ_UNSIGNED #(.width(7)) u_eq_1045 (
        .y(_node_982),
        .a(7'd79),
        .b(_T_1091)
    );
    wire _node_983;
    MUX_UNSIGNED #(.width(1)) u_mux_1046 (
        .y(_node_983),
        .sel(_node_982),
        .a(_T_777_79),
        .b(_node_981)
    );
    wire _node_984;
    EQ_UNSIGNED #(.width(7)) u_eq_1047 (
        .y(_node_984),
        .a(7'd80),
        .b(_T_1091)
    );
    wire _node_985;
    MUX_UNSIGNED #(.width(1)) u_mux_1048 (
        .y(_node_985),
        .sel(_node_984),
        .a(_T_777_80),
        .b(_node_983)
    );
    wire _node_986;
    EQ_UNSIGNED #(.width(7)) u_eq_1049 (
        .y(_node_986),
        .a(7'd81),
        .b(_T_1091)
    );
    wire _node_987;
    MUX_UNSIGNED #(.width(1)) u_mux_1050 (
        .y(_node_987),
        .sel(_node_986),
        .a(_T_777_81),
        .b(_node_985)
    );
    wire _node_988;
    EQ_UNSIGNED #(.width(7)) u_eq_1051 (
        .y(_node_988),
        .a(7'd82),
        .b(_T_1091)
    );
    wire _node_989;
    MUX_UNSIGNED #(.width(1)) u_mux_1052 (
        .y(_node_989),
        .sel(_node_988),
        .a(_T_777_82),
        .b(_node_987)
    );
    wire _node_990;
    EQ_UNSIGNED #(.width(7)) u_eq_1053 (
        .y(_node_990),
        .a(7'd83),
        .b(_T_1091)
    );
    wire _node_991;
    MUX_UNSIGNED #(.width(1)) u_mux_1054 (
        .y(_node_991),
        .sel(_node_990),
        .a(_T_777_83),
        .b(_node_989)
    );
    wire _node_992;
    EQ_UNSIGNED #(.width(7)) u_eq_1055 (
        .y(_node_992),
        .a(7'd84),
        .b(_T_1091)
    );
    wire _node_993;
    MUX_UNSIGNED #(.width(1)) u_mux_1056 (
        .y(_node_993),
        .sel(_node_992),
        .a(_T_777_84),
        .b(_node_991)
    );
    wire _node_994;
    EQ_UNSIGNED #(.width(7)) u_eq_1057 (
        .y(_node_994),
        .a(7'd85),
        .b(_T_1091)
    );
    wire _node_995;
    MUX_UNSIGNED #(.width(1)) u_mux_1058 (
        .y(_node_995),
        .sel(_node_994),
        .a(_T_777_85),
        .b(_node_993)
    );
    wire _node_996;
    EQ_UNSIGNED #(.width(7)) u_eq_1059 (
        .y(_node_996),
        .a(7'd86),
        .b(_T_1091)
    );
    wire _node_997;
    MUX_UNSIGNED #(.width(1)) u_mux_1060 (
        .y(_node_997),
        .sel(_node_996),
        .a(_T_777_86),
        .b(_node_995)
    );
    wire _node_998;
    EQ_UNSIGNED #(.width(7)) u_eq_1061 (
        .y(_node_998),
        .a(7'd87),
        .b(_T_1091)
    );
    wire _node_999;
    MUX_UNSIGNED #(.width(1)) u_mux_1062 (
        .y(_node_999),
        .sel(_node_998),
        .a(_T_777_87),
        .b(_node_997)
    );
    wire _node_1000;
    EQ_UNSIGNED #(.width(7)) u_eq_1063 (
        .y(_node_1000),
        .a(7'd88),
        .b(_T_1091)
    );
    wire _node_1001;
    MUX_UNSIGNED #(.width(1)) u_mux_1064 (
        .y(_node_1001),
        .sel(_node_1000),
        .a(_T_777_88),
        .b(_node_999)
    );
    wire _node_1002;
    EQ_UNSIGNED #(.width(7)) u_eq_1065 (
        .y(_node_1002),
        .a(7'd89),
        .b(_T_1091)
    );
    wire _node_1003;
    MUX_UNSIGNED #(.width(1)) u_mux_1066 (
        .y(_node_1003),
        .sel(_node_1002),
        .a(_T_777_89),
        .b(_node_1001)
    );
    wire _node_1004;
    EQ_UNSIGNED #(.width(7)) u_eq_1067 (
        .y(_node_1004),
        .a(7'd90),
        .b(_T_1091)
    );
    wire _node_1005;
    MUX_UNSIGNED #(.width(1)) u_mux_1068 (
        .y(_node_1005),
        .sel(_node_1004),
        .a(_T_777_90),
        .b(_node_1003)
    );
    wire _node_1006;
    EQ_UNSIGNED #(.width(7)) u_eq_1069 (
        .y(_node_1006),
        .a(7'd91),
        .b(_T_1091)
    );
    wire _node_1007;
    MUX_UNSIGNED #(.width(1)) u_mux_1070 (
        .y(_node_1007),
        .sel(_node_1006),
        .a(_T_777_91),
        .b(_node_1005)
    );
    wire _node_1008;
    EQ_UNSIGNED #(.width(7)) u_eq_1071 (
        .y(_node_1008),
        .a(7'd92),
        .b(_T_1091)
    );
    wire _node_1009;
    MUX_UNSIGNED #(.width(1)) u_mux_1072 (
        .y(_node_1009),
        .sel(_node_1008),
        .a(_T_777_92),
        .b(_node_1007)
    );
    wire _node_1010;
    EQ_UNSIGNED #(.width(7)) u_eq_1073 (
        .y(_node_1010),
        .a(7'd93),
        .b(_T_1091)
    );
    wire _node_1011;
    MUX_UNSIGNED #(.width(1)) u_mux_1074 (
        .y(_node_1011),
        .sel(_node_1010),
        .a(_T_777_93),
        .b(_node_1009)
    );
    wire _node_1012;
    EQ_UNSIGNED #(.width(7)) u_eq_1075 (
        .y(_node_1012),
        .a(7'd94),
        .b(_T_1091)
    );
    wire _node_1013;
    MUX_UNSIGNED #(.width(1)) u_mux_1076 (
        .y(_node_1013),
        .sel(_node_1012),
        .a(_T_777_94),
        .b(_node_1011)
    );
    wire _node_1014;
    EQ_UNSIGNED #(.width(7)) u_eq_1077 (
        .y(_node_1014),
        .a(7'd95),
        .b(_T_1091)
    );
    wire _node_1015;
    MUX_UNSIGNED #(.width(1)) u_mux_1078 (
        .y(_node_1015),
        .sel(_node_1014),
        .a(_T_777_95),
        .b(_node_1013)
    );
    wire _node_1016;
    EQ_UNSIGNED #(.width(7)) u_eq_1079 (
        .y(_node_1016),
        .a(7'd96),
        .b(_T_1091)
    );
    wire _node_1017;
    MUX_UNSIGNED #(.width(1)) u_mux_1080 (
        .y(_node_1017),
        .sel(_node_1016),
        .a(_T_777_96),
        .b(_node_1015)
    );
    wire _node_1018;
    EQ_UNSIGNED #(.width(7)) u_eq_1081 (
        .y(_node_1018),
        .a(7'd97),
        .b(_T_1091)
    );
    wire _node_1019;
    MUX_UNSIGNED #(.width(1)) u_mux_1082 (
        .y(_node_1019),
        .sel(_node_1018),
        .a(_T_777_97),
        .b(_node_1017)
    );
    wire _node_1020;
    EQ_UNSIGNED #(.width(7)) u_eq_1083 (
        .y(_node_1020),
        .a(7'd98),
        .b(_T_1091)
    );
    wire _node_1021;
    MUX_UNSIGNED #(.width(1)) u_mux_1084 (
        .y(_node_1021),
        .sel(_node_1020),
        .a(_T_777_98),
        .b(_node_1019)
    );
    wire _node_1022;
    EQ_UNSIGNED #(.width(7)) u_eq_1085 (
        .y(_node_1022),
        .a(7'd99),
        .b(_T_1091)
    );
    wire _node_1023;
    MUX_UNSIGNED #(.width(1)) u_mux_1086 (
        .y(_node_1023),
        .sel(_node_1022),
        .a(_T_777_99),
        .b(_node_1021)
    );
    wire _node_1024;
    EQ_UNSIGNED #(.width(7)) u_eq_1087 (
        .y(_node_1024),
        .a(7'd100),
        .b(_T_1091)
    );
    wire _node_1025;
    MUX_UNSIGNED #(.width(1)) u_mux_1088 (
        .y(_node_1025),
        .sel(_node_1024),
        .a(_T_777_100),
        .b(_node_1023)
    );
    wire [8:0] _node_1026;
    MUX_UNSIGNED #(.width(9)) u_mux_1089 (
        .y(_node_1026),
        .sel(_c__io_out_valid),
        .a(_node_821),
        .b(__T_10__q)
    );
    wire _node_1027;
    MUX_UNSIGNED #(.width(1)) u_mux_1090 (
        .y(_node_1027),
        .sel(_c__io_out_valid),
        .a(_node_822),
        .b(__T_13__q)
    );
    wire [6:0] _node_1028;
    MUX_UNSIGNED #(.width(7)) u_mux_1091 (
        .y(_node_1028),
        .sel(_c__io_out_valid),
        .a(_node_823),
        .b(_value_1__q)
    );
    MUX_UNSIGNED #(.width(9)) u_mux_1092 (
        .y(_WTEMP_6),
        .sel(_node_1025),
        .a(_node_1026),
        .b(__T_10__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_1093 (
        .y(_WTEMP_7),
        .sel(_node_1025),
        .a(_node_1027),
        .b(__T_13__q)
    );
    assign _T_135_0 = 1'h1;
    assign _T_135_1 = 1'h1;
    assign _T_135_10 = 1'h1;
    assign _T_135_100 = 1'h0;
    assign _T_135_11 = 1'h1;
    assign _T_135_12 = 1'h1;
    assign _T_135_13 = 1'h1;
    assign _T_135_14 = 1'h1;
    assign _T_135_15 = 1'h1;
    assign _T_135_16 = 1'h1;
    assign _T_135_17 = 1'h1;
    assign _T_135_18 = 1'h1;
    assign _T_135_19 = 1'h1;
    assign _T_135_2 = 1'h1;
    assign _T_135_20 = 1'h1;
    assign _T_135_21 = 1'h1;
    assign _T_135_22 = 1'h1;
    assign _T_135_23 = 1'h1;
    assign _T_135_24 = 1'h1;
    assign _T_135_25 = 1'h1;
    assign _T_135_26 = 1'h1;
    assign _T_135_27 = 1'h1;
    assign _T_135_28 = 1'h1;
    assign _T_135_29 = 1'h1;
    assign _T_135_3 = 1'h1;
    assign _T_135_30 = 1'h1;
    assign _T_135_31 = 1'h1;
    assign _T_135_32 = 1'h1;
    assign _T_135_33 = 1'h1;
    assign _T_135_34 = 1'h1;
    assign _T_135_35 = 1'h1;
    assign _T_135_36 = 1'h1;
    assign _T_135_37 = 1'h1;
    assign _T_135_38 = 1'h1;
    assign _T_135_39 = 1'h1;
    assign _T_135_4 = 1'h1;
    assign _T_135_40 = 1'h1;
    assign _T_135_41 = 1'h1;
    assign _T_135_42 = 1'h1;
    assign _T_135_43 = 1'h1;
    assign _T_135_44 = 1'h1;
    assign _T_135_45 = 1'h1;
    assign _T_135_46 = 1'h1;
    assign _T_135_47 = 1'h1;
    assign _T_135_48 = 1'h1;
    assign _T_135_49 = 1'h1;
    assign _T_135_5 = 1'h1;
    assign _T_135_50 = 1'h1;
    assign _T_135_51 = 1'h1;
    assign _T_135_52 = 1'h1;
    assign _T_135_53 = 1'h1;
    assign _T_135_54 = 1'h1;
    assign _T_135_55 = 1'h1;
    assign _T_135_56 = 1'h1;
    assign _T_135_57 = 1'h1;
    assign _T_135_58 = 1'h1;
    assign _T_135_59 = 1'h1;
    assign _T_135_6 = 1'h1;
    assign _T_135_60 = 1'h1;
    assign _T_135_61 = 1'h1;
    assign _T_135_62 = 1'h1;
    assign _T_135_63 = 1'h1;
    assign _T_135_64 = 1'h1;
    assign _T_135_65 = 1'h1;
    assign _T_135_66 = 1'h1;
    assign _T_135_67 = 1'h1;
    assign _T_135_68 = 1'h1;
    assign _T_135_69 = 1'h1;
    assign _T_135_7 = 1'h1;
    assign _T_135_70 = 1'h1;
    assign _T_135_71 = 1'h1;
    assign _T_135_72 = 1'h1;
    assign _T_135_73 = 1'h1;
    assign _T_135_74 = 1'h1;
    assign _T_135_75 = 1'h1;
    assign _T_135_76 = 1'h1;
    assign _T_135_77 = 1'h1;
    assign _T_135_78 = 1'h1;
    assign _T_135_79 = 1'h1;
    assign _T_135_8 = 1'h1;
    assign _T_135_80 = 1'h1;
    assign _T_135_81 = 1'h1;
    assign _T_135_82 = 1'h1;
    assign _T_135_83 = 1'h1;
    assign _T_135_84 = 1'h1;
    assign _T_135_85 = 1'h1;
    assign _T_135_86 = 1'h1;
    assign _T_135_87 = 1'h1;
    assign _T_135_88 = 1'h1;
    assign _T_135_89 = 1'h1;
    assign _T_135_9 = 1'h1;
    assign _T_135_90 = 1'h1;
    assign _T_135_91 = 1'h1;
    assign _T_135_92 = 1'h1;
    assign _T_135_93 = 1'h1;
    assign _T_135_94 = 1'h1;
    assign _T_135_95 = 1'h1;
    assign _T_135_96 = 1'h1;
    assign _T_135_97 = 1'h1;
    assign _T_135_98 = 1'h1;
    assign _T_135_99 = 1'h1;
    assign _WTEMP_8 = _T_24;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1094 (
        .y(_T_344_0),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1095 (
        .y(_T_344_1),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1096 (
        .y(_T_344_10),
        .in(2'h2)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1097 (
        .y(_T_344_100),
        .in(1'h0)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1098 (
        .y(_T_344_11),
        .in(2'h2)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1099 (
        .y(_T_344_12),
        .in(2'h2)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1100 (
        .y(_T_344_13),
        .in(2'h2)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1101 (
        .y(_T_344_14),
        .in(2'h2)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1102 (
        .y(_T_344_15),
        .in(2'h2)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1103 (
        .y(_T_344_16),
        .in(2'h2)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1104 (
        .y(_T_344_17),
        .in(2'h2)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1105 (
        .y(_T_344_18),
        .in(2'h2)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1106 (
        .y(_T_344_19),
        .in(2'h2)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1107 (
        .y(_T_344_2),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1108 (
        .y(_T_344_20),
        .in(2'h3)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1109 (
        .y(_T_344_21),
        .in(2'h3)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1110 (
        .y(_T_344_22),
        .in(2'h3)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1111 (
        .y(_T_344_23),
        .in(2'h3)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1112 (
        .y(_T_344_24),
        .in(2'h3)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1113 (
        .y(_T_344_25),
        .in(2'h3)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1114 (
        .y(_T_344_26),
        .in(2'h3)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1115 (
        .y(_T_344_27),
        .in(2'h3)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1116 (
        .y(_T_344_28),
        .in(2'h3)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1117 (
        .y(_T_344_29),
        .in(2'h3)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1118 (
        .y(_T_344_3),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1119 (
        .y(_T_344_30),
        .in(3'h4)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1120 (
        .y(_T_344_31),
        .in(3'h4)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1121 (
        .y(_T_344_32),
        .in(3'h4)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1122 (
        .y(_T_344_33),
        .in(3'h4)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1123 (
        .y(_T_344_34),
        .in(3'h4)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1124 (
        .y(_T_344_35),
        .in(3'h4)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1125 (
        .y(_T_344_36),
        .in(3'h4)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1126 (
        .y(_T_344_37),
        .in(3'h4)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1127 (
        .y(_T_344_38),
        .in(3'h4)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1128 (
        .y(_T_344_39),
        .in(3'h4)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1129 (
        .y(_T_344_4),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1130 (
        .y(_T_344_40),
        .in(3'h5)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1131 (
        .y(_T_344_41),
        .in(3'h5)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1132 (
        .y(_T_344_42),
        .in(3'h5)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1133 (
        .y(_T_344_43),
        .in(3'h5)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1134 (
        .y(_T_344_44),
        .in(3'h5)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1135 (
        .y(_T_344_45),
        .in(3'h5)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1136 (
        .y(_T_344_46),
        .in(3'h5)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1137 (
        .y(_T_344_47),
        .in(3'h5)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1138 (
        .y(_T_344_48),
        .in(3'h5)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1139 (
        .y(_T_344_49),
        .in(3'h5)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1140 (
        .y(_T_344_5),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1141 (
        .y(_T_344_50),
        .in(3'h6)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1142 (
        .y(_T_344_51),
        .in(3'h6)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1143 (
        .y(_T_344_52),
        .in(3'h6)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1144 (
        .y(_T_344_53),
        .in(3'h6)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1145 (
        .y(_T_344_54),
        .in(3'h6)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1146 (
        .y(_T_344_55),
        .in(3'h6)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1147 (
        .y(_T_344_56),
        .in(3'h6)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1148 (
        .y(_T_344_57),
        .in(3'h6)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1149 (
        .y(_T_344_58),
        .in(3'h6)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1150 (
        .y(_T_344_59),
        .in(3'h6)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1151 (
        .y(_T_344_6),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1152 (
        .y(_T_344_60),
        .in(3'h7)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1153 (
        .y(_T_344_61),
        .in(3'h7)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1154 (
        .y(_T_344_62),
        .in(3'h7)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1155 (
        .y(_T_344_63),
        .in(3'h7)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1156 (
        .y(_T_344_64),
        .in(3'h7)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1157 (
        .y(_T_344_65),
        .in(3'h7)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1158 (
        .y(_T_344_66),
        .in(3'h7)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1159 (
        .y(_T_344_67),
        .in(3'h7)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1160 (
        .y(_T_344_68),
        .in(3'h7)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1161 (
        .y(_T_344_69),
        .in(3'h7)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1162 (
        .y(_T_344_7),
        .in(1'h1)
    );
    assign _T_344_70 = 4'h8;
    assign _T_344_71 = 4'h8;
    assign _T_344_72 = 4'h8;
    assign _T_344_73 = 4'h8;
    assign _T_344_74 = 4'h8;
    assign _T_344_75 = 4'h8;
    assign _T_344_76 = 4'h8;
    assign _T_344_77 = 4'h8;
    assign _T_344_78 = 4'h8;
    assign _T_344_79 = 4'h8;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1163 (
        .y(_T_344_8),
        .in(1'h1)
    );
    assign _T_344_80 = 4'h9;
    assign _T_344_81 = 4'h9;
    assign _T_344_82 = 4'h9;
    assign _T_344_83 = 4'h9;
    assign _T_344_84 = 4'h9;
    assign _T_344_85 = 4'h9;
    assign _T_344_86 = 4'h9;
    assign _T_344_87 = 4'h9;
    assign _T_344_88 = 4'h9;
    assign _T_344_89 = 4'h9;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1164 (
        .y(_T_344_9),
        .in(1'h1)
    );
    assign _T_344_90 = 4'hA;
    assign _T_344_91 = 4'hA;
    assign _T_344_92 = 4'hA;
    assign _T_344_93 = 4'hA;
    assign _T_344_94 = 4'hA;
    assign _T_344_95 = 4'hA;
    assign _T_344_96 = 4'hA;
    assign _T_344_97 = 4'hA;
    assign _T_344_98 = 4'hA;
    assign _T_344_99 = 4'hA;
    MUX_UNSIGNED #(.width(9)) u_mux_1165 (
        .y(_WTEMP_4),
        .sel(_T_659),
        .a(_node_615),
        .b(__T_4__q)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1166 (
        .y(_T_551_0),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1167 (
        .y(_T_551_1),
        .in(2'h2)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1168 (
        .y(_T_551_10),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1169 (
        .y(_T_551_100),
        .in(1'h0)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1170 (
        .y(_T_551_11),
        .in(2'h2)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1171 (
        .y(_T_551_12),
        .in(2'h3)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1172 (
        .y(_T_551_13),
        .in(3'h4)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1173 (
        .y(_T_551_14),
        .in(3'h5)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1174 (
        .y(_T_551_15),
        .in(3'h6)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1175 (
        .y(_T_551_16),
        .in(3'h7)
    );
    assign _T_551_17 = 4'h8;
    assign _T_551_18 = 4'h9;
    assign _T_551_19 = 4'hA;
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1176 (
        .y(_T_551_2),
        .in(2'h3)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1177 (
        .y(_T_551_20),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1178 (
        .y(_T_551_21),
        .in(2'h2)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1179 (
        .y(_T_551_22),
        .in(2'h3)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1180 (
        .y(_T_551_23),
        .in(3'h4)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1181 (
        .y(_T_551_24),
        .in(3'h5)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1182 (
        .y(_T_551_25),
        .in(3'h6)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1183 (
        .y(_T_551_26),
        .in(3'h7)
    );
    assign _T_551_27 = 4'h8;
    assign _T_551_28 = 4'h9;
    assign _T_551_29 = 4'hA;
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1184 (
        .y(_T_551_3),
        .in(3'h4)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1185 (
        .y(_T_551_30),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1186 (
        .y(_T_551_31),
        .in(2'h2)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1187 (
        .y(_T_551_32),
        .in(2'h3)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1188 (
        .y(_T_551_33),
        .in(3'h4)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1189 (
        .y(_T_551_34),
        .in(3'h5)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1190 (
        .y(_T_551_35),
        .in(3'h6)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1191 (
        .y(_T_551_36),
        .in(3'h7)
    );
    assign _T_551_37 = 4'h8;
    assign _T_551_38 = 4'h9;
    assign _T_551_39 = 4'hA;
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1192 (
        .y(_T_551_4),
        .in(3'h5)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1193 (
        .y(_T_551_40),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1194 (
        .y(_T_551_41),
        .in(2'h2)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1195 (
        .y(_T_551_42),
        .in(2'h3)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1196 (
        .y(_T_551_43),
        .in(3'h4)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1197 (
        .y(_T_551_44),
        .in(3'h5)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1198 (
        .y(_T_551_45),
        .in(3'h6)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1199 (
        .y(_T_551_46),
        .in(3'h7)
    );
    assign _T_551_47 = 4'h8;
    assign _T_551_48 = 4'h9;
    assign _T_551_49 = 4'hA;
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1200 (
        .y(_T_551_5),
        .in(3'h6)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1201 (
        .y(_T_551_50),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1202 (
        .y(_T_551_51),
        .in(2'h2)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1203 (
        .y(_T_551_52),
        .in(2'h3)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1204 (
        .y(_T_551_53),
        .in(3'h4)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1205 (
        .y(_T_551_54),
        .in(3'h5)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1206 (
        .y(_T_551_55),
        .in(3'h6)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1207 (
        .y(_T_551_56),
        .in(3'h7)
    );
    assign _T_551_57 = 4'h8;
    assign _T_551_58 = 4'h9;
    assign _T_551_59 = 4'hA;
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1208 (
        .y(_T_551_6),
        .in(3'h7)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1209 (
        .y(_T_551_60),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1210 (
        .y(_T_551_61),
        .in(2'h2)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1211 (
        .y(_T_551_62),
        .in(2'h3)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1212 (
        .y(_T_551_63),
        .in(3'h4)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1213 (
        .y(_T_551_64),
        .in(3'h5)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1214 (
        .y(_T_551_65),
        .in(3'h6)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1215 (
        .y(_T_551_66),
        .in(3'h7)
    );
    assign _T_551_67 = 4'h8;
    assign _T_551_68 = 4'h9;
    assign _T_551_69 = 4'hA;
    assign _T_551_7 = 4'h8;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1216 (
        .y(_T_551_70),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1217 (
        .y(_T_551_71),
        .in(2'h2)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1218 (
        .y(_T_551_72),
        .in(2'h3)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1219 (
        .y(_T_551_73),
        .in(3'h4)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1220 (
        .y(_T_551_74),
        .in(3'h5)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1221 (
        .y(_T_551_75),
        .in(3'h6)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1222 (
        .y(_T_551_76),
        .in(3'h7)
    );
    assign _T_551_77 = 4'h8;
    assign _T_551_78 = 4'h9;
    assign _T_551_79 = 4'hA;
    assign _T_551_8 = 4'h9;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1223 (
        .y(_T_551_80),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1224 (
        .y(_T_551_81),
        .in(2'h2)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1225 (
        .y(_T_551_82),
        .in(2'h3)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1226 (
        .y(_T_551_83),
        .in(3'h4)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1227 (
        .y(_T_551_84),
        .in(3'h5)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1228 (
        .y(_T_551_85),
        .in(3'h6)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1229 (
        .y(_T_551_86),
        .in(3'h7)
    );
    assign _T_551_87 = 4'h8;
    assign _T_551_88 = 4'h9;
    assign _T_551_89 = 4'hA;
    assign _T_551_9 = 4'hA;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1230 (
        .y(_T_551_90),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1231 (
        .y(_T_551_91),
        .in(2'h2)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1232 (
        .y(_T_551_92),
        .in(2'h3)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1233 (
        .y(_T_551_93),
        .in(3'h4)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1234 (
        .y(_T_551_94),
        .in(3'h5)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1235 (
        .y(_T_551_95),
        .in(3'h6)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1236 (
        .y(_T_551_96),
        .in(3'h7)
    );
    assign _T_551_97 = 4'h8;
    assign _T_551_98 = 4'h9;
    assign _T_551_99 = 4'hA;
    MUX_UNSIGNED #(.width(1)) u_mux_1237 (
        .y(_WTEMP_5),
        .sel(_T_659),
        .a(_node_616),
        .b(__T_7__q)
    );
    assign _T_777_0 = 1'h1;
    assign _T_777_1 = 1'h1;
    assign _T_777_10 = 1'h1;
    assign _T_777_100 = 1'h0;
    assign _T_777_11 = 1'h1;
    assign _T_777_12 = 1'h1;
    assign _T_777_13 = 1'h1;
    assign _T_777_14 = 1'h1;
    assign _T_777_15 = 1'h1;
    assign _T_777_16 = 1'h1;
    assign _T_777_17 = 1'h1;
    assign _T_777_18 = 1'h1;
    assign _T_777_19 = 1'h1;
    assign _T_777_2 = 1'h1;
    assign _T_777_20 = 1'h1;
    assign _T_777_21 = 1'h1;
    assign _T_777_22 = 1'h1;
    assign _T_777_23 = 1'h1;
    assign _T_777_24 = 1'h1;
    assign _T_777_25 = 1'h1;
    assign _T_777_26 = 1'h1;
    assign _T_777_27 = 1'h1;
    assign _T_777_28 = 1'h1;
    assign _T_777_29 = 1'h1;
    assign _T_777_3 = 1'h1;
    assign _T_777_30 = 1'h1;
    assign _T_777_31 = 1'h1;
    assign _T_777_32 = 1'h1;
    assign _T_777_33 = 1'h1;
    assign _T_777_34 = 1'h1;
    assign _T_777_35 = 1'h1;
    assign _T_777_36 = 1'h1;
    assign _T_777_37 = 1'h1;
    assign _T_777_38 = 1'h1;
    assign _T_777_39 = 1'h1;
    assign _T_777_4 = 1'h1;
    assign _T_777_40 = 1'h1;
    assign _T_777_41 = 1'h1;
    assign _T_777_42 = 1'h1;
    assign _T_777_43 = 1'h1;
    assign _T_777_44 = 1'h1;
    assign _T_777_45 = 1'h1;
    assign _T_777_46 = 1'h1;
    assign _T_777_47 = 1'h1;
    assign _T_777_48 = 1'h1;
    assign _T_777_49 = 1'h1;
    assign _T_777_5 = 1'h1;
    assign _T_777_50 = 1'h1;
    assign _T_777_51 = 1'h1;
    assign _T_777_52 = 1'h1;
    assign _T_777_53 = 1'h1;
    assign _T_777_54 = 1'h1;
    assign _T_777_55 = 1'h1;
    assign _T_777_56 = 1'h1;
    assign _T_777_57 = 1'h1;
    assign _T_777_58 = 1'h1;
    assign _T_777_59 = 1'h1;
    assign _T_777_6 = 1'h1;
    assign _T_777_60 = 1'h1;
    assign _T_777_61 = 1'h1;
    assign _T_777_62 = 1'h1;
    assign _T_777_63 = 1'h1;
    assign _T_777_64 = 1'h1;
    assign _T_777_65 = 1'h1;
    assign _T_777_66 = 1'h1;
    assign _T_777_67 = 1'h1;
    assign _T_777_68 = 1'h1;
    assign _T_777_69 = 1'h1;
    assign _T_777_7 = 1'h1;
    assign _T_777_70 = 1'h1;
    assign _T_777_71 = 1'h1;
    assign _T_777_72 = 1'h1;
    assign _T_777_73 = 1'h1;
    assign _T_777_74 = 1'h1;
    assign _T_777_75 = 1'h1;
    assign _T_777_76 = 1'h1;
    assign _T_777_77 = 1'h1;
    assign _T_777_78 = 1'h1;
    assign _T_777_79 = 1'h1;
    assign _T_777_8 = 1'h1;
    assign _T_777_80 = 1'h1;
    assign _T_777_81 = 1'h1;
    assign _T_777_82 = 1'h1;
    assign _T_777_83 = 1'h1;
    assign _T_777_84 = 1'h1;
    assign _T_777_85 = 1'h1;
    assign _T_777_86 = 1'h1;
    assign _T_777_87 = 1'h1;
    assign _T_777_88 = 1'h1;
    assign _T_777_89 = 1'h1;
    assign _T_777_9 = 1'h1;
    assign _T_777_90 = 1'h1;
    assign _T_777_91 = 1'h1;
    assign _T_777_92 = 1'h1;
    assign _T_777_93 = 1'h1;
    assign _T_777_94 = 1'h1;
    assign _T_777_95 = 1'h1;
    assign _T_777_96 = 1'h1;
    assign _T_777_97 = 1'h1;
    assign _T_777_98 = 1'h1;
    assign _T_777_99 = 1'h1;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1238 (
        .y(_T_986_0),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1239 (
        .y(_T_986_1),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1240 (
        .y(_T_986_10),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1241 (
        .y(_T_986_100),
        .in(1'h0)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1242 (
        .y(_T_986_11),
        .in(2'h2)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1243 (
        .y(_T_986_12),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1244 (
        .y(_T_986_13),
        .in(2'h2)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1245 (
        .y(_T_986_14),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1246 (
        .y(_T_986_15),
        .in(2'h2)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1247 (
        .y(_T_986_16),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1248 (
        .y(_T_986_17),
        .in(2'h2)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1249 (
        .y(_T_986_18),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1250 (
        .y(_T_986_19),
        .in(2'h2)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1251 (
        .y(_T_986_2),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1252 (
        .y(_T_986_20),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1253 (
        .y(_T_986_21),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1254 (
        .y(_T_986_22),
        .in(2'h3)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1255 (
        .y(_T_986_23),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1256 (
        .y(_T_986_24),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1257 (
        .y(_T_986_25),
        .in(2'h3)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1258 (
        .y(_T_986_26),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1259 (
        .y(_T_986_27),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1260 (
        .y(_T_986_28),
        .in(2'h3)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1261 (
        .y(_T_986_29),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1262 (
        .y(_T_986_3),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1263 (
        .y(_T_986_30),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1264 (
        .y(_T_986_31),
        .in(2'h2)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1265 (
        .y(_T_986_32),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1266 (
        .y(_T_986_33),
        .in(3'h4)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1267 (
        .y(_T_986_34),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1268 (
        .y(_T_986_35),
        .in(2'h2)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1269 (
        .y(_T_986_36),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1270 (
        .y(_T_986_37),
        .in(3'h4)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1271 (
        .y(_T_986_38),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1272 (
        .y(_T_986_39),
        .in(2'h2)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1273 (
        .y(_T_986_4),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1274 (
        .y(_T_986_40),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1275 (
        .y(_T_986_41),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1276 (
        .y(_T_986_42),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1277 (
        .y(_T_986_43),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1278 (
        .y(_T_986_44),
        .in(3'h5)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1279 (
        .y(_T_986_45),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1280 (
        .y(_T_986_46),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1281 (
        .y(_T_986_47),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1282 (
        .y(_T_986_48),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1283 (
        .y(_T_986_49),
        .in(3'h5)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1284 (
        .y(_T_986_5),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1285 (
        .y(_T_986_50),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1286 (
        .y(_T_986_51),
        .in(2'h2)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1287 (
        .y(_T_986_52),
        .in(2'h3)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1288 (
        .y(_T_986_53),
        .in(2'h2)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1289 (
        .y(_T_986_54),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1290 (
        .y(_T_986_55),
        .in(3'h6)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1291 (
        .y(_T_986_56),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1292 (
        .y(_T_986_57),
        .in(2'h2)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1293 (
        .y(_T_986_58),
        .in(2'h3)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1294 (
        .y(_T_986_59),
        .in(2'h2)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1295 (
        .y(_T_986_6),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1296 (
        .y(_T_986_60),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1297 (
        .y(_T_986_61),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1298 (
        .y(_T_986_62),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1299 (
        .y(_T_986_63),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1300 (
        .y(_T_986_64),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1301 (
        .y(_T_986_65),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1302 (
        .y(_T_986_66),
        .in(3'h7)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1303 (
        .y(_T_986_67),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1304 (
        .y(_T_986_68),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1305 (
        .y(_T_986_69),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1306 (
        .y(_T_986_7),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1307 (
        .y(_T_986_70),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1308 (
        .y(_T_986_71),
        .in(2'h2)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1309 (
        .y(_T_986_72),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1310 (
        .y(_T_986_73),
        .in(3'h4)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1311 (
        .y(_T_986_74),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1312 (
        .y(_T_986_75),
        .in(2'h2)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1313 (
        .y(_T_986_76),
        .in(1'h1)
    );
    assign _T_986_77 = 4'h8;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1314 (
        .y(_T_986_78),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1315 (
        .y(_T_986_79),
        .in(2'h2)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1316 (
        .y(_T_986_8),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1317 (
        .y(_T_986_80),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1318 (
        .y(_T_986_81),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1319 (
        .y(_T_986_82),
        .in(2'h3)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1320 (
        .y(_T_986_83),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1321 (
        .y(_T_986_84),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1322 (
        .y(_T_986_85),
        .in(2'h3)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1323 (
        .y(_T_986_86),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1324 (
        .y(_T_986_87),
        .in(1'h1)
    );
    assign _T_986_88 = 4'h9;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1325 (
        .y(_T_986_89),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1326 (
        .y(_T_986_9),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1327 (
        .y(_T_986_90),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1328 (
        .y(_T_986_91),
        .in(2'h2)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1329 (
        .y(_T_986_92),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1330 (
        .y(_T_986_93),
        .in(2'h2)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1331 (
        .y(_T_986_94),
        .in(3'h5)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1332 (
        .y(_T_986_95),
        .in(2'h2)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1333 (
        .y(_T_986_96),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1334 (
        .y(_T_986_97),
        .in(2'h2)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1335 (
        .y(_T_986_98),
        .in(1'h1)
    );
    assign _T_986_99 = 4'hA;
    assign _c__clock = clock;
    PAD_UNSIGNED #(.width(4), .n(16)) u_pad_1336 (
        .y(_c__io_in_bits_a),
        .in(_node_209)
    );
    PAD_UNSIGNED #(.width(4), .n(16)) u_pad_1337 (
        .y(_c__io_in_bits_b),
        .in(_node_411)
    );
    assign _c__io_in_valid = _node_613;
    assign _c__reset = reset;
    MUX_UNSIGNED #(.width(7)) u_mux_1338 (
        .y(_WTEMP_10),
        .sel(_T_659),
        .a(_node_617),
        .b(_value__q)
    );
    MUX_UNSIGNED #(.width(7)) u_mux_1339 (
        .y(_WTEMP_15),
        .sel(_node_1025),
        .a(_node_1028),
        .b(_value_1__q)
    );
endmodule //DecoupledRealGCDTests4
module RealGCD(
    input clock,
    input reset,
    output io_in_ready,
    input io_in_valid,
    input [15:0] io_in_bits_a,
    input [15:0] io_in_bits_b,
    output io_out_valid,
    output [15:0] io_out_bits
);
    wire [15:0] _x__q;
    wire [15:0] _x__d;
    DFF_POSCLK #(.width(16)) x (
        .q(_x__q),
        .d(_x__d),
        .clk(clock)
    );
    wire [15:0] _y__q;
    wire [15:0] _y__d;
    DFF_POSCLK #(.width(16)) y (
        .q(_y__q),
        .d(_y__d),
        .clk(clock)
    );
    wire _p__q;
    wire _p__d;
    DFF_POSCLK #(.width(1)) p (
        .q(_p__q),
        .d(_p__d),
        .clk(clock)
    );
    wire _WTEMP_0;
    MUX_UNSIGNED #(.width(1)) u_mux_1 (
        .y(_p__d),
        .sel(reset),
        .a(1'h0),
        .b(_WTEMP_0)
    );
    wire [15:0] _ti__q;
    wire [15:0] _ti__d;
    DFF_POSCLK #(.width(16)) ti (
        .q(_ti__q),
        .d(_ti__d),
        .clk(clock)
    );
    wire [15:0] _WTEMP_1;
    MUX_UNSIGNED #(.width(16)) u_mux_2 (
        .y(_ti__d),
        .sel(reset),
        .a(16'h0),
        .b(_WTEMP_1)
    );
    wire [16:0] _T_20;
    wire [15:0] _WTEMP_2;
    PAD_UNSIGNED #(.width(1), .n(16)) u_pad_3 (
        .y(_WTEMP_2),
        .in(1'h1)
    );
    ADD_UNSIGNED #(.width(16)) u_add_4 (
        .y(_T_20),
        .a(_ti__q),
        .b(_WTEMP_2)
    );
    wire [15:0] _T_21;
    TAIL #(.width(17), .n(1)) tail_5 (
        .y(_T_21),
        .in(_T_20)
    );
    wire _T_23;
    EQ_UNSIGNED #(.width(1)) u_eq_6 (
        .y(_T_23),
        .a(_p__q),
        .b(1'h0)
    );
    wire _T_25;
    EQ_UNSIGNED #(.width(1)) u_eq_7 (
        .y(_T_25),
        .a(_p__q),
        .b(1'h0)
    );
    wire _T_26;
    BITWISEAND #(.width(1)) bitwiseand_8 (
        .y(_T_26),
        .a(io_in_valid),
        .b(_T_25)
    );
    wire _T_28;
    GT_UNSIGNED #(.width(16)) u_gt_9 (
        .y(_T_28),
        .a(_x__q),
        .b(_y__q)
    );
    wire [15:0] _node_0;
    MUX_UNSIGNED #(.width(16)) u_mux_10 (
        .y(_node_0),
        .sel(_T_26),
        .a(io_in_bits_a),
        .b(_x__q)
    );
    wire [15:0] _node_1;
    MUX_UNSIGNED #(.width(16)) u_mux_11 (
        .y(_node_1),
        .sel(_T_26),
        .a(io_in_bits_b),
        .b(_y__q)
    );
    wire _T_30;
    EQ_UNSIGNED #(.width(1)) u_eq_12 (
        .y(_T_30),
        .a(_T_28),
        .b(1'h0)
    );
    wire [16:0] _T_31;
    SUB_UNSIGNED #(.width(16)) u_sub_13 (
        .y(_T_31),
        .a(_y__q),
        .b(_x__q)
    );
    wire [16:0] _T_32;
    ASUINT #(.width(17)) asuint_14 (
        .y(_T_32),
        .in(_T_31)
    );
    wire [15:0] _T_33;
    TAIL #(.width(17), .n(1)) tail_15 (
        .y(_T_33),
        .in(_T_32)
    );
    wire [15:0] _node_2;
    MUX_UNSIGNED #(.width(16)) u_mux_16 (
        .y(_node_2),
        .sel(_T_28),
        .a(_x__q),
        .b(_node_1)
    );
    wire [15:0] _node_3;
    MUX_UNSIGNED #(.width(16)) u_mux_17 (
        .y(_node_3),
        .sel(_T_28),
        .a(_y__q),
        .b(_node_0)
    );
    wire [15:0] _node_4;
    MUX_UNSIGNED #(.width(16)) u_mux_18 (
        .y(_node_4),
        .sel(_T_26),
        .a(io_in_bits_a),
        .b(_x__q)
    );
    wire [15:0] _node_5;
    MUX_UNSIGNED #(.width(16)) u_mux_19 (
        .y(_node_5),
        .sel(_T_30),
        .a(_T_33),
        .b(_node_2)
    );
    wire [15:0] _node_6;
    MUX_UNSIGNED #(.width(16)) u_mux_20 (
        .y(_node_6),
        .sel(_T_26),
        .a(io_in_bits_b),
        .b(_y__q)
    );
    wire _T_36;
    EQ_UNSIGNED #(.width(1)) u_eq_21 (
        .y(_T_36),
        .a(reset),
        .b(1'h0)
    );
    wire _T_38;
    wire [15:0] _WTEMP_3;
    PAD_UNSIGNED #(.width(1), .n(16)) u_pad_22 (
        .y(_WTEMP_3),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(16)) u_eq_23 (
        .y(_T_38),
        .a(_y__q),
        .b(_WTEMP_3)
    );
    wire _T_39;
    BITWISEAND #(.width(1)) bitwiseand_24 (
        .y(_T_39),
        .a(_T_38),
        .b(_p__q)
    );
    wire _node_7;
    MUX_UNSIGNED #(.width(1)) u_mux_25 (
        .y(_node_7),
        .sel(_T_26),
        .a(1'h1),
        .b(_p__q)
    );
    assign io_in_ready = _T_23;
    assign io_out_bits = _x__q;
    assign io_out_valid = _T_39;
    MUX_UNSIGNED #(.width(1)) u_mux_26 (
        .y(_WTEMP_0),
        .sel(io_out_valid),
        .a(1'h0),
        .b(_node_7)
    );
    assign _WTEMP_1 = _T_21;
    MUX_UNSIGNED #(.width(16)) u_mux_27 (
        .y(_x__d),
        .sel(_p__q),
        .a(_node_3),
        .b(_node_4)
    );
    MUX_UNSIGNED #(.width(16)) u_mux_28 (
        .y(_y__d),
        .sel(_p__q),
        .a(_node_5),
        .b(_node_6)
    );
endmodule //RealGCD
module DFF_POSCLK(q, d, clk);
    parameter width = 4;
    output reg [width-1:0] q;
    input [width-1:0] d;
    input clk;
    always @(posedge clk) begin
        q <= d;
    end
endmodule // DFF_POSCLK
module MUX_UNSIGNED(y, sel, a, b);
    parameter width = 4;
    output [width-1:0] y;
    input sel;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = sel ? a : b;
endmodule // MUX_UNSIGNED
module PAD_UNSIGNED(y, in);
    parameter width = 4;
    parameter n = 4;
    output [(n > width ? n : width)-1:0] y;
    input [width-1:0] in;
    assign y = (n > width) ? {{(n - width){1'b0}}, in} : in;
endmodule // PAD_UNSIGNED
module ADD_UNSIGNED(y, a, b);
    parameter width = 4;
    output [width:0] y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a + b;
endmodule // ADD_UNSIGNED
module TAIL(y, in);
    parameter width = 4;
    parameter n = 2;
    output [width-n-1:0] y;
    input [width-1:0] in;
    assign y = in[width-n-1:0];
endmodule // TAIL
module EQ_UNSIGNED(y, a, b);
    parameter width = 4;
    output y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a == b;
endmodule // EQ_UNSIGNED
module BITWISEAND(y, a, b);
    parameter width = 4;
    output [width-1:0] y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a & b;
endmodule // BITWISEAND
module GT_UNSIGNED(y, a, b);
    parameter width = 4;
    output y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a > b;
endmodule // GT_UNSIGNED
module SUB_UNSIGNED(y, a, b);
    parameter width = 4;
    output [width:0] y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a - b;
endmodule // SUB_UNSIGNED
module ASUINT(y, in);
    parameter width = 4;
    output [width-1:0] y;
    input [width-1:0] in;
    assign y = $unsigned(in);
endmodule // ASUINT
module BITS(y, in);
    parameter width = 4;
    parameter high = 2;
    parameter low = 0;
    output [high-low:0] y;
    input [width-1:0] in;
    assign y = in[high:low];
endmodule // BITS
module NEQ_UNSIGNED(y, a, b);
    parameter width = 4;
    output y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a != b;
endmodule // NEQ_UNSIGNED
module BITWISEOR(y, a, b);
    parameter width = 4;
    output [width-1:0] y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a | b;
endmodule // BITWISEOR
