module DynamicMemorySearch(
  input        clock,
  input        reset,
  input        io_isWr,
  input  [2:0] io_wrAddr,
  input  [3:0] io_data,
  input        io_en,
  output [2:0] io_target,
  output       io_done
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] list [0:7]; // @[DynamicMemorySearch.scala 19:19]
  wire  list_memVal_en; // @[DynamicMemorySearch.scala 19:19]
  wire [2:0] list_memVal_addr; // @[DynamicMemorySearch.scala 19:19]
  wire [3:0] list_memVal_data; // @[DynamicMemorySearch.scala 19:19]
  wire [3:0] list__T_19_data; // @[DynamicMemorySearch.scala 19:19]
  wire [2:0] list__T_19_addr; // @[DynamicMemorySearch.scala 19:19]
  wire  list__T_19_mask; // @[DynamicMemorySearch.scala 19:19]
  wire  list__T_19_en; // @[DynamicMemorySearch.scala 19:19]
  wire [3:0] list__T_22_data; // @[DynamicMemorySearch.scala 19:19]
  wire [2:0] list__T_22_addr; // @[DynamicMemorySearch.scala 19:19]
  wire  list__T_22_mask; // @[DynamicMemorySearch.scala 19:19]
  wire  list__T_22_en; // @[DynamicMemorySearch.scala 19:19]
  wire [3:0] list__T_25_data; // @[DynamicMemorySearch.scala 19:19]
  wire [2:0] list__T_25_addr; // @[DynamicMemorySearch.scala 19:19]
  wire  list__T_25_mask; // @[DynamicMemorySearch.scala 19:19]
  wire  list__T_25_en; // @[DynamicMemorySearch.scala 19:19]
  wire [3:0] list__T_28_data; // @[DynamicMemorySearch.scala 19:19]
  wire [2:0] list__T_28_addr; // @[DynamicMemorySearch.scala 19:19]
  wire  list__T_28_mask; // @[DynamicMemorySearch.scala 19:19]
  wire  list__T_28_en; // @[DynamicMemorySearch.scala 19:19]
  wire [3:0] list__T_31_data; // @[DynamicMemorySearch.scala 19:19]
  wire [2:0] list__T_31_addr; // @[DynamicMemorySearch.scala 19:19]
  wire  list__T_31_mask; // @[DynamicMemorySearch.scala 19:19]
  wire  list__T_31_en; // @[DynamicMemorySearch.scala 19:19]
  wire [3:0] list__T_34_data; // @[DynamicMemorySearch.scala 19:19]
  wire [2:0] list__T_34_addr; // @[DynamicMemorySearch.scala 19:19]
  wire  list__T_34_mask; // @[DynamicMemorySearch.scala 19:19]
  wire  list__T_34_en; // @[DynamicMemorySearch.scala 19:19]
  wire [3:0] list__T_37_data; // @[DynamicMemorySearch.scala 19:19]
  wire [2:0] list__T_37_addr; // @[DynamicMemorySearch.scala 19:19]
  wire  list__T_37_mask; // @[DynamicMemorySearch.scala 19:19]
  wire  list__T_37_en; // @[DynamicMemorySearch.scala 19:19]
  wire [3:0] list__T_40_data; // @[DynamicMemorySearch.scala 19:19]
  wire [2:0] list__T_40_addr; // @[DynamicMemorySearch.scala 19:19]
  wire  list__T_40_mask; // @[DynamicMemorySearch.scala 19:19]
  wire  list__T_40_en; // @[DynamicMemorySearch.scala 19:19]
  wire [3:0] list__T_42_data; // @[DynamicMemorySearch.scala 19:19]
  wire [2:0] list__T_42_addr; // @[DynamicMemorySearch.scala 19:19]
  wire  list__T_42_mask; // @[DynamicMemorySearch.scala 19:19]
  wire  list__T_42_en; // @[DynamicMemorySearch.scala 19:19]
  reg [2:0] index; // @[DynamicMemorySearch.scala 18:23]
  wire  _T_13 = ~io_en; // @[DynamicMemorySearch.scala 21:16]
  wire  over = ~io_en & (list_memVal_data == io_data | index == 3'h7); // @[DynamicMemorySearch.scala 21:23]
  wire  _T_44 = ~io_isWr; // @[DynamicMemorySearch.scala 28:18]
  wire  _T_53 = _T_44 & _T_13; // @[DynamicMemorySearch.scala 30:23]
  wire [2:0] _T_57 = index + 3'h1; // @[DynamicMemorySearch.scala 33:20]
  assign list_memVal_en = 1'h1;
  assign list_memVal_addr = index;
  assign list_memVal_data = list[list_memVal_addr]; // @[DynamicMemorySearch.scala 19:19]
  assign list__T_19_data = 4'h0;
  assign list__T_19_addr = 3'h0;
  assign list__T_19_mask = 1'h1;
  assign list__T_19_en = reset;
  assign list__T_22_data = 4'h0;
  assign list__T_22_addr = 3'h1;
  assign list__T_22_mask = 1'h1;
  assign list__T_22_en = reset;
  assign list__T_25_data = 4'h0;
  assign list__T_25_addr = 3'h2;
  assign list__T_25_mask = 1'h1;
  assign list__T_25_en = reset;
  assign list__T_28_data = 4'h0;
  assign list__T_28_addr = 3'h3;
  assign list__T_28_mask = 1'h1;
  assign list__T_28_en = reset;
  assign list__T_31_data = 4'h0;
  assign list__T_31_addr = 3'h4;
  assign list__T_31_mask = 1'h1;
  assign list__T_31_en = reset;
  assign list__T_34_data = 4'h0;
  assign list__T_34_addr = 3'h5;
  assign list__T_34_mask = 1'h1;
  assign list__T_34_en = reset;
  assign list__T_37_data = 4'h0;
  assign list__T_37_addr = 3'h6;
  assign list__T_37_mask = 1'h1;
  assign list__T_37_en = reset;
  assign list__T_40_data = 4'h0;
  assign list__T_40_addr = 3'h7;
  assign list__T_40_mask = 1'h1;
  assign list__T_40_en = reset;
  assign list__T_42_data = io_data;
  assign list__T_42_addr = io_wrAddr;
  assign list__T_42_mask = 1'h1;
  assign list__T_42_en = io_isWr;
  assign io_target = index; // @[DynamicMemorySearch.scala 36:13]
  assign io_done = ~io_en & (list_memVal_data == io_data | index == 3'h7); // @[DynamicMemorySearch.scala 21:23]
  always @(posedge clock) begin
    if (list__T_19_en & list__T_19_mask) begin
      list[list__T_19_addr] <= list__T_19_data; // @[DynamicMemorySearch.scala 19:19]
    end
    if (list__T_22_en & list__T_22_mask) begin
      list[list__T_22_addr] <= list__T_22_data; // @[DynamicMemorySearch.scala 19:19]
    end
    if (list__T_25_en & list__T_25_mask) begin
      list[list__T_25_addr] <= list__T_25_data; // @[DynamicMemorySearch.scala 19:19]
    end
    if (list__T_28_en & list__T_28_mask) begin
      list[list__T_28_addr] <= list__T_28_data; // @[DynamicMemorySearch.scala 19:19]
    end
    if (list__T_31_en & list__T_31_mask) begin
      list[list__T_31_addr] <= list__T_31_data; // @[DynamicMemorySearch.scala 19:19]
    end
    if (list__T_34_en & list__T_34_mask) begin
      list[list__T_34_addr] <= list__T_34_data; // @[DynamicMemorySearch.scala 19:19]
    end
    if (list__T_37_en & list__T_37_mask) begin
      list[list__T_37_addr] <= list__T_37_data; // @[DynamicMemorySearch.scala 19:19]
    end
    if (list__T_40_en & list__T_40_mask) begin
      list[list__T_40_addr] <= list__T_40_data; // @[DynamicMemorySearch.scala 19:19]
    end
    if (list__T_42_en & list__T_42_mask) begin
      list[list__T_42_addr] <= list__T_42_data; // @[DynamicMemorySearch.scala 19:19]
    end
    if (reset) begin // @[DynamicMemorySearch.scala 18:23]
      index <= 3'h0; // @[DynamicMemorySearch.scala 18:23]
    end else if (_T_53 & ~over) begin // @[DynamicMemorySearch.scala 32:34]
      index <= _T_57; // @[DynamicMemorySearch.scala 33:11]
    end else if (_T_44 & io_en) begin // @[DynamicMemorySearch.scala 30:23]
      index <= 3'h0; // @[DynamicMemorySearch.scala 31:11]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    list[initvar] = _RAND_0[3:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  index = _RAND_1[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DynamicMemorySearchTests(
  input   clock,
  input   reset
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  c_clock; // @[DynamicMemorySearch.scala 40:33]
  wire  c_reset; // @[DynamicMemorySearch.scala 40:33]
  wire  c_io_isWr; // @[DynamicMemorySearch.scala 40:33]
  wire [2:0] c_io_wrAddr; // @[DynamicMemorySearch.scala 40:33]
  wire [3:0] c_io_data; // @[DynamicMemorySearch.scala 40:33]
  wire  c_io_en; // @[DynamicMemorySearch.scala 40:33]
  wire [2:0] c_io_target; // @[DynamicMemorySearch.scala 40:33]
  wire  c_io_done; // @[DynamicMemorySearch.scala 40:33]
  reg [6:0] value; // @[Counter.scala 17:33]
  reg  _T_6; // @[SteppedHWIOTester.scala 177:33]
  wire  _T_8 = ~_T_6; // @[SteppedHWIOTester.scala 179:10]
  wire [2:0] _GEN_9 = 7'h9 == value ? 3'h4 : 3'h5; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_10 = 7'ha == value ? 3'h4 : _GEN_9; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_11 = 7'hb == value ? 3'h4 : _GEN_10; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_12 = 7'hc == value ? 3'h4 : _GEN_11; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_13 = 7'hd == value ? 3'h4 : _GEN_12; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_14 = 7'he == value ? 3'h4 : _GEN_13; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_15 = 7'hf == value ? 3'h4 : _GEN_14; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_16 = 7'h10 == value ? 3'h4 : _GEN_15; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_17 = 7'h11 == value ? 3'h4 : _GEN_16; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_18 = 7'h12 == value ? 3'h4 : _GEN_17; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_19 = 7'h13 == value ? 3'h4 : _GEN_18; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_20 = 7'h14 == value ? 3'h4 : _GEN_19; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_21 = 7'h15 == value ? 3'h4 : _GEN_20; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_22 = 7'h16 == value ? 3'h4 : _GEN_21; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_23 = 7'h17 == value ? 3'h4 : _GEN_22; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_24 = 7'h18 == value ? 3'h4 : _GEN_23; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_25 = 7'h19 == value ? 3'h2 : _GEN_24; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_26 = 7'h1a == value ? 3'h2 : _GEN_25; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_27 = 7'h1b == value ? 3'h2 : _GEN_26; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_28 = 7'h1c == value ? 3'h2 : _GEN_27; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_29 = 7'h1d == value ? 3'h2 : _GEN_28; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_30 = 7'h1e == value ? 3'h2 : _GEN_29; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_31 = 7'h1f == value ? 3'h6 : _GEN_30; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_32 = 7'h20 == value ? 3'h6 : _GEN_31; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_33 = 7'h21 == value ? 3'h6 : _GEN_32; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_34 = 7'h22 == value ? 3'h6 : _GEN_33; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_35 = 7'h23 == value ? 3'h6 : _GEN_34; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_36 = 7'h24 == value ? 3'h6 : _GEN_35; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_37 = 7'h25 == value ? 3'h6 : _GEN_36; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_38 = 7'h26 == value ? 3'h6 : _GEN_37; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_39 = 7'h27 == value ? 3'h6 : _GEN_38; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_40 = 7'h28 == value ? 3'h6 : _GEN_39; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_41 = 7'h29 == value ? 3'h1 : _GEN_40; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_42 = 7'h2a == value ? 3'h1 : _GEN_41; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_43 = 7'h2b == value ? 3'h1 : _GEN_42; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_44 = 7'h2c == value ? 3'h1 : _GEN_43; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_45 = 7'h2d == value ? 3'h1 : _GEN_44; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_46 = 7'h2e == value ? 3'h0 : _GEN_45; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_47 = 7'h2f == value ? 3'h0 : _GEN_46; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_48 = 7'h30 == value ? 3'h0 : _GEN_47; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_49 = 7'h31 == value ? 3'h0 : _GEN_48; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_50 = 7'h32 == value ? 3'h4 : _GEN_49; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_51 = 7'h33 == value ? 3'h4 : _GEN_50; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_52 = 7'h34 == value ? 3'h4 : _GEN_51; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_53 = 7'h35 == value ? 3'h4 : _GEN_52; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_54 = 7'h36 == value ? 3'h4 : _GEN_53; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_55 = 7'h37 == value ? 3'h4 : _GEN_54; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_56 = 7'h38 == value ? 3'h4 : _GEN_55; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_57 = 7'h39 == value ? 3'h4 : _GEN_56; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_58 = 7'h3a == value ? 3'h3 : _GEN_57; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_59 = 7'h3b == value ? 3'h3 : _GEN_58; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_60 = 7'h3c == value ? 3'h3 : _GEN_59; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_61 = 7'h3d == value ? 3'h3 : _GEN_60; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_62 = 7'h3e == value ? 3'h3 : _GEN_61; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_63 = 7'h3f == value ? 3'h3 : _GEN_62; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_64 = 7'h40 == value ? 3'h3 : _GEN_63; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_65 = 7'h41 == value ? 3'h6 : _GEN_64; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_66 = 7'h42 == value ? 3'h6 : _GEN_65; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_67 = 7'h43 == value ? 3'h6 : _GEN_66; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_68 = 7'h44 == value ? 3'h6 : _GEN_67; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_69 = 7'h45 == value ? 3'h6 : _GEN_68; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_70 = 7'h46 == value ? 3'h6 : _GEN_69; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_71 = 7'h47 == value ? 3'h6 : _GEN_70; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_72 = 7'h48 == value ? 3'h6 : _GEN_71; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_73 = 7'h49 == value ? 3'h6 : _GEN_72; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_74 = 7'h4a == value ? 3'h6 : _GEN_73; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_75 = 7'h4b == value ? 3'h1 : _GEN_74; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_76 = 7'h4c == value ? 3'h1 : _GEN_75; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_77 = 7'h4d == value ? 3'h1 : _GEN_76; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_78 = 7'h4e == value ? 3'h1 : _GEN_77; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_79 = 7'h4f == value ? 3'h1 : _GEN_78; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_80 = 7'h50 == value ? 3'h3 : _GEN_79; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_81 = 7'h51 == value ? 3'h3 : _GEN_80; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_82 = 7'h52 == value ? 3'h3 : _GEN_81; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_83 = 7'h53 == value ? 3'h3 : _GEN_82; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_84 = 7'h54 == value ? 3'h3 : _GEN_83; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_85 = 7'h55 == value ? 3'h3 : _GEN_84; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_86 = 7'h56 == value ? 3'h3 : _GEN_85; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_87 = 7'h57 == value ? 3'h2 : _GEN_86; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_88 = 7'h58 == value ? 3'h2 : _GEN_87; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_89 = 7'h59 == value ? 3'h2 : _GEN_88; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_90 = 7'h5a == value ? 3'h2 : _GEN_89; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_91 = 7'h5b == value ? 3'h2 : _GEN_90; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_92 = 7'h5c == value ? 3'h2 : _GEN_91; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_93 = 7'h5d == value ? 3'h6 : _GEN_92; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_94 = 7'h5e == value ? 3'h6 : _GEN_93; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_95 = 7'h5f == value ? 3'h6 : _GEN_94; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_96 = 7'h60 == value ? 3'h6 : _GEN_95; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_97 = 7'h61 == value ? 3'h6 : _GEN_96; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_98 = 7'h62 == value ? 3'h6 : _GEN_97; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_99 = 7'h63 == value ? 3'h6 : _GEN_98; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_100 = 7'h64 == value ? 3'h6 : _GEN_99; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_101 = 7'h65 == value ? 3'h6 : _GEN_100; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_102 = 7'h66 == value ? 3'h6 : _GEN_101; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_103 = 7'h67 == value ? 3'h6 : _GEN_102; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_104 = 7'h68 == value ? 3'h6 : _GEN_103; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_105 = 7'h69 == value ? 3'h6 : _GEN_104; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_106 = 7'h6a == value ? 3'h6 : _GEN_105; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_107 = 7'h6b == value ? 3'h6 : _GEN_106; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_108 = 7'h6c == value ? 3'h2 : _GEN_107; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_109 = 7'h6d == value ? 3'h2 : _GEN_108; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_110 = 7'h6e == value ? 3'h2 : _GEN_109; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_111 = 7'h6f == value ? 3'h2 : _GEN_110; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_112 = 7'h70 == value ? 3'h2 : _GEN_111; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_113 = 7'h71 == value ? 3'h2 : _GEN_112; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_114 = 7'h72 == value ? 3'h2 : _GEN_113; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_115 = 7'h73 == value ? 3'h2 : _GEN_114; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_116 = 7'h74 == value ? 3'h2 : _GEN_115; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_117 = 7'h75 == value ? 3'h2 : _GEN_116; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [2:0] _GEN_118 = 7'h76 == value ? 3'h2 : _GEN_117; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_122 = 7'h2 == value ? 1'h0 : 7'h1 == value; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_123 = 7'h3 == value ? 1'h0 : _GEN_122; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_124 = 7'h4 == value ? 1'h0 : _GEN_123; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_125 = 7'h5 == value ? 1'h0 : _GEN_124; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_126 = 7'h6 == value ? 1'h0 : _GEN_125; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_127 = 7'h7 == value ? 1'h0 : _GEN_126; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_128 = 7'h8 == value ? 1'h0 : _GEN_127; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_129 = 7'h9 == value ? 1'h0 : _GEN_128; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_131 = 7'hb == value ? 1'h0 : 7'ha == value | _GEN_129; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_132 = 7'hc == value ? 1'h0 : _GEN_131; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_133 = 7'hd == value ? 1'h0 : _GEN_132; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_134 = 7'he == value ? 1'h0 : _GEN_133; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_135 = 7'hf == value ? 1'h0 : _GEN_134; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_136 = 7'h10 == value ? 1'h0 : _GEN_135; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_137 = 7'h11 == value ? 1'h0 : _GEN_136; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_139 = 7'h13 == value ? 1'h0 : 7'h12 == value | _GEN_137; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_140 = 7'h14 == value ? 1'h0 : _GEN_139; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_141 = 7'h15 == value ? 1'h0 : _GEN_140; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_142 = 7'h16 == value ? 1'h0 : _GEN_141; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_143 = 7'h17 == value ? 1'h0 : _GEN_142; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_144 = 7'h18 == value ? 1'h0 : _GEN_143; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_145 = 7'h19 == value ? 1'h0 : _GEN_144; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_147 = 7'h1b == value ? 1'h0 : 7'h1a == value | _GEN_145; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_148 = 7'h1c == value ? 1'h0 : _GEN_147; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_149 = 7'h1d == value ? 1'h0 : _GEN_148; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_150 = 7'h1e == value ? 1'h0 : _GEN_149; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_151 = 7'h1f == value ? 1'h0 : _GEN_150; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_153 = 7'h21 == value ? 1'h0 : 7'h20 == value | _GEN_151; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_154 = 7'h22 == value ? 1'h0 : _GEN_153; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_155 = 7'h23 == value ? 1'h0 : _GEN_154; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_156 = 7'h24 == value ? 1'h0 : _GEN_155; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_157 = 7'h25 == value ? 1'h0 : _GEN_156; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_158 = 7'h26 == value ? 1'h0 : _GEN_157; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_159 = 7'h27 == value ? 1'h0 : _GEN_158; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_160 = 7'h28 == value ? 1'h0 : _GEN_159; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_161 = 7'h29 == value ? 1'h0 : _GEN_160; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_163 = 7'h2b == value ? 1'h0 : 7'h2a == value | _GEN_161; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_164 = 7'h2c == value ? 1'h0 : _GEN_163; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_165 = 7'h2d == value ? 1'h0 : _GEN_164; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_166 = 7'h2e == value ? 1'h0 : _GEN_165; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_168 = 7'h30 == value ? 1'h0 : 7'h2f == value | _GEN_166; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_169 = 7'h31 == value ? 1'h0 : _GEN_168; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_170 = 7'h32 == value ? 1'h0 : _GEN_169; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_172 = 7'h34 == value ? 1'h0 : 7'h33 == value | _GEN_170; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_173 = 7'h35 == value ? 1'h0 : _GEN_172; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_174 = 7'h36 == value ? 1'h0 : _GEN_173; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_175 = 7'h37 == value ? 1'h0 : _GEN_174; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_176 = 7'h38 == value ? 1'h0 : _GEN_175; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_177 = 7'h39 == value ? 1'h0 : _GEN_176; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_178 = 7'h3a == value ? 1'h0 : _GEN_177; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_180 = 7'h3c == value ? 1'h0 : 7'h3b == value | _GEN_178; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_181 = 7'h3d == value ? 1'h0 : _GEN_180; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_182 = 7'h3e == value ? 1'h0 : _GEN_181; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_183 = 7'h3f == value ? 1'h0 : _GEN_182; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_184 = 7'h40 == value ? 1'h0 : _GEN_183; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_185 = 7'h41 == value ? 1'h0 : _GEN_184; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_187 = 7'h43 == value ? 1'h0 : 7'h42 == value | _GEN_185; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_188 = 7'h44 == value ? 1'h0 : _GEN_187; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_189 = 7'h45 == value ? 1'h0 : _GEN_188; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_190 = 7'h46 == value ? 1'h0 : _GEN_189; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_191 = 7'h47 == value ? 1'h0 : _GEN_190; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_192 = 7'h48 == value ? 1'h0 : _GEN_191; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_193 = 7'h49 == value ? 1'h0 : _GEN_192; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_194 = 7'h4a == value ? 1'h0 : _GEN_193; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_195 = 7'h4b == value ? 1'h0 : _GEN_194; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_197 = 7'h4d == value ? 1'h0 : 7'h4c == value | _GEN_195; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_198 = 7'h4e == value ? 1'h0 : _GEN_197; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_199 = 7'h4f == value ? 1'h0 : _GEN_198; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_200 = 7'h50 == value ? 1'h0 : _GEN_199; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_202 = 7'h52 == value ? 1'h0 : 7'h51 == value | _GEN_200; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_203 = 7'h53 == value ? 1'h0 : _GEN_202; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_204 = 7'h54 == value ? 1'h0 : _GEN_203; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_205 = 7'h55 == value ? 1'h0 : _GEN_204; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_206 = 7'h56 == value ? 1'h0 : _GEN_205; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_207 = 7'h57 == value ? 1'h0 : _GEN_206; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_209 = 7'h59 == value ? 1'h0 : 7'h58 == value | _GEN_207; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_210 = 7'h5a == value ? 1'h0 : _GEN_209; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_211 = 7'h5b == value ? 1'h0 : _GEN_210; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_212 = 7'h5c == value ? 1'h0 : _GEN_211; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_213 = 7'h5d == value ? 1'h0 : _GEN_212; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_215 = 7'h5f == value ? 1'h0 : 7'h5e == value | _GEN_213; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_216 = 7'h60 == value ? 1'h0 : _GEN_215; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_217 = 7'h61 == value ? 1'h0 : _GEN_216; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_219 = 7'h63 == value ? 1'h0 : 7'h62 == value | _GEN_217; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_220 = 7'h64 == value ? 1'h0 : _GEN_219; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_221 = 7'h65 == value ? 1'h0 : _GEN_220; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_222 = 7'h66 == value ? 1'h0 : _GEN_221; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_223 = 7'h67 == value ? 1'h0 : _GEN_222; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_224 = 7'h68 == value ? 1'h0 : _GEN_223; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_225 = 7'h69 == value ? 1'h0 : _GEN_224; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_226 = 7'h6a == value ? 1'h0 : _GEN_225; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_227 = 7'h6b == value ? 1'h0 : _GEN_226; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_228 = 7'h6c == value ? 1'h0 : _GEN_227; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_230 = 7'h6e == value ? 1'h0 : 7'h6d == value | _GEN_228; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_231 = 7'h6f == value ? 1'h0 : _GEN_230; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_232 = 7'h70 == value ? 1'h0 : _GEN_231; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_233 = 7'h71 == value ? 1'h0 : _GEN_232; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_234 = 7'h72 == value ? 1'h0 : _GEN_233; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_235 = 7'h73 == value ? 1'h0 : _GEN_234; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_236 = 7'h74 == value ? 1'h0 : _GEN_235; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_237 = 7'h75 == value ? 1'h0 : _GEN_236; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_238 = 7'h76 == value ? 1'h0 : _GEN_237; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_241 = 7'h1 == value ? 1'h0 : 1'h1; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_242 = 7'h2 == value ? 1'h0 : _GEN_241; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_243 = 7'h3 == value ? 1'h0 : _GEN_242; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_244 = 7'h4 == value ? 1'h0 : _GEN_243; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_245 = 7'h5 == value ? 1'h0 : _GEN_244; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_246 = 7'h6 == value ? 1'h0 : _GEN_245; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_247 = 7'h7 == value ? 1'h0 : _GEN_246; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_248 = 7'h8 == value ? 1'h0 : _GEN_247; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_250 = 7'ha == value ? 1'h0 : 7'h9 == value | _GEN_248; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_251 = 7'hb == value ? 1'h0 : _GEN_250; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_252 = 7'hc == value ? 1'h0 : _GEN_251; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_253 = 7'hd == value ? 1'h0 : _GEN_252; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_254 = 7'he == value ? 1'h0 : _GEN_253; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_255 = 7'hf == value ? 1'h0 : _GEN_254; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_256 = 7'h10 == value ? 1'h0 : _GEN_255; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_258 = 7'h12 == value ? 1'h0 : 7'h11 == value | _GEN_256; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_259 = 7'h13 == value ? 1'h0 : _GEN_258; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_260 = 7'h14 == value ? 1'h0 : _GEN_259; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_261 = 7'h15 == value ? 1'h0 : _GEN_260; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_262 = 7'h16 == value ? 1'h0 : _GEN_261; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_263 = 7'h17 == value ? 1'h0 : _GEN_262; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_264 = 7'h18 == value ? 1'h0 : _GEN_263; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_266 = 7'h1a == value ? 1'h0 : 7'h19 == value | _GEN_264; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_267 = 7'h1b == value ? 1'h0 : _GEN_266; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_268 = 7'h1c == value ? 1'h0 : _GEN_267; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_269 = 7'h1d == value ? 1'h0 : _GEN_268; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_270 = 7'h1e == value ? 1'h0 : _GEN_269; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_272 = 7'h20 == value ? 1'h0 : 7'h1f == value | _GEN_270; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_273 = 7'h21 == value ? 1'h0 : _GEN_272; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_274 = 7'h22 == value ? 1'h0 : _GEN_273; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_275 = 7'h23 == value ? 1'h0 : _GEN_274; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_276 = 7'h24 == value ? 1'h0 : _GEN_275; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_277 = 7'h25 == value ? 1'h0 : _GEN_276; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_278 = 7'h26 == value ? 1'h0 : _GEN_277; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_279 = 7'h27 == value ? 1'h0 : _GEN_278; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_280 = 7'h28 == value ? 1'h0 : _GEN_279; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_282 = 7'h2a == value ? 1'h0 : 7'h29 == value | _GEN_280; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_283 = 7'h2b == value ? 1'h0 : _GEN_282; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_284 = 7'h2c == value ? 1'h0 : _GEN_283; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_285 = 7'h2d == value ? 1'h0 : _GEN_284; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_287 = 7'h2f == value ? 1'h0 : 7'h2e == value | _GEN_285; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_288 = 7'h30 == value ? 1'h0 : _GEN_287; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_289 = 7'h31 == value ? 1'h0 : _GEN_288; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_291 = 7'h33 == value ? 1'h0 : 7'h32 == value | _GEN_289; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_292 = 7'h34 == value ? 1'h0 : _GEN_291; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_293 = 7'h35 == value ? 1'h0 : _GEN_292; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_294 = 7'h36 == value ? 1'h0 : _GEN_293; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_295 = 7'h37 == value ? 1'h0 : _GEN_294; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_296 = 7'h38 == value ? 1'h0 : _GEN_295; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_297 = 7'h39 == value ? 1'h0 : _GEN_296; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_299 = 7'h3b == value ? 1'h0 : 7'h3a == value | _GEN_297; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_300 = 7'h3c == value ? 1'h0 : _GEN_299; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_301 = 7'h3d == value ? 1'h0 : _GEN_300; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_302 = 7'h3e == value ? 1'h0 : _GEN_301; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_303 = 7'h3f == value ? 1'h0 : _GEN_302; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_304 = 7'h40 == value ? 1'h0 : _GEN_303; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_306 = 7'h42 == value ? 1'h0 : 7'h41 == value | _GEN_304; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_307 = 7'h43 == value ? 1'h0 : _GEN_306; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_308 = 7'h44 == value ? 1'h0 : _GEN_307; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_309 = 7'h45 == value ? 1'h0 : _GEN_308; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_310 = 7'h46 == value ? 1'h0 : _GEN_309; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_311 = 7'h47 == value ? 1'h0 : _GEN_310; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_312 = 7'h48 == value ? 1'h0 : _GEN_311; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_313 = 7'h49 == value ? 1'h0 : _GEN_312; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_314 = 7'h4a == value ? 1'h0 : _GEN_313; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_316 = 7'h4c == value ? 1'h0 : 7'h4b == value | _GEN_314; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_317 = 7'h4d == value ? 1'h0 : _GEN_316; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_318 = 7'h4e == value ? 1'h0 : _GEN_317; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_319 = 7'h4f == value ? 1'h0 : _GEN_318; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_321 = 7'h51 == value ? 1'h0 : 7'h50 == value | _GEN_319; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_322 = 7'h52 == value ? 1'h0 : _GEN_321; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_323 = 7'h53 == value ? 1'h0 : _GEN_322; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_324 = 7'h54 == value ? 1'h0 : _GEN_323; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_325 = 7'h55 == value ? 1'h0 : _GEN_324; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_326 = 7'h56 == value ? 1'h0 : _GEN_325; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_328 = 7'h58 == value ? 1'h0 : 7'h57 == value | _GEN_326; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_329 = 7'h59 == value ? 1'h0 : _GEN_328; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_330 = 7'h5a == value ? 1'h0 : _GEN_329; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_331 = 7'h5b == value ? 1'h0 : _GEN_330; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_332 = 7'h5c == value ? 1'h0 : _GEN_331; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_334 = 7'h5e == value ? 1'h0 : 7'h5d == value | _GEN_332; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_335 = 7'h5f == value ? 1'h0 : _GEN_334; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_336 = 7'h60 == value ? 1'h0 : _GEN_335; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_338 = 7'h62 == value ? 1'h0 : 7'h61 == value | _GEN_336; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_339 = 7'h63 == value ? 1'h0 : _GEN_338; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_340 = 7'h64 == value ? 1'h0 : _GEN_339; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_341 = 7'h65 == value ? 1'h0 : _GEN_340; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_342 = 7'h66 == value ? 1'h0 : _GEN_341; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_343 = 7'h67 == value ? 1'h0 : _GEN_342; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_344 = 7'h68 == value ? 1'h0 : _GEN_343; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_345 = 7'h69 == value ? 1'h0 : _GEN_344; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_346 = 7'h6a == value ? 1'h0 : _GEN_345; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_347 = 7'h6b == value ? 1'h0 : _GEN_346; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_349 = 7'h6d == value ? 1'h0 : 7'h6c == value | _GEN_347; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_350 = 7'h6e == value ? 1'h0 : _GEN_349; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_351 = 7'h6f == value ? 1'h0 : _GEN_350; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_352 = 7'h70 == value ? 1'h0 : _GEN_351; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_353 = 7'h71 == value ? 1'h0 : _GEN_352; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_354 = 7'h72 == value ? 1'h0 : _GEN_353; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_355 = 7'h73 == value ? 1'h0 : _GEN_354; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_356 = 7'h74 == value ? 1'h0 : _GEN_355; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_357 = 7'h75 == value ? 1'h0 : _GEN_356; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_358 = 7'h76 == value ? 1'h0 : _GEN_357; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_369 = 7'h9 == value ? 4'h3 : 4'he; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_370 = 7'ha == value ? 4'h3 : _GEN_369; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_371 = 7'hb == value ? 4'h3 : _GEN_370; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_372 = 7'hc == value ? 4'h3 : _GEN_371; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_373 = 7'hd == value ? 4'h3 : _GEN_372; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_374 = 7'he == value ? 4'h3 : _GEN_373; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_375 = 7'hf == value ? 4'h3 : _GEN_374; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_376 = 7'h10 == value ? 4'h3 : _GEN_375; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_377 = 7'h11 == value ? 4'h9 : _GEN_376; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_378 = 7'h12 == value ? 4'h9 : _GEN_377; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_379 = 7'h13 == value ? 4'h9 : _GEN_378; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_380 = 7'h14 == value ? 4'h9 : _GEN_379; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_381 = 7'h15 == value ? 4'h9 : _GEN_380; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_382 = 7'h16 == value ? 4'h9 : _GEN_381; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_383 = 7'h17 == value ? 4'h9 : _GEN_382; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_384 = 7'h18 == value ? 4'h9 : _GEN_383; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_385 = 7'h19 == value ? 4'h7 : _GEN_384; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_386 = 7'h1a == value ? 4'h7 : _GEN_385; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_387 = 7'h1b == value ? 4'h7 : _GEN_386; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_388 = 7'h1c == value ? 4'h7 : _GEN_387; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_389 = 7'h1d == value ? 4'h7 : _GEN_388; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_390 = 7'h1e == value ? 4'h7 : _GEN_389; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_391 = 7'h1f == value ? 4'hf : _GEN_390; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_392 = 7'h20 == value ? 4'hf : _GEN_391; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_393 = 7'h21 == value ? 4'hf : _GEN_392; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_394 = 7'h22 == value ? 4'hf : _GEN_393; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_395 = 7'h23 == value ? 4'hf : _GEN_394; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_396 = 7'h24 == value ? 4'hf : _GEN_395; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_397 = 7'h25 == value ? 4'hf : _GEN_396; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_398 = 7'h26 == value ? 4'hf : _GEN_397; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_399 = 7'h27 == value ? 4'hf : _GEN_398; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_400 = 7'h28 == value ? 4'hf : _GEN_399; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_401 = 7'h29 == value ? 4'h3 : _GEN_400; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_402 = 7'h2a == value ? 4'h3 : _GEN_401; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_403 = 7'h2b == value ? 4'h3 : _GEN_402; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_404 = 7'h2c == value ? 4'h3 : _GEN_403; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_405 = 7'h2d == value ? 4'h3 : _GEN_404; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_406 = 7'h2e == value ? 4'h8 : _GEN_405; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_407 = 7'h2f == value ? 4'h8 : _GEN_406; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_408 = 7'h30 == value ? 4'h8 : _GEN_407; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_409 = 7'h31 == value ? 4'h8 : _GEN_408; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_410 = 7'h32 == value ? 4'hf : _GEN_409; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_411 = 7'h33 == value ? 4'hf : _GEN_410; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_412 = 7'h34 == value ? 4'hf : _GEN_411; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_413 = 7'h35 == value ? 4'hf : _GEN_412; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_414 = 7'h36 == value ? 4'hf : _GEN_413; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_415 = 7'h37 == value ? 4'hf : _GEN_414; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_416 = 7'h38 == value ? 4'hf : _GEN_415; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_417 = 7'h39 == value ? 4'hf : _GEN_416; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_418 = 7'h3a == value ? 4'h1 : _GEN_417; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_419 = 7'h3b == value ? 4'h1 : _GEN_418; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_420 = 7'h3c == value ? 4'h1 : _GEN_419; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_421 = 7'h3d == value ? 4'h1 : _GEN_420; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_422 = 7'h3e == value ? 4'h1 : _GEN_421; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_423 = 7'h3f == value ? 4'h1 : _GEN_422; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_424 = 7'h40 == value ? 4'h1 : _GEN_423; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_425 = 7'h41 == value ? 4'h6 : _GEN_424; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_426 = 7'h42 == value ? 4'h6 : _GEN_425; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_427 = 7'h43 == value ? 4'h6 : _GEN_426; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_428 = 7'h44 == value ? 4'h6 : _GEN_427; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_429 = 7'h45 == value ? 4'h6 : _GEN_428; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_430 = 7'h46 == value ? 4'h6 : _GEN_429; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_431 = 7'h47 == value ? 4'h6 : _GEN_430; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_432 = 7'h48 == value ? 4'h6 : _GEN_431; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_433 = 7'h49 == value ? 4'h6 : _GEN_432; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_434 = 7'h4a == value ? 4'h6 : _GEN_433; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_435 = 7'h4b == value ? 4'h4 : _GEN_434; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_436 = 7'h4c == value ? 4'h4 : _GEN_435; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_437 = 7'h4d == value ? 4'h4 : _GEN_436; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_438 = 7'h4e == value ? 4'h4 : _GEN_437; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_439 = 7'h4f == value ? 4'h4 : _GEN_438; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_440 = 7'h50 == value ? 4'h3 : _GEN_439; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_441 = 7'h51 == value ? 4'h3 : _GEN_440; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_442 = 7'h52 == value ? 4'h3 : _GEN_441; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_443 = 7'h53 == value ? 4'h3 : _GEN_442; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_444 = 7'h54 == value ? 4'h3 : _GEN_443; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_445 = 7'h55 == value ? 4'h3 : _GEN_444; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_446 = 7'h56 == value ? 4'h3 : _GEN_445; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_447 = 7'h57 == value ? 4'hb : _GEN_446; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_448 = 7'h58 == value ? 4'hb : _GEN_447; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_449 = 7'h59 == value ? 4'hb : _GEN_448; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_450 = 7'h5a == value ? 4'hb : _GEN_449; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_451 = 7'h5b == value ? 4'hb : _GEN_450; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_452 = 7'h5c == value ? 4'hb : _GEN_451; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_453 = 7'h5d == value ? 4'h8 : _GEN_452; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_454 = 7'h5e == value ? 4'h8 : _GEN_453; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_455 = 7'h5f == value ? 4'h8 : _GEN_454; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_456 = 7'h60 == value ? 4'h8 : _GEN_455; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_457 = 7'h61 == value ? 4'h6 : _GEN_456; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_458 = 7'h62 == value ? 4'h9 : _GEN_457; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_459 = 7'h63 == value ? 4'h9 : _GEN_458; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_460 = 7'h64 == value ? 4'h9 : _GEN_459; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_461 = 7'h65 == value ? 4'h9 : _GEN_460; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_462 = 7'h66 == value ? 4'h9 : _GEN_461; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_463 = 7'h67 == value ? 4'h9 : _GEN_462; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_464 = 7'h68 == value ? 4'h9 : _GEN_463; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_465 = 7'h69 == value ? 4'h9 : _GEN_464; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_466 = 7'h6a == value ? 4'h9 : _GEN_465; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_467 = 7'h6b == value ? 4'h9 : _GEN_466; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_468 = 7'h6c == value ? 4'h3 : _GEN_467; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_469 = 7'h6d == value ? 4'ha : _GEN_468; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_470 = 7'h6e == value ? 4'ha : _GEN_469; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_471 = 7'h6f == value ? 4'ha : _GEN_470; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_472 = 7'h70 == value ? 4'ha : _GEN_471; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_473 = 7'h71 == value ? 4'ha : _GEN_472; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_474 = 7'h72 == value ? 4'ha : _GEN_473; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_475 = 7'h73 == value ? 4'ha : _GEN_474; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_476 = 7'h74 == value ? 4'ha : _GEN_475; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_477 = 7'h75 == value ? 4'ha : _GEN_476; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire [3:0] _GEN_478 = 7'h76 == value ? 4'ha : _GEN_477; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  wire  _GEN_489 = 7'h9 == value ? 1'h0 : 7'h8 == value; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_490 = 7'ha == value ? 1'h0 : _GEN_489; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_491 = 7'hb == value ? 1'h0 : _GEN_490; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_492 = 7'hc == value ? 1'h0 : _GEN_491; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_493 = 7'hd == value ? 1'h0 : _GEN_492; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_494 = 7'he == value ? 1'h0 : _GEN_493; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_495 = 7'hf == value ? 1'h0 : _GEN_494; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_497 = 7'h11 == value ? 1'h0 : 7'h10 == value | _GEN_495; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_498 = 7'h12 == value ? 1'h0 : _GEN_497; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_499 = 7'h13 == value ? 1'h0 : _GEN_498; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_500 = 7'h14 == value ? 1'h0 : _GEN_499; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_501 = 7'h15 == value ? 1'h0 : _GEN_500; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_502 = 7'h16 == value ? 1'h0 : _GEN_501; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_503 = 7'h17 == value ? 1'h0 : _GEN_502; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_505 = 7'h19 == value ? 1'h0 : 7'h18 == value | _GEN_503; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_506 = 7'h1a == value ? 1'h0 : _GEN_505; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_507 = 7'h1b == value ? 1'h0 : _GEN_506; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_508 = 7'h1c == value ? 1'h0 : _GEN_507; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_509 = 7'h1d == value ? 1'h0 : _GEN_508; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_511 = 7'h1f == value ? 1'h0 : 7'h1e == value | _GEN_509; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_512 = 7'h20 == value ? 1'h0 : _GEN_511; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_513 = 7'h21 == value ? 1'h0 : _GEN_512; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_514 = 7'h22 == value ? 1'h0 : _GEN_513; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_515 = 7'h23 == value ? 1'h0 : _GEN_514; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_516 = 7'h24 == value ? 1'h0 : _GEN_515; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_517 = 7'h25 == value ? 1'h0 : _GEN_516; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_518 = 7'h26 == value ? 1'h0 : _GEN_517; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_519 = 7'h27 == value ? 1'h0 : _GEN_518; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_521 = 7'h29 == value ? 1'h0 : 7'h28 == value | _GEN_519; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_522 = 7'h2a == value ? 1'h0 : _GEN_521; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_523 = 7'h2b == value ? 1'h0 : _GEN_522; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_524 = 7'h2c == value ? 1'h0 : _GEN_523; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_526 = 7'h2e == value ? 1'h0 : 7'h2d == value | _GEN_524; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_527 = 7'h2f == value ? 1'h0 : _GEN_526; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_528 = 7'h30 == value ? 1'h0 : _GEN_527; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_530 = 7'h32 == value ? 1'h0 : 7'h31 == value | _GEN_528; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_531 = 7'h33 == value ? 1'h0 : _GEN_530; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_532 = 7'h34 == value ? 1'h0 : _GEN_531; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_533 = 7'h35 == value ? 1'h0 : _GEN_532; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_534 = 7'h36 == value ? 1'h0 : _GEN_533; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_535 = 7'h37 == value ? 1'h0 : _GEN_534; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_536 = 7'h38 == value ? 1'h0 : _GEN_535; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_538 = 7'h3a == value ? 1'h0 : 7'h39 == value | _GEN_536; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_539 = 7'h3b == value ? 1'h0 : _GEN_538; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_540 = 7'h3c == value ? 1'h0 : _GEN_539; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_541 = 7'h3d == value ? 1'h0 : _GEN_540; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_542 = 7'h3e == value ? 1'h0 : _GEN_541; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_543 = 7'h3f == value ? 1'h0 : _GEN_542; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_545 = 7'h41 == value ? 1'h0 : 7'h40 == value | _GEN_543; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_546 = 7'h42 == value ? 1'h0 : _GEN_545; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_547 = 7'h43 == value ? 1'h0 : _GEN_546; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_548 = 7'h44 == value ? 1'h0 : _GEN_547; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_549 = 7'h45 == value ? 1'h0 : _GEN_548; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_550 = 7'h46 == value ? 1'h0 : _GEN_549; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_551 = 7'h47 == value ? 1'h0 : _GEN_550; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_552 = 7'h48 == value ? 1'h0 : _GEN_551; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_553 = 7'h49 == value ? 1'h0 : _GEN_552; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_555 = 7'h4b == value ? 1'h0 : 7'h4a == value | _GEN_553; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_556 = 7'h4c == value ? 1'h0 : _GEN_555; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_557 = 7'h4d == value ? 1'h0 : _GEN_556; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_558 = 7'h4e == value ? 1'h0 : _GEN_557; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_560 = 7'h50 == value ? 1'h0 : 7'h4f == value | _GEN_558; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_561 = 7'h51 == value ? 1'h0 : _GEN_560; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_562 = 7'h52 == value ? 1'h0 : _GEN_561; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_563 = 7'h53 == value ? 1'h0 : _GEN_562; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_564 = 7'h54 == value ? 1'h0 : _GEN_563; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_565 = 7'h55 == value ? 1'h0 : _GEN_564; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_567 = 7'h57 == value ? 1'h0 : 7'h56 == value | _GEN_565; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_568 = 7'h58 == value ? 1'h0 : _GEN_567; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_569 = 7'h59 == value ? 1'h0 : _GEN_568; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_570 = 7'h5a == value ? 1'h0 : _GEN_569; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_571 = 7'h5b == value ? 1'h0 : _GEN_570; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_573 = 7'h5d == value ? 1'h0 : 7'h5c == value | _GEN_571; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_574 = 7'h5e == value ? 1'h0 : _GEN_573; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_575 = 7'h5f == value ? 1'h0 : _GEN_574; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_577 = 7'h61 == value ? 1'h0 : 7'h60 == value | _GEN_575; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_578 = 7'h62 == value ? 1'h0 : _GEN_577; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_579 = 7'h63 == value ? 1'h0 : _GEN_578; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_580 = 7'h64 == value ? 1'h0 : _GEN_579; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_581 = 7'h65 == value ? 1'h0 : _GEN_580; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_582 = 7'h66 == value ? 1'h0 : _GEN_581; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_583 = 7'h67 == value ? 1'h0 : _GEN_582; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_584 = 7'h68 == value ? 1'h0 : _GEN_583; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_585 = 7'h69 == value ? 1'h0 : _GEN_584; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_586 = 7'h6a == value ? 1'h0 : _GEN_585; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_588 = 7'h6c == value ? 1'h0 : 7'h6b == value | _GEN_586; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_589 = 7'h6d == value ? 1'h0 : _GEN_588; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_590 = 7'h6e == value ? 1'h0 : _GEN_589; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_591 = 7'h6f == value ? 1'h0 : _GEN_590; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_592 = 7'h70 == value ? 1'h0 : _GEN_591; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_593 = 7'h71 == value ? 1'h0 : _GEN_592; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_594 = 7'h72 == value ? 1'h0 : _GEN_593; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_595 = 7'h73 == value ? 1'h0 : _GEN_594; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_596 = 7'h74 == value ? 1'h0 : _GEN_595; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_597 = 7'h75 == value ? 1'h0 : _GEN_596; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire  _GEN_599 = 7'h77 == value ? 1'h0 : 7'h76 == value | _GEN_597; // @[SteppedHWIOTester.scala 144:51 SteppedHWIOTester.scala 144:51]
  wire [2:0] _GEN_608 = 7'h8 == value ? 3'h5 : 3'h0; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_609 = 7'h9 == value ? 3'h0 : _GEN_608; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_610 = 7'ha == value ? 3'h0 : _GEN_609; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_611 = 7'hb == value ? 3'h0 : _GEN_610; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_612 = 7'hc == value ? 3'h0 : _GEN_611; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_613 = 7'hd == value ? 3'h0 : _GEN_612; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_614 = 7'he == value ? 3'h0 : _GEN_613; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_615 = 7'hf == value ? 3'h0 : _GEN_614; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_616 = 7'h10 == value ? 3'h4 : _GEN_615; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_617 = 7'h11 == value ? 3'h0 : _GEN_616; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_618 = 7'h12 == value ? 3'h0 : _GEN_617; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_619 = 7'h13 == value ? 3'h0 : _GEN_618; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_620 = 7'h14 == value ? 3'h0 : _GEN_619; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_621 = 7'h15 == value ? 3'h0 : _GEN_620; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_622 = 7'h16 == value ? 3'h0 : _GEN_621; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_623 = 7'h17 == value ? 3'h0 : _GEN_622; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_624 = 7'h18 == value ? 3'h4 : _GEN_623; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_625 = 7'h19 == value ? 3'h0 : _GEN_624; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_626 = 7'h1a == value ? 3'h0 : _GEN_625; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_627 = 7'h1b == value ? 3'h0 : _GEN_626; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_628 = 7'h1c == value ? 3'h0 : _GEN_627; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_629 = 7'h1d == value ? 3'h0 : _GEN_628; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_630 = 7'h1e == value ? 3'h2 : _GEN_629; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_631 = 7'h1f == value ? 3'h0 : _GEN_630; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_632 = 7'h20 == value ? 3'h0 : _GEN_631; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_633 = 7'h21 == value ? 3'h0 : _GEN_632; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_634 = 7'h22 == value ? 3'h0 : _GEN_633; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_635 = 7'h23 == value ? 3'h0 : _GEN_634; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_636 = 7'h24 == value ? 3'h0 : _GEN_635; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_637 = 7'h25 == value ? 3'h0 : _GEN_636; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_638 = 7'h26 == value ? 3'h0 : _GEN_637; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_639 = 7'h27 == value ? 3'h0 : _GEN_638; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_640 = 7'h28 == value ? 3'h6 : _GEN_639; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_641 = 7'h29 == value ? 3'h0 : _GEN_640; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_642 = 7'h2a == value ? 3'h0 : _GEN_641; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_643 = 7'h2b == value ? 3'h0 : _GEN_642; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_644 = 7'h2c == value ? 3'h0 : _GEN_643; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_645 = 7'h2d == value ? 3'h1 : _GEN_644; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_646 = 7'h2e == value ? 3'h0 : _GEN_645; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_647 = 7'h2f == value ? 3'h0 : _GEN_646; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_648 = 7'h30 == value ? 3'h0 : _GEN_647; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_649 = 7'h31 == value ? 3'h0 : _GEN_648; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_650 = 7'h32 == value ? 3'h0 : _GEN_649; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_651 = 7'h33 == value ? 3'h0 : _GEN_650; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_652 = 7'h34 == value ? 3'h0 : _GEN_651; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_653 = 7'h35 == value ? 3'h0 : _GEN_652; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_654 = 7'h36 == value ? 3'h0 : _GEN_653; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_655 = 7'h37 == value ? 3'h0 : _GEN_654; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_656 = 7'h38 == value ? 3'h0 : _GEN_655; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_657 = 7'h39 == value ? 3'h4 : _GEN_656; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_658 = 7'h3a == value ? 3'h0 : _GEN_657; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_659 = 7'h3b == value ? 3'h0 : _GEN_658; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_660 = 7'h3c == value ? 3'h0 : _GEN_659; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_661 = 7'h3d == value ? 3'h0 : _GEN_660; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_662 = 7'h3e == value ? 3'h0 : _GEN_661; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_663 = 7'h3f == value ? 3'h0 : _GEN_662; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_664 = 7'h40 == value ? 3'h3 : _GEN_663; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_665 = 7'h41 == value ? 3'h0 : _GEN_664; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_666 = 7'h42 == value ? 3'h0 : _GEN_665; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_667 = 7'h43 == value ? 3'h0 : _GEN_666; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_668 = 7'h44 == value ? 3'h0 : _GEN_667; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_669 = 7'h45 == value ? 3'h0 : _GEN_668; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_670 = 7'h46 == value ? 3'h0 : _GEN_669; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_671 = 7'h47 == value ? 3'h0 : _GEN_670; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_672 = 7'h48 == value ? 3'h0 : _GEN_671; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_673 = 7'h49 == value ? 3'h0 : _GEN_672; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_674 = 7'h4a == value ? 3'h6 : _GEN_673; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_675 = 7'h4b == value ? 3'h0 : _GEN_674; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_676 = 7'h4c == value ? 3'h0 : _GEN_675; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_677 = 7'h4d == value ? 3'h0 : _GEN_676; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_678 = 7'h4e == value ? 3'h0 : _GEN_677; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_679 = 7'h4f == value ? 3'h1 : _GEN_678; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_680 = 7'h50 == value ? 3'h0 : _GEN_679; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_681 = 7'h51 == value ? 3'h0 : _GEN_680; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_682 = 7'h52 == value ? 3'h0 : _GEN_681; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_683 = 7'h53 == value ? 3'h0 : _GEN_682; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_684 = 7'h54 == value ? 3'h0 : _GEN_683; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_685 = 7'h55 == value ? 3'h0 : _GEN_684; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_686 = 7'h56 == value ? 3'h3 : _GEN_685; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_687 = 7'h57 == value ? 3'h0 : _GEN_686; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_688 = 7'h58 == value ? 3'h0 : _GEN_687; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_689 = 7'h59 == value ? 3'h0 : _GEN_688; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_690 = 7'h5a == value ? 3'h0 : _GEN_689; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_691 = 7'h5b == value ? 3'h0 : _GEN_690; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_692 = 7'h5c == value ? 3'h2 : _GEN_691; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_693 = 7'h5d == value ? 3'h0 : _GEN_692; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_694 = 7'h5e == value ? 3'h0 : _GEN_693; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_695 = 7'h5f == value ? 3'h0 : _GEN_694; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_696 = 7'h60 == value ? 3'h0 : _GEN_695; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_697 = 7'h61 == value ? 3'h0 : _GEN_696; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_698 = 7'h62 == value ? 3'h0 : _GEN_697; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_699 = 7'h63 == value ? 3'h0 : _GEN_698; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_700 = 7'h64 == value ? 3'h0 : _GEN_699; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_701 = 7'h65 == value ? 3'h0 : _GEN_700; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_702 = 7'h66 == value ? 3'h0 : _GEN_701; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_703 = 7'h67 == value ? 3'h0 : _GEN_702; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_704 = 7'h68 == value ? 3'h0 : _GEN_703; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_705 = 7'h69 == value ? 3'h0 : _GEN_704; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_706 = 7'h6a == value ? 3'h0 : _GEN_705; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_707 = 7'h6b == value ? 3'h7 : _GEN_706; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_708 = 7'h6c == value ? 3'h0 : _GEN_707; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_709 = 7'h6d == value ? 3'h0 : _GEN_708; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_710 = 7'h6e == value ? 3'h0 : _GEN_709; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_711 = 7'h6f == value ? 3'h0 : _GEN_710; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_712 = 7'h70 == value ? 3'h0 : _GEN_711; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_713 = 7'h71 == value ? 3'h0 : _GEN_712; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_714 = 7'h72 == value ? 3'h0 : _GEN_713; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_715 = 7'h73 == value ? 3'h0 : _GEN_714; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_716 = 7'h74 == value ? 3'h0 : _GEN_715; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_717 = 7'h75 == value ? 3'h0 : _GEN_716; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_718 = 7'h76 == value ? 3'h7 : _GEN_717; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire [2:0] _GEN_719 = 7'h77 == value ? 3'h0 : _GEN_718; // @[SteppedHWIOTester.scala 145:31 SteppedHWIOTester.scala 145:31]
  wire  _T_1845 = c_io_target == _GEN_719; // @[SteppedHWIOTester.scala 145:31]
  wire  _T_1847 = ~reset; // @[HWIOTester.scala 30:55]
  wire  _T_1849 = ~(c_io_target == _GEN_719); // @[SteppedHWIOTester.scala 145:72]
  wire  _T_2711 = c_io_done == _GEN_599; // @[SteppedHWIOTester.scala 145:31]
  wire  _T_2715 = ~(c_io_done == _GEN_599); // @[SteppedHWIOTester.scala 145:72]
  wire  _T_2726 = value == 7'h77; // @[Counter.scala 25:24]
  wire [6:0] _T_2729 = value + 7'h1; // @[Counter.scala 26:22]
  wire  _GEN_961 = _T_2726 | _T_6; // @[SteppedHWIOTester.scala 183:22 SteppedHWIOTester.scala 185:14 SteppedHWIOTester.scala 177:33]
  wire  _GEN_1043 = _T_8 & _GEN_599; // @[HWIOTester.scala 30:55]
  wire  _GEN_1046 = _GEN_1043 & _T_1849; // @[SteppedHWIOTester.scala 151:15]
  wire  _GEN_1056 = _GEN_1043 & _T_2715; // @[SteppedHWIOTester.scala 151:15]
  wire  _GEN_1063 = _T_8 & _T_2726; // @[SteppedHWIOTester.scala 184:15]
  DynamicMemorySearch c ( // @[DynamicMemorySearch.scala 40:33]
    .clock(c_clock),
    .reset(c_reset),
    .io_isWr(c_io_isWr),
    .io_wrAddr(c_io_wrAddr),
    .io_data(c_io_data),
    .io_en(c_io_en),
    .io_target(c_io_target),
    .io_done(c_io_done)
  );
  assign c_clock = clock;
  assign c_reset = reset;
  assign c_io_isWr = 7'h77 == value ? 1'h0 : _GEN_358; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  assign c_io_wrAddr = 7'h77 == value ? 3'h2 : _GEN_118; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  assign c_io_data = 7'h77 == value ? 4'ha : _GEN_478; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  assign c_io_en = 7'h77 == value ? 1'h0 : _GEN_238; // @[SteppedHWIOTester.scala 129:16 SteppedHWIOTester.scala 129:16]
  always @(posedge clock) begin
    if (reset) begin // @[Counter.scala 17:33]
      value <= 7'h0; // @[Counter.scala 17:33]
    end else if (~_T_6) begin // @[SteppedHWIOTester.scala 179:17]
      if (_T_2726) begin // @[Counter.scala 28:21]
        value <= 7'h0; // @[Counter.scala 28:29]
      end else begin
        value <= _T_2729; // @[Counter.scala 26:13]
      end
    end
    if (reset) begin // @[SteppedHWIOTester.scala 177:33]
      _T_6 <= 1'h0; // @[SteppedHWIOTester.scala 177:33]
    end else if (~_T_6) begin // @[SteppedHWIOTester.scala 179:17]
      _T_6 <= _GEN_961;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8 & _GEN_599 & _T_1845 & ~reset) begin
          $fwrite(32'h80000002,"    passed step %d -- target:  %d\n",value,c_io_target); // @[HWIOTester.scala 30:55]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_1043 & _T_1849 & _T_1847) begin
          $fwrite(32'h80000002,"    failed on step %d -- port target:  %d expected %d\n",value,c_io_target,_GEN_719); // @[SteppedHWIOTester.scala 151:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_1046 & _T_1847) begin
          $fwrite(32'h80000002,"Assertion failed\n    at SteppedHWIOTester.scala:158 assert(false.B)\n"); // @[SteppedHWIOTester.scala 158:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_1046 & _T_1847) begin
          $fatal; // @[SteppedHWIOTester.scala 158:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_1046 & _T_1847) begin
          $finish; // @[SteppedHWIOTester.scala 159:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8 & _GEN_599 & _T_2711 & ~reset) begin
          $fwrite(32'h80000002,"    passed step %d -- done:  %d\n",value,c_io_done); // @[HWIOTester.scala 30:55]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_1043 & _T_2715 & _T_1847) begin
          $fwrite(32'h80000002,"    failed on step %d -- port done:  %d expected %d\n",value,c_io_done,_GEN_599); // @[SteppedHWIOTester.scala 151:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_1056 & _T_1847) begin
          $fwrite(32'h80000002,"Assertion failed\n    at SteppedHWIOTester.scala:158 assert(false.B)\n"); // @[SteppedHWIOTester.scala 158:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_1056 & _T_1847) begin
          $fatal; // @[SteppedHWIOTester.scala 158:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_1056 & _T_1847) begin
          $finish; // @[SteppedHWIOTester.scala 159:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8 & _T_2726 & _T_1847) begin
          $fwrite(32'h80000002,"Stopping, end of tests, 120 steps\n"); // @[SteppedHWIOTester.scala 184:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_1063 & _T_1847) begin
          $finish; // @[SteppedHWIOTester.scala 186:13]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[6:0];
  _RAND_1 = {1{`RANDOM}};
  _T_6 = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
