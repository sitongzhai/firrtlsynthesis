module MaxNTests(
    input clock,
    input reset
);
    wire _c__clock;
    wire _c__reset;
    wire [15:0] _c__io_ins_0;
    wire [15:0] _c__io_ins_1;
    wire [15:0] _c__io_ins_2;
    wire [15:0] _c__io_ins_3;
    wire [15:0] _c__io_ins_4;
    wire [15:0] _c__io_ins_5;
    wire [15:0] _c__io_ins_6;
    wire [15:0] _c__io_ins_7;
    wire [15:0] _c__io_ins_8;
    wire [15:0] _c__io_ins_9;
    wire [15:0] _c__io_out;
    MaxN c (
        .clock(_c__clock),
        .reset(_c__reset),
        .io_ins_0(_c__io_ins_0),
        .io_ins_1(_c__io_ins_1),
        .io_ins_2(_c__io_ins_2),
        .io_ins_3(_c__io_ins_3),
        .io_ins_4(_c__io_ins_4),
        .io_ins_5(_c__io_ins_5),
        .io_ins_6(_c__io_ins_6),
        .io_ins_7(_c__io_ins_7),
        .io_ins_8(_c__io_ins_8),
        .io_ins_9(_c__io_ins_9),
        .io_out(_c__io_out)
    );
    wire [3:0] _value__q;
    wire [3:0] _value__d;
    DFF_POSCLK #(.width(4)) value (
        .q(_value__q),
        .d(_value__d),
        .clk(clock)
    );
    wire [3:0] _WTEMP_0;
    MUX_UNSIGNED #(.width(4)) u_mux_19 (
        .y(_value__d),
        .sel(reset),
        .a(4'h0),
        .b(_WTEMP_0)
    );
    wire __T_6__q;
    wire __T_6__d;
    DFF_POSCLK #(.width(1)) _T_6 (
        .q(__T_6__q),
        .d(__T_6__d),
        .clk(clock)
    );
    wire _WTEMP_1;
    MUX_UNSIGNED #(.width(1)) u_mux_20 (
        .y(__T_6__d),
        .sel(reset),
        .a(1'h0),
        .b(_WTEMP_1)
    );
    wire _T_8;
    EQ_UNSIGNED #(.width(1)) u_eq_21 (
        .y(_T_8),
        .a(__T_6__q),
        .b(1'h0)
    );
    wire [15:0] _T_22_0;
    wire [15:0] _T_22_1;
    wire [15:0] _T_22_2;
    wire [15:0] _T_22_3;
    wire [15:0] _T_22_4;
    wire [15:0] _T_22_5;
    wire [15:0] _T_22_6;
    wire [15:0] _T_22_7;
    wire [15:0] _T_22_8;
    wire [15:0] _T_22_9;
    wire [15:0] _T_22_10;
    wire _node_0;
    EQ_UNSIGNED #(.width(4)) u_eq_22 (
        .y(_node_0),
        .a(4'd0),
        .b(_value__q)
    );
    wire [15:0] _node_1;
    assign _node_1 = _T_22_0;
    wire _node_2;
    EQ_UNSIGNED #(.width(4)) u_eq_23 (
        .y(_node_2),
        .a(4'd1),
        .b(_value__q)
    );
    wire [15:0] _node_3;
    MUX_UNSIGNED #(.width(16)) u_mux_24 (
        .y(_node_3),
        .sel(_node_2),
        .a(_T_22_1),
        .b(_node_1)
    );
    wire _node_4;
    EQ_UNSIGNED #(.width(4)) u_eq_25 (
        .y(_node_4),
        .a(4'd2),
        .b(_value__q)
    );
    wire [15:0] _node_5;
    MUX_UNSIGNED #(.width(16)) u_mux_26 (
        .y(_node_5),
        .sel(_node_4),
        .a(_T_22_2),
        .b(_node_3)
    );
    wire _node_6;
    EQ_UNSIGNED #(.width(4)) u_eq_27 (
        .y(_node_6),
        .a(4'd3),
        .b(_value__q)
    );
    wire [15:0] _node_7;
    MUX_UNSIGNED #(.width(16)) u_mux_28 (
        .y(_node_7),
        .sel(_node_6),
        .a(_T_22_3),
        .b(_node_5)
    );
    wire _node_8;
    EQ_UNSIGNED #(.width(4)) u_eq_29 (
        .y(_node_8),
        .a(4'd4),
        .b(_value__q)
    );
    wire [15:0] _node_9;
    MUX_UNSIGNED #(.width(16)) u_mux_30 (
        .y(_node_9),
        .sel(_node_8),
        .a(_T_22_4),
        .b(_node_7)
    );
    wire _node_10;
    EQ_UNSIGNED #(.width(4)) u_eq_31 (
        .y(_node_10),
        .a(4'd5),
        .b(_value__q)
    );
    wire [15:0] _node_11;
    MUX_UNSIGNED #(.width(16)) u_mux_32 (
        .y(_node_11),
        .sel(_node_10),
        .a(_T_22_5),
        .b(_node_9)
    );
    wire _node_12;
    EQ_UNSIGNED #(.width(4)) u_eq_33 (
        .y(_node_12),
        .a(4'd6),
        .b(_value__q)
    );
    wire [15:0] _node_13;
    MUX_UNSIGNED #(.width(16)) u_mux_34 (
        .y(_node_13),
        .sel(_node_12),
        .a(_T_22_6),
        .b(_node_11)
    );
    wire _node_14;
    EQ_UNSIGNED #(.width(4)) u_eq_35 (
        .y(_node_14),
        .a(4'd7),
        .b(_value__q)
    );
    wire [15:0] _node_15;
    MUX_UNSIGNED #(.width(16)) u_mux_36 (
        .y(_node_15),
        .sel(_node_14),
        .a(_T_22_7),
        .b(_node_13)
    );
    wire _node_16;
    EQ_UNSIGNED #(.width(4)) u_eq_37 (
        .y(_node_16),
        .a(4'd8),
        .b(_value__q)
    );
    wire [15:0] _node_17;
    MUX_UNSIGNED #(.width(16)) u_mux_38 (
        .y(_node_17),
        .sel(_node_16),
        .a(_T_22_8),
        .b(_node_15)
    );
    wire _node_18;
    EQ_UNSIGNED #(.width(4)) u_eq_39 (
        .y(_node_18),
        .a(4'd9),
        .b(_value__q)
    );
    wire [15:0] _node_19;
    MUX_UNSIGNED #(.width(16)) u_mux_40 (
        .y(_node_19),
        .sel(_node_18),
        .a(_T_22_9),
        .b(_node_17)
    );
    wire _node_20;
    EQ_UNSIGNED #(.width(4)) u_eq_41 (
        .y(_node_20),
        .a(4'd10),
        .b(_value__q)
    );
    wire [15:0] _node_21;
    MUX_UNSIGNED #(.width(16)) u_mux_42 (
        .y(_node_21),
        .sel(_node_20),
        .a(_T_22_10),
        .b(_node_19)
    );
    wire [15:0] _T_50_0;
    wire [15:0] _T_50_1;
    wire [15:0] _T_50_2;
    wire [15:0] _T_50_3;
    wire [15:0] _T_50_4;
    wire [15:0] _T_50_5;
    wire [15:0] _T_50_6;
    wire [15:0] _T_50_7;
    wire [15:0] _T_50_8;
    wire [15:0] _T_50_9;
    wire [15:0] _T_50_10;
    wire _node_22;
    EQ_UNSIGNED #(.width(4)) u_eq_43 (
        .y(_node_22),
        .a(4'd0),
        .b(_value__q)
    );
    wire [15:0] _node_23;
    assign _node_23 = _T_50_0;
    wire _node_24;
    EQ_UNSIGNED #(.width(4)) u_eq_44 (
        .y(_node_24),
        .a(4'd1),
        .b(_value__q)
    );
    wire [15:0] _node_25;
    MUX_UNSIGNED #(.width(16)) u_mux_45 (
        .y(_node_25),
        .sel(_node_24),
        .a(_T_50_1),
        .b(_node_23)
    );
    wire _node_26;
    EQ_UNSIGNED #(.width(4)) u_eq_46 (
        .y(_node_26),
        .a(4'd2),
        .b(_value__q)
    );
    wire [15:0] _node_27;
    MUX_UNSIGNED #(.width(16)) u_mux_47 (
        .y(_node_27),
        .sel(_node_26),
        .a(_T_50_2),
        .b(_node_25)
    );
    wire _node_28;
    EQ_UNSIGNED #(.width(4)) u_eq_48 (
        .y(_node_28),
        .a(4'd3),
        .b(_value__q)
    );
    wire [15:0] _node_29;
    MUX_UNSIGNED #(.width(16)) u_mux_49 (
        .y(_node_29),
        .sel(_node_28),
        .a(_T_50_3),
        .b(_node_27)
    );
    wire _node_30;
    EQ_UNSIGNED #(.width(4)) u_eq_50 (
        .y(_node_30),
        .a(4'd4),
        .b(_value__q)
    );
    wire [15:0] _node_31;
    MUX_UNSIGNED #(.width(16)) u_mux_51 (
        .y(_node_31),
        .sel(_node_30),
        .a(_T_50_4),
        .b(_node_29)
    );
    wire _node_32;
    EQ_UNSIGNED #(.width(4)) u_eq_52 (
        .y(_node_32),
        .a(4'd5),
        .b(_value__q)
    );
    wire [15:0] _node_33;
    MUX_UNSIGNED #(.width(16)) u_mux_53 (
        .y(_node_33),
        .sel(_node_32),
        .a(_T_50_5),
        .b(_node_31)
    );
    wire _node_34;
    EQ_UNSIGNED #(.width(4)) u_eq_54 (
        .y(_node_34),
        .a(4'd6),
        .b(_value__q)
    );
    wire [15:0] _node_35;
    MUX_UNSIGNED #(.width(16)) u_mux_55 (
        .y(_node_35),
        .sel(_node_34),
        .a(_T_50_6),
        .b(_node_33)
    );
    wire _node_36;
    EQ_UNSIGNED #(.width(4)) u_eq_56 (
        .y(_node_36),
        .a(4'd7),
        .b(_value__q)
    );
    wire [15:0] _node_37;
    MUX_UNSIGNED #(.width(16)) u_mux_57 (
        .y(_node_37),
        .sel(_node_36),
        .a(_T_50_7),
        .b(_node_35)
    );
    wire _node_38;
    EQ_UNSIGNED #(.width(4)) u_eq_58 (
        .y(_node_38),
        .a(4'd8),
        .b(_value__q)
    );
    wire [15:0] _node_39;
    MUX_UNSIGNED #(.width(16)) u_mux_59 (
        .y(_node_39),
        .sel(_node_38),
        .a(_T_50_8),
        .b(_node_37)
    );
    wire _node_40;
    EQ_UNSIGNED #(.width(4)) u_eq_60 (
        .y(_node_40),
        .a(4'd9),
        .b(_value__q)
    );
    wire [15:0] _node_41;
    MUX_UNSIGNED #(.width(16)) u_mux_61 (
        .y(_node_41),
        .sel(_node_40),
        .a(_T_50_9),
        .b(_node_39)
    );
    wire _node_42;
    EQ_UNSIGNED #(.width(4)) u_eq_62 (
        .y(_node_42),
        .a(4'd10),
        .b(_value__q)
    );
    wire [15:0] _node_43;
    MUX_UNSIGNED #(.width(16)) u_mux_63 (
        .y(_node_43),
        .sel(_node_42),
        .a(_T_50_10),
        .b(_node_41)
    );
    wire [15:0] _T_78_0;
    wire [15:0] _T_78_1;
    wire [15:0] _T_78_2;
    wire [15:0] _T_78_3;
    wire [15:0] _T_78_4;
    wire [15:0] _T_78_5;
    wire [15:0] _T_78_6;
    wire [15:0] _T_78_7;
    wire [15:0] _T_78_8;
    wire [15:0] _T_78_9;
    wire [15:0] _T_78_10;
    wire _node_44;
    EQ_UNSIGNED #(.width(4)) u_eq_64 (
        .y(_node_44),
        .a(4'd0),
        .b(_value__q)
    );
    wire [15:0] _node_45;
    assign _node_45 = _T_78_0;
    wire _node_46;
    EQ_UNSIGNED #(.width(4)) u_eq_65 (
        .y(_node_46),
        .a(4'd1),
        .b(_value__q)
    );
    wire [15:0] _node_47;
    MUX_UNSIGNED #(.width(16)) u_mux_66 (
        .y(_node_47),
        .sel(_node_46),
        .a(_T_78_1),
        .b(_node_45)
    );
    wire _node_48;
    EQ_UNSIGNED #(.width(4)) u_eq_67 (
        .y(_node_48),
        .a(4'd2),
        .b(_value__q)
    );
    wire [15:0] _node_49;
    MUX_UNSIGNED #(.width(16)) u_mux_68 (
        .y(_node_49),
        .sel(_node_48),
        .a(_T_78_2),
        .b(_node_47)
    );
    wire _node_50;
    EQ_UNSIGNED #(.width(4)) u_eq_69 (
        .y(_node_50),
        .a(4'd3),
        .b(_value__q)
    );
    wire [15:0] _node_51;
    MUX_UNSIGNED #(.width(16)) u_mux_70 (
        .y(_node_51),
        .sel(_node_50),
        .a(_T_78_3),
        .b(_node_49)
    );
    wire _node_52;
    EQ_UNSIGNED #(.width(4)) u_eq_71 (
        .y(_node_52),
        .a(4'd4),
        .b(_value__q)
    );
    wire [15:0] _node_53;
    MUX_UNSIGNED #(.width(16)) u_mux_72 (
        .y(_node_53),
        .sel(_node_52),
        .a(_T_78_4),
        .b(_node_51)
    );
    wire _node_54;
    EQ_UNSIGNED #(.width(4)) u_eq_73 (
        .y(_node_54),
        .a(4'd5),
        .b(_value__q)
    );
    wire [15:0] _node_55;
    MUX_UNSIGNED #(.width(16)) u_mux_74 (
        .y(_node_55),
        .sel(_node_54),
        .a(_T_78_5),
        .b(_node_53)
    );
    wire _node_56;
    EQ_UNSIGNED #(.width(4)) u_eq_75 (
        .y(_node_56),
        .a(4'd6),
        .b(_value__q)
    );
    wire [15:0] _node_57;
    MUX_UNSIGNED #(.width(16)) u_mux_76 (
        .y(_node_57),
        .sel(_node_56),
        .a(_T_78_6),
        .b(_node_55)
    );
    wire _node_58;
    EQ_UNSIGNED #(.width(4)) u_eq_77 (
        .y(_node_58),
        .a(4'd7),
        .b(_value__q)
    );
    wire [15:0] _node_59;
    MUX_UNSIGNED #(.width(16)) u_mux_78 (
        .y(_node_59),
        .sel(_node_58),
        .a(_T_78_7),
        .b(_node_57)
    );
    wire _node_60;
    EQ_UNSIGNED #(.width(4)) u_eq_79 (
        .y(_node_60),
        .a(4'd8),
        .b(_value__q)
    );
    wire [15:0] _node_61;
    MUX_UNSIGNED #(.width(16)) u_mux_80 (
        .y(_node_61),
        .sel(_node_60),
        .a(_T_78_8),
        .b(_node_59)
    );
    wire _node_62;
    EQ_UNSIGNED #(.width(4)) u_eq_81 (
        .y(_node_62),
        .a(4'd9),
        .b(_value__q)
    );
    wire [15:0] _node_63;
    MUX_UNSIGNED #(.width(16)) u_mux_82 (
        .y(_node_63),
        .sel(_node_62),
        .a(_T_78_9),
        .b(_node_61)
    );
    wire _node_64;
    EQ_UNSIGNED #(.width(4)) u_eq_83 (
        .y(_node_64),
        .a(4'd10),
        .b(_value__q)
    );
    wire [15:0] _node_65;
    MUX_UNSIGNED #(.width(16)) u_mux_84 (
        .y(_node_65),
        .sel(_node_64),
        .a(_T_78_10),
        .b(_node_63)
    );
    wire [15:0] _T_106_0;
    wire [15:0] _T_106_1;
    wire [15:0] _T_106_2;
    wire [15:0] _T_106_3;
    wire [15:0] _T_106_4;
    wire [15:0] _T_106_5;
    wire [15:0] _T_106_6;
    wire [15:0] _T_106_7;
    wire [15:0] _T_106_8;
    wire [15:0] _T_106_9;
    wire [15:0] _T_106_10;
    wire _node_66;
    EQ_UNSIGNED #(.width(4)) u_eq_85 (
        .y(_node_66),
        .a(4'd0),
        .b(_value__q)
    );
    wire [15:0] _node_67;
    assign _node_67 = _T_106_0;
    wire _node_68;
    EQ_UNSIGNED #(.width(4)) u_eq_86 (
        .y(_node_68),
        .a(4'd1),
        .b(_value__q)
    );
    wire [15:0] _node_69;
    MUX_UNSIGNED #(.width(16)) u_mux_87 (
        .y(_node_69),
        .sel(_node_68),
        .a(_T_106_1),
        .b(_node_67)
    );
    wire _node_70;
    EQ_UNSIGNED #(.width(4)) u_eq_88 (
        .y(_node_70),
        .a(4'd2),
        .b(_value__q)
    );
    wire [15:0] _node_71;
    MUX_UNSIGNED #(.width(16)) u_mux_89 (
        .y(_node_71),
        .sel(_node_70),
        .a(_T_106_2),
        .b(_node_69)
    );
    wire _node_72;
    EQ_UNSIGNED #(.width(4)) u_eq_90 (
        .y(_node_72),
        .a(4'd3),
        .b(_value__q)
    );
    wire [15:0] _node_73;
    MUX_UNSIGNED #(.width(16)) u_mux_91 (
        .y(_node_73),
        .sel(_node_72),
        .a(_T_106_3),
        .b(_node_71)
    );
    wire _node_74;
    EQ_UNSIGNED #(.width(4)) u_eq_92 (
        .y(_node_74),
        .a(4'd4),
        .b(_value__q)
    );
    wire [15:0] _node_75;
    MUX_UNSIGNED #(.width(16)) u_mux_93 (
        .y(_node_75),
        .sel(_node_74),
        .a(_T_106_4),
        .b(_node_73)
    );
    wire _node_76;
    EQ_UNSIGNED #(.width(4)) u_eq_94 (
        .y(_node_76),
        .a(4'd5),
        .b(_value__q)
    );
    wire [15:0] _node_77;
    MUX_UNSIGNED #(.width(16)) u_mux_95 (
        .y(_node_77),
        .sel(_node_76),
        .a(_T_106_5),
        .b(_node_75)
    );
    wire _node_78;
    EQ_UNSIGNED #(.width(4)) u_eq_96 (
        .y(_node_78),
        .a(4'd6),
        .b(_value__q)
    );
    wire [15:0] _node_79;
    MUX_UNSIGNED #(.width(16)) u_mux_97 (
        .y(_node_79),
        .sel(_node_78),
        .a(_T_106_6),
        .b(_node_77)
    );
    wire _node_80;
    EQ_UNSIGNED #(.width(4)) u_eq_98 (
        .y(_node_80),
        .a(4'd7),
        .b(_value__q)
    );
    wire [15:0] _node_81;
    MUX_UNSIGNED #(.width(16)) u_mux_99 (
        .y(_node_81),
        .sel(_node_80),
        .a(_T_106_7),
        .b(_node_79)
    );
    wire _node_82;
    EQ_UNSIGNED #(.width(4)) u_eq_100 (
        .y(_node_82),
        .a(4'd8),
        .b(_value__q)
    );
    wire [15:0] _node_83;
    MUX_UNSIGNED #(.width(16)) u_mux_101 (
        .y(_node_83),
        .sel(_node_82),
        .a(_T_106_8),
        .b(_node_81)
    );
    wire _node_84;
    EQ_UNSIGNED #(.width(4)) u_eq_102 (
        .y(_node_84),
        .a(4'd9),
        .b(_value__q)
    );
    wire [15:0] _node_85;
    MUX_UNSIGNED #(.width(16)) u_mux_103 (
        .y(_node_85),
        .sel(_node_84),
        .a(_T_106_9),
        .b(_node_83)
    );
    wire _node_86;
    EQ_UNSIGNED #(.width(4)) u_eq_104 (
        .y(_node_86),
        .a(4'd10),
        .b(_value__q)
    );
    wire [15:0] _node_87;
    MUX_UNSIGNED #(.width(16)) u_mux_105 (
        .y(_node_87),
        .sel(_node_86),
        .a(_T_106_10),
        .b(_node_85)
    );
    wire [15:0] _T_134_0;
    wire [15:0] _T_134_1;
    wire [15:0] _T_134_2;
    wire [15:0] _T_134_3;
    wire [15:0] _T_134_4;
    wire [15:0] _T_134_5;
    wire [15:0] _T_134_6;
    wire [15:0] _T_134_7;
    wire [15:0] _T_134_8;
    wire [15:0] _T_134_9;
    wire [15:0] _T_134_10;
    wire _node_88;
    EQ_UNSIGNED #(.width(4)) u_eq_106 (
        .y(_node_88),
        .a(4'd0),
        .b(_value__q)
    );
    wire [15:0] _node_89;
    assign _node_89 = _T_134_0;
    wire _node_90;
    EQ_UNSIGNED #(.width(4)) u_eq_107 (
        .y(_node_90),
        .a(4'd1),
        .b(_value__q)
    );
    wire [15:0] _node_91;
    MUX_UNSIGNED #(.width(16)) u_mux_108 (
        .y(_node_91),
        .sel(_node_90),
        .a(_T_134_1),
        .b(_node_89)
    );
    wire _node_92;
    EQ_UNSIGNED #(.width(4)) u_eq_109 (
        .y(_node_92),
        .a(4'd2),
        .b(_value__q)
    );
    wire [15:0] _node_93;
    MUX_UNSIGNED #(.width(16)) u_mux_110 (
        .y(_node_93),
        .sel(_node_92),
        .a(_T_134_2),
        .b(_node_91)
    );
    wire _node_94;
    EQ_UNSIGNED #(.width(4)) u_eq_111 (
        .y(_node_94),
        .a(4'd3),
        .b(_value__q)
    );
    wire [15:0] _node_95;
    MUX_UNSIGNED #(.width(16)) u_mux_112 (
        .y(_node_95),
        .sel(_node_94),
        .a(_T_134_3),
        .b(_node_93)
    );
    wire _node_96;
    EQ_UNSIGNED #(.width(4)) u_eq_113 (
        .y(_node_96),
        .a(4'd4),
        .b(_value__q)
    );
    wire [15:0] _node_97;
    MUX_UNSIGNED #(.width(16)) u_mux_114 (
        .y(_node_97),
        .sel(_node_96),
        .a(_T_134_4),
        .b(_node_95)
    );
    wire _node_98;
    EQ_UNSIGNED #(.width(4)) u_eq_115 (
        .y(_node_98),
        .a(4'd5),
        .b(_value__q)
    );
    wire [15:0] _node_99;
    MUX_UNSIGNED #(.width(16)) u_mux_116 (
        .y(_node_99),
        .sel(_node_98),
        .a(_T_134_5),
        .b(_node_97)
    );
    wire _node_100;
    EQ_UNSIGNED #(.width(4)) u_eq_117 (
        .y(_node_100),
        .a(4'd6),
        .b(_value__q)
    );
    wire [15:0] _node_101;
    MUX_UNSIGNED #(.width(16)) u_mux_118 (
        .y(_node_101),
        .sel(_node_100),
        .a(_T_134_6),
        .b(_node_99)
    );
    wire _node_102;
    EQ_UNSIGNED #(.width(4)) u_eq_119 (
        .y(_node_102),
        .a(4'd7),
        .b(_value__q)
    );
    wire [15:0] _node_103;
    MUX_UNSIGNED #(.width(16)) u_mux_120 (
        .y(_node_103),
        .sel(_node_102),
        .a(_T_134_7),
        .b(_node_101)
    );
    wire _node_104;
    EQ_UNSIGNED #(.width(4)) u_eq_121 (
        .y(_node_104),
        .a(4'd8),
        .b(_value__q)
    );
    wire [15:0] _node_105;
    MUX_UNSIGNED #(.width(16)) u_mux_122 (
        .y(_node_105),
        .sel(_node_104),
        .a(_T_134_8),
        .b(_node_103)
    );
    wire _node_106;
    EQ_UNSIGNED #(.width(4)) u_eq_123 (
        .y(_node_106),
        .a(4'd9),
        .b(_value__q)
    );
    wire [15:0] _node_107;
    MUX_UNSIGNED #(.width(16)) u_mux_124 (
        .y(_node_107),
        .sel(_node_106),
        .a(_T_134_9),
        .b(_node_105)
    );
    wire _node_108;
    EQ_UNSIGNED #(.width(4)) u_eq_125 (
        .y(_node_108),
        .a(4'd10),
        .b(_value__q)
    );
    wire [15:0] _node_109;
    MUX_UNSIGNED #(.width(16)) u_mux_126 (
        .y(_node_109),
        .sel(_node_108),
        .a(_T_134_10),
        .b(_node_107)
    );
    wire [15:0] _T_162_0;
    wire [15:0] _T_162_1;
    wire [15:0] _T_162_2;
    wire [15:0] _T_162_3;
    wire [15:0] _T_162_4;
    wire [15:0] _T_162_5;
    wire [15:0] _T_162_6;
    wire [15:0] _T_162_7;
    wire [15:0] _T_162_8;
    wire [15:0] _T_162_9;
    wire [15:0] _T_162_10;
    wire _node_110;
    EQ_UNSIGNED #(.width(4)) u_eq_127 (
        .y(_node_110),
        .a(4'd0),
        .b(_value__q)
    );
    wire [15:0] _node_111;
    assign _node_111 = _T_162_0;
    wire _node_112;
    EQ_UNSIGNED #(.width(4)) u_eq_128 (
        .y(_node_112),
        .a(4'd1),
        .b(_value__q)
    );
    wire [15:0] _node_113;
    MUX_UNSIGNED #(.width(16)) u_mux_129 (
        .y(_node_113),
        .sel(_node_112),
        .a(_T_162_1),
        .b(_node_111)
    );
    wire _node_114;
    EQ_UNSIGNED #(.width(4)) u_eq_130 (
        .y(_node_114),
        .a(4'd2),
        .b(_value__q)
    );
    wire [15:0] _node_115;
    MUX_UNSIGNED #(.width(16)) u_mux_131 (
        .y(_node_115),
        .sel(_node_114),
        .a(_T_162_2),
        .b(_node_113)
    );
    wire _node_116;
    EQ_UNSIGNED #(.width(4)) u_eq_132 (
        .y(_node_116),
        .a(4'd3),
        .b(_value__q)
    );
    wire [15:0] _node_117;
    MUX_UNSIGNED #(.width(16)) u_mux_133 (
        .y(_node_117),
        .sel(_node_116),
        .a(_T_162_3),
        .b(_node_115)
    );
    wire _node_118;
    EQ_UNSIGNED #(.width(4)) u_eq_134 (
        .y(_node_118),
        .a(4'd4),
        .b(_value__q)
    );
    wire [15:0] _node_119;
    MUX_UNSIGNED #(.width(16)) u_mux_135 (
        .y(_node_119),
        .sel(_node_118),
        .a(_T_162_4),
        .b(_node_117)
    );
    wire _node_120;
    EQ_UNSIGNED #(.width(4)) u_eq_136 (
        .y(_node_120),
        .a(4'd5),
        .b(_value__q)
    );
    wire [15:0] _node_121;
    MUX_UNSIGNED #(.width(16)) u_mux_137 (
        .y(_node_121),
        .sel(_node_120),
        .a(_T_162_5),
        .b(_node_119)
    );
    wire _node_122;
    EQ_UNSIGNED #(.width(4)) u_eq_138 (
        .y(_node_122),
        .a(4'd6),
        .b(_value__q)
    );
    wire [15:0] _node_123;
    MUX_UNSIGNED #(.width(16)) u_mux_139 (
        .y(_node_123),
        .sel(_node_122),
        .a(_T_162_6),
        .b(_node_121)
    );
    wire _node_124;
    EQ_UNSIGNED #(.width(4)) u_eq_140 (
        .y(_node_124),
        .a(4'd7),
        .b(_value__q)
    );
    wire [15:0] _node_125;
    MUX_UNSIGNED #(.width(16)) u_mux_141 (
        .y(_node_125),
        .sel(_node_124),
        .a(_T_162_7),
        .b(_node_123)
    );
    wire _node_126;
    EQ_UNSIGNED #(.width(4)) u_eq_142 (
        .y(_node_126),
        .a(4'd8),
        .b(_value__q)
    );
    wire [15:0] _node_127;
    MUX_UNSIGNED #(.width(16)) u_mux_143 (
        .y(_node_127),
        .sel(_node_126),
        .a(_T_162_8),
        .b(_node_125)
    );
    wire _node_128;
    EQ_UNSIGNED #(.width(4)) u_eq_144 (
        .y(_node_128),
        .a(4'd9),
        .b(_value__q)
    );
    wire [15:0] _node_129;
    MUX_UNSIGNED #(.width(16)) u_mux_145 (
        .y(_node_129),
        .sel(_node_128),
        .a(_T_162_9),
        .b(_node_127)
    );
    wire _node_130;
    EQ_UNSIGNED #(.width(4)) u_eq_146 (
        .y(_node_130),
        .a(4'd10),
        .b(_value__q)
    );
    wire [15:0] _node_131;
    MUX_UNSIGNED #(.width(16)) u_mux_147 (
        .y(_node_131),
        .sel(_node_130),
        .a(_T_162_10),
        .b(_node_129)
    );
    wire [15:0] _T_190_0;
    wire [15:0] _T_190_1;
    wire [15:0] _T_190_2;
    wire [15:0] _T_190_3;
    wire [15:0] _T_190_4;
    wire [15:0] _T_190_5;
    wire [15:0] _T_190_6;
    wire [15:0] _T_190_7;
    wire [15:0] _T_190_8;
    wire [15:0] _T_190_9;
    wire [15:0] _T_190_10;
    wire _node_132;
    EQ_UNSIGNED #(.width(4)) u_eq_148 (
        .y(_node_132),
        .a(4'd0),
        .b(_value__q)
    );
    wire [15:0] _node_133;
    assign _node_133 = _T_190_0;
    wire _node_134;
    EQ_UNSIGNED #(.width(4)) u_eq_149 (
        .y(_node_134),
        .a(4'd1),
        .b(_value__q)
    );
    wire [15:0] _node_135;
    MUX_UNSIGNED #(.width(16)) u_mux_150 (
        .y(_node_135),
        .sel(_node_134),
        .a(_T_190_1),
        .b(_node_133)
    );
    wire _node_136;
    EQ_UNSIGNED #(.width(4)) u_eq_151 (
        .y(_node_136),
        .a(4'd2),
        .b(_value__q)
    );
    wire [15:0] _node_137;
    MUX_UNSIGNED #(.width(16)) u_mux_152 (
        .y(_node_137),
        .sel(_node_136),
        .a(_T_190_2),
        .b(_node_135)
    );
    wire _node_138;
    EQ_UNSIGNED #(.width(4)) u_eq_153 (
        .y(_node_138),
        .a(4'd3),
        .b(_value__q)
    );
    wire [15:0] _node_139;
    MUX_UNSIGNED #(.width(16)) u_mux_154 (
        .y(_node_139),
        .sel(_node_138),
        .a(_T_190_3),
        .b(_node_137)
    );
    wire _node_140;
    EQ_UNSIGNED #(.width(4)) u_eq_155 (
        .y(_node_140),
        .a(4'd4),
        .b(_value__q)
    );
    wire [15:0] _node_141;
    MUX_UNSIGNED #(.width(16)) u_mux_156 (
        .y(_node_141),
        .sel(_node_140),
        .a(_T_190_4),
        .b(_node_139)
    );
    wire _node_142;
    EQ_UNSIGNED #(.width(4)) u_eq_157 (
        .y(_node_142),
        .a(4'd5),
        .b(_value__q)
    );
    wire [15:0] _node_143;
    MUX_UNSIGNED #(.width(16)) u_mux_158 (
        .y(_node_143),
        .sel(_node_142),
        .a(_T_190_5),
        .b(_node_141)
    );
    wire _node_144;
    EQ_UNSIGNED #(.width(4)) u_eq_159 (
        .y(_node_144),
        .a(4'd6),
        .b(_value__q)
    );
    wire [15:0] _node_145;
    MUX_UNSIGNED #(.width(16)) u_mux_160 (
        .y(_node_145),
        .sel(_node_144),
        .a(_T_190_6),
        .b(_node_143)
    );
    wire _node_146;
    EQ_UNSIGNED #(.width(4)) u_eq_161 (
        .y(_node_146),
        .a(4'd7),
        .b(_value__q)
    );
    wire [15:0] _node_147;
    MUX_UNSIGNED #(.width(16)) u_mux_162 (
        .y(_node_147),
        .sel(_node_146),
        .a(_T_190_7),
        .b(_node_145)
    );
    wire _node_148;
    EQ_UNSIGNED #(.width(4)) u_eq_163 (
        .y(_node_148),
        .a(4'd8),
        .b(_value__q)
    );
    wire [15:0] _node_149;
    MUX_UNSIGNED #(.width(16)) u_mux_164 (
        .y(_node_149),
        .sel(_node_148),
        .a(_T_190_8),
        .b(_node_147)
    );
    wire _node_150;
    EQ_UNSIGNED #(.width(4)) u_eq_165 (
        .y(_node_150),
        .a(4'd9),
        .b(_value__q)
    );
    wire [15:0] _node_151;
    MUX_UNSIGNED #(.width(16)) u_mux_166 (
        .y(_node_151),
        .sel(_node_150),
        .a(_T_190_9),
        .b(_node_149)
    );
    wire _node_152;
    EQ_UNSIGNED #(.width(4)) u_eq_167 (
        .y(_node_152),
        .a(4'd10),
        .b(_value__q)
    );
    wire [15:0] _node_153;
    MUX_UNSIGNED #(.width(16)) u_mux_168 (
        .y(_node_153),
        .sel(_node_152),
        .a(_T_190_10),
        .b(_node_151)
    );
    wire [15:0] _T_218_0;
    wire [15:0] _T_218_1;
    wire [15:0] _T_218_2;
    wire [15:0] _T_218_3;
    wire [15:0] _T_218_4;
    wire [15:0] _T_218_5;
    wire [15:0] _T_218_6;
    wire [15:0] _T_218_7;
    wire [15:0] _T_218_8;
    wire [15:0] _T_218_9;
    wire [15:0] _T_218_10;
    wire _node_154;
    EQ_UNSIGNED #(.width(4)) u_eq_169 (
        .y(_node_154),
        .a(4'd0),
        .b(_value__q)
    );
    wire [15:0] _node_155;
    assign _node_155 = _T_218_0;
    wire _node_156;
    EQ_UNSIGNED #(.width(4)) u_eq_170 (
        .y(_node_156),
        .a(4'd1),
        .b(_value__q)
    );
    wire [15:0] _node_157;
    MUX_UNSIGNED #(.width(16)) u_mux_171 (
        .y(_node_157),
        .sel(_node_156),
        .a(_T_218_1),
        .b(_node_155)
    );
    wire _node_158;
    EQ_UNSIGNED #(.width(4)) u_eq_172 (
        .y(_node_158),
        .a(4'd2),
        .b(_value__q)
    );
    wire [15:0] _node_159;
    MUX_UNSIGNED #(.width(16)) u_mux_173 (
        .y(_node_159),
        .sel(_node_158),
        .a(_T_218_2),
        .b(_node_157)
    );
    wire _node_160;
    EQ_UNSIGNED #(.width(4)) u_eq_174 (
        .y(_node_160),
        .a(4'd3),
        .b(_value__q)
    );
    wire [15:0] _node_161;
    MUX_UNSIGNED #(.width(16)) u_mux_175 (
        .y(_node_161),
        .sel(_node_160),
        .a(_T_218_3),
        .b(_node_159)
    );
    wire _node_162;
    EQ_UNSIGNED #(.width(4)) u_eq_176 (
        .y(_node_162),
        .a(4'd4),
        .b(_value__q)
    );
    wire [15:0] _node_163;
    MUX_UNSIGNED #(.width(16)) u_mux_177 (
        .y(_node_163),
        .sel(_node_162),
        .a(_T_218_4),
        .b(_node_161)
    );
    wire _node_164;
    EQ_UNSIGNED #(.width(4)) u_eq_178 (
        .y(_node_164),
        .a(4'd5),
        .b(_value__q)
    );
    wire [15:0] _node_165;
    MUX_UNSIGNED #(.width(16)) u_mux_179 (
        .y(_node_165),
        .sel(_node_164),
        .a(_T_218_5),
        .b(_node_163)
    );
    wire _node_166;
    EQ_UNSIGNED #(.width(4)) u_eq_180 (
        .y(_node_166),
        .a(4'd6),
        .b(_value__q)
    );
    wire [15:0] _node_167;
    MUX_UNSIGNED #(.width(16)) u_mux_181 (
        .y(_node_167),
        .sel(_node_166),
        .a(_T_218_6),
        .b(_node_165)
    );
    wire _node_168;
    EQ_UNSIGNED #(.width(4)) u_eq_182 (
        .y(_node_168),
        .a(4'd7),
        .b(_value__q)
    );
    wire [15:0] _node_169;
    MUX_UNSIGNED #(.width(16)) u_mux_183 (
        .y(_node_169),
        .sel(_node_168),
        .a(_T_218_7),
        .b(_node_167)
    );
    wire _node_170;
    EQ_UNSIGNED #(.width(4)) u_eq_184 (
        .y(_node_170),
        .a(4'd8),
        .b(_value__q)
    );
    wire [15:0] _node_171;
    MUX_UNSIGNED #(.width(16)) u_mux_185 (
        .y(_node_171),
        .sel(_node_170),
        .a(_T_218_8),
        .b(_node_169)
    );
    wire _node_172;
    EQ_UNSIGNED #(.width(4)) u_eq_186 (
        .y(_node_172),
        .a(4'd9),
        .b(_value__q)
    );
    wire [15:0] _node_173;
    MUX_UNSIGNED #(.width(16)) u_mux_187 (
        .y(_node_173),
        .sel(_node_172),
        .a(_T_218_9),
        .b(_node_171)
    );
    wire _node_174;
    EQ_UNSIGNED #(.width(4)) u_eq_188 (
        .y(_node_174),
        .a(4'd10),
        .b(_value__q)
    );
    wire [15:0] _node_175;
    MUX_UNSIGNED #(.width(16)) u_mux_189 (
        .y(_node_175),
        .sel(_node_174),
        .a(_T_218_10),
        .b(_node_173)
    );
    wire [15:0] _T_246_0;
    wire [15:0] _T_246_1;
    wire [15:0] _T_246_2;
    wire [15:0] _T_246_3;
    wire [15:0] _T_246_4;
    wire [15:0] _T_246_5;
    wire [15:0] _T_246_6;
    wire [15:0] _T_246_7;
    wire [15:0] _T_246_8;
    wire [15:0] _T_246_9;
    wire [15:0] _T_246_10;
    wire _node_176;
    EQ_UNSIGNED #(.width(4)) u_eq_190 (
        .y(_node_176),
        .a(4'd0),
        .b(_value__q)
    );
    wire [15:0] _node_177;
    assign _node_177 = _T_246_0;
    wire _node_178;
    EQ_UNSIGNED #(.width(4)) u_eq_191 (
        .y(_node_178),
        .a(4'd1),
        .b(_value__q)
    );
    wire [15:0] _node_179;
    MUX_UNSIGNED #(.width(16)) u_mux_192 (
        .y(_node_179),
        .sel(_node_178),
        .a(_T_246_1),
        .b(_node_177)
    );
    wire _node_180;
    EQ_UNSIGNED #(.width(4)) u_eq_193 (
        .y(_node_180),
        .a(4'd2),
        .b(_value__q)
    );
    wire [15:0] _node_181;
    MUX_UNSIGNED #(.width(16)) u_mux_194 (
        .y(_node_181),
        .sel(_node_180),
        .a(_T_246_2),
        .b(_node_179)
    );
    wire _node_182;
    EQ_UNSIGNED #(.width(4)) u_eq_195 (
        .y(_node_182),
        .a(4'd3),
        .b(_value__q)
    );
    wire [15:0] _node_183;
    MUX_UNSIGNED #(.width(16)) u_mux_196 (
        .y(_node_183),
        .sel(_node_182),
        .a(_T_246_3),
        .b(_node_181)
    );
    wire _node_184;
    EQ_UNSIGNED #(.width(4)) u_eq_197 (
        .y(_node_184),
        .a(4'd4),
        .b(_value__q)
    );
    wire [15:0] _node_185;
    MUX_UNSIGNED #(.width(16)) u_mux_198 (
        .y(_node_185),
        .sel(_node_184),
        .a(_T_246_4),
        .b(_node_183)
    );
    wire _node_186;
    EQ_UNSIGNED #(.width(4)) u_eq_199 (
        .y(_node_186),
        .a(4'd5),
        .b(_value__q)
    );
    wire [15:0] _node_187;
    MUX_UNSIGNED #(.width(16)) u_mux_200 (
        .y(_node_187),
        .sel(_node_186),
        .a(_T_246_5),
        .b(_node_185)
    );
    wire _node_188;
    EQ_UNSIGNED #(.width(4)) u_eq_201 (
        .y(_node_188),
        .a(4'd6),
        .b(_value__q)
    );
    wire [15:0] _node_189;
    MUX_UNSIGNED #(.width(16)) u_mux_202 (
        .y(_node_189),
        .sel(_node_188),
        .a(_T_246_6),
        .b(_node_187)
    );
    wire _node_190;
    EQ_UNSIGNED #(.width(4)) u_eq_203 (
        .y(_node_190),
        .a(4'd7),
        .b(_value__q)
    );
    wire [15:0] _node_191;
    MUX_UNSIGNED #(.width(16)) u_mux_204 (
        .y(_node_191),
        .sel(_node_190),
        .a(_T_246_7),
        .b(_node_189)
    );
    wire _node_192;
    EQ_UNSIGNED #(.width(4)) u_eq_205 (
        .y(_node_192),
        .a(4'd8),
        .b(_value__q)
    );
    wire [15:0] _node_193;
    MUX_UNSIGNED #(.width(16)) u_mux_206 (
        .y(_node_193),
        .sel(_node_192),
        .a(_T_246_8),
        .b(_node_191)
    );
    wire _node_194;
    EQ_UNSIGNED #(.width(4)) u_eq_207 (
        .y(_node_194),
        .a(4'd9),
        .b(_value__q)
    );
    wire [15:0] _node_195;
    MUX_UNSIGNED #(.width(16)) u_mux_208 (
        .y(_node_195),
        .sel(_node_194),
        .a(_T_246_9),
        .b(_node_193)
    );
    wire _node_196;
    EQ_UNSIGNED #(.width(4)) u_eq_209 (
        .y(_node_196),
        .a(4'd10),
        .b(_value__q)
    );
    wire [15:0] _node_197;
    MUX_UNSIGNED #(.width(16)) u_mux_210 (
        .y(_node_197),
        .sel(_node_196),
        .a(_T_246_10),
        .b(_node_195)
    );
    wire [15:0] _T_274_0;
    wire [15:0] _T_274_1;
    wire [15:0] _T_274_2;
    wire [15:0] _T_274_3;
    wire [15:0] _T_274_4;
    wire [15:0] _T_274_5;
    wire [15:0] _T_274_6;
    wire [15:0] _T_274_7;
    wire [15:0] _T_274_8;
    wire [15:0] _T_274_9;
    wire [15:0] _T_274_10;
    wire _node_198;
    EQ_UNSIGNED #(.width(4)) u_eq_211 (
        .y(_node_198),
        .a(4'd0),
        .b(_value__q)
    );
    wire [15:0] _node_199;
    assign _node_199 = _T_274_0;
    wire _node_200;
    EQ_UNSIGNED #(.width(4)) u_eq_212 (
        .y(_node_200),
        .a(4'd1),
        .b(_value__q)
    );
    wire [15:0] _node_201;
    MUX_UNSIGNED #(.width(16)) u_mux_213 (
        .y(_node_201),
        .sel(_node_200),
        .a(_T_274_1),
        .b(_node_199)
    );
    wire _node_202;
    EQ_UNSIGNED #(.width(4)) u_eq_214 (
        .y(_node_202),
        .a(4'd2),
        .b(_value__q)
    );
    wire [15:0] _node_203;
    MUX_UNSIGNED #(.width(16)) u_mux_215 (
        .y(_node_203),
        .sel(_node_202),
        .a(_T_274_2),
        .b(_node_201)
    );
    wire _node_204;
    EQ_UNSIGNED #(.width(4)) u_eq_216 (
        .y(_node_204),
        .a(4'd3),
        .b(_value__q)
    );
    wire [15:0] _node_205;
    MUX_UNSIGNED #(.width(16)) u_mux_217 (
        .y(_node_205),
        .sel(_node_204),
        .a(_T_274_3),
        .b(_node_203)
    );
    wire _node_206;
    EQ_UNSIGNED #(.width(4)) u_eq_218 (
        .y(_node_206),
        .a(4'd4),
        .b(_value__q)
    );
    wire [15:0] _node_207;
    MUX_UNSIGNED #(.width(16)) u_mux_219 (
        .y(_node_207),
        .sel(_node_206),
        .a(_T_274_4),
        .b(_node_205)
    );
    wire _node_208;
    EQ_UNSIGNED #(.width(4)) u_eq_220 (
        .y(_node_208),
        .a(4'd5),
        .b(_value__q)
    );
    wire [15:0] _node_209;
    MUX_UNSIGNED #(.width(16)) u_mux_221 (
        .y(_node_209),
        .sel(_node_208),
        .a(_T_274_5),
        .b(_node_207)
    );
    wire _node_210;
    EQ_UNSIGNED #(.width(4)) u_eq_222 (
        .y(_node_210),
        .a(4'd6),
        .b(_value__q)
    );
    wire [15:0] _node_211;
    MUX_UNSIGNED #(.width(16)) u_mux_223 (
        .y(_node_211),
        .sel(_node_210),
        .a(_T_274_6),
        .b(_node_209)
    );
    wire _node_212;
    EQ_UNSIGNED #(.width(4)) u_eq_224 (
        .y(_node_212),
        .a(4'd7),
        .b(_value__q)
    );
    wire [15:0] _node_213;
    MUX_UNSIGNED #(.width(16)) u_mux_225 (
        .y(_node_213),
        .sel(_node_212),
        .a(_T_274_7),
        .b(_node_211)
    );
    wire _node_214;
    EQ_UNSIGNED #(.width(4)) u_eq_226 (
        .y(_node_214),
        .a(4'd8),
        .b(_value__q)
    );
    wire [15:0] _node_215;
    MUX_UNSIGNED #(.width(16)) u_mux_227 (
        .y(_node_215),
        .sel(_node_214),
        .a(_T_274_8),
        .b(_node_213)
    );
    wire _node_216;
    EQ_UNSIGNED #(.width(4)) u_eq_228 (
        .y(_node_216),
        .a(4'd9),
        .b(_value__q)
    );
    wire [15:0] _node_217;
    MUX_UNSIGNED #(.width(16)) u_mux_229 (
        .y(_node_217),
        .sel(_node_216),
        .a(_T_274_9),
        .b(_node_215)
    );
    wire _node_218;
    EQ_UNSIGNED #(.width(4)) u_eq_230 (
        .y(_node_218),
        .a(4'd10),
        .b(_value__q)
    );
    wire [15:0] _node_219;
    MUX_UNSIGNED #(.width(16)) u_mux_231 (
        .y(_node_219),
        .sel(_node_218),
        .a(_T_274_10),
        .b(_node_217)
    );
    wire [15:0] _T_292;
    wire [15:0] _T_296;
    wire [15:0] _T_300;
    wire [15:0] _T_304;
    wire [15:0] _T_308;
    wire [15:0] _T_312;
    wire [15:0] _T_316;
    wire [15:0] _T_320;
    wire [15:0] _T_324;
    wire [15:0] _T_328;
    wire [15:0] _T_332;
    wire [15:0] _T_335_0;
    wire [15:0] _T_335_1;
    wire [15:0] _T_335_2;
    wire [15:0] _T_335_3;
    wire [15:0] _T_335_4;
    wire [15:0] _T_335_5;
    wire [15:0] _T_335_6;
    wire [15:0] _T_335_7;
    wire [15:0] _T_335_8;
    wire [15:0] _T_335_9;
    wire [15:0] _T_335_10;
    wire _T_362_0;
    wire _T_362_1;
    wire _T_362_2;
    wire _T_362_3;
    wire _T_362_4;
    wire _T_362_5;
    wire _T_362_6;
    wire _T_362_7;
    wire _T_362_8;
    wire _T_362_9;
    wire _T_362_10;
    wire _node_220;
    EQ_UNSIGNED #(.width(4)) u_eq_232 (
        .y(_node_220),
        .a(4'd0),
        .b(_value__q)
    );
    wire [15:0] _node_221;
    assign _node_221 = _T_335_0;
    wire _node_222;
    EQ_UNSIGNED #(.width(4)) u_eq_233 (
        .y(_node_222),
        .a(4'd1),
        .b(_value__q)
    );
    wire [15:0] _node_223;
    MUX_UNSIGNED #(.width(16)) u_mux_234 (
        .y(_node_223),
        .sel(_node_222),
        .a(_T_335_1),
        .b(_node_221)
    );
    wire _node_224;
    EQ_UNSIGNED #(.width(4)) u_eq_235 (
        .y(_node_224),
        .a(4'd2),
        .b(_value__q)
    );
    wire [15:0] _node_225;
    MUX_UNSIGNED #(.width(16)) u_mux_236 (
        .y(_node_225),
        .sel(_node_224),
        .a(_T_335_2),
        .b(_node_223)
    );
    wire _node_226;
    EQ_UNSIGNED #(.width(4)) u_eq_237 (
        .y(_node_226),
        .a(4'd3),
        .b(_value__q)
    );
    wire [15:0] _node_227;
    MUX_UNSIGNED #(.width(16)) u_mux_238 (
        .y(_node_227),
        .sel(_node_226),
        .a(_T_335_3),
        .b(_node_225)
    );
    wire _node_228;
    EQ_UNSIGNED #(.width(4)) u_eq_239 (
        .y(_node_228),
        .a(4'd4),
        .b(_value__q)
    );
    wire [15:0] _node_229;
    MUX_UNSIGNED #(.width(16)) u_mux_240 (
        .y(_node_229),
        .sel(_node_228),
        .a(_T_335_4),
        .b(_node_227)
    );
    wire _node_230;
    EQ_UNSIGNED #(.width(4)) u_eq_241 (
        .y(_node_230),
        .a(4'd5),
        .b(_value__q)
    );
    wire [15:0] _node_231;
    MUX_UNSIGNED #(.width(16)) u_mux_242 (
        .y(_node_231),
        .sel(_node_230),
        .a(_T_335_5),
        .b(_node_229)
    );
    wire _node_232;
    EQ_UNSIGNED #(.width(4)) u_eq_243 (
        .y(_node_232),
        .a(4'd6),
        .b(_value__q)
    );
    wire [15:0] _node_233;
    MUX_UNSIGNED #(.width(16)) u_mux_244 (
        .y(_node_233),
        .sel(_node_232),
        .a(_T_335_6),
        .b(_node_231)
    );
    wire _node_234;
    EQ_UNSIGNED #(.width(4)) u_eq_245 (
        .y(_node_234),
        .a(4'd7),
        .b(_value__q)
    );
    wire [15:0] _node_235;
    MUX_UNSIGNED #(.width(16)) u_mux_246 (
        .y(_node_235),
        .sel(_node_234),
        .a(_T_335_7),
        .b(_node_233)
    );
    wire _node_236;
    EQ_UNSIGNED #(.width(4)) u_eq_247 (
        .y(_node_236),
        .a(4'd8),
        .b(_value__q)
    );
    wire [15:0] _node_237;
    MUX_UNSIGNED #(.width(16)) u_mux_248 (
        .y(_node_237),
        .sel(_node_236),
        .a(_T_335_8),
        .b(_node_235)
    );
    wire _node_238;
    EQ_UNSIGNED #(.width(4)) u_eq_249 (
        .y(_node_238),
        .a(4'd9),
        .b(_value__q)
    );
    wire [15:0] _node_239;
    MUX_UNSIGNED #(.width(16)) u_mux_250 (
        .y(_node_239),
        .sel(_node_238),
        .a(_T_335_9),
        .b(_node_237)
    );
    wire _node_240;
    EQ_UNSIGNED #(.width(4)) u_eq_251 (
        .y(_node_240),
        .a(4'd10),
        .b(_value__q)
    );
    wire [15:0] _node_241;
    MUX_UNSIGNED #(.width(16)) u_mux_252 (
        .y(_node_241),
        .sel(_node_240),
        .a(_T_335_10),
        .b(_node_239)
    );
    wire _T_378;
    EQ_UNSIGNED #(.width(16)) u_eq_253 (
        .y(_T_378),
        .a(_c__io_out),
        .b(_node_241)
    );
    wire _T_380;
    EQ_UNSIGNED #(.width(1)) u_eq_254 (
        .y(_T_380),
        .a(_T_378),
        .b(1'h0)
    );
    wire _T_383;
    EQ_UNSIGNED #(.width(1)) u_eq_255 (
        .y(_T_383),
        .a(reset),
        .b(1'h0)
    );
    wire _T_385;
    BITWISEOR #(.width(1)) bitwiseor_256 (
        .y(_T_385),
        .a(1'h0),
        .b(reset)
    );
    wire _T_387;
    EQ_UNSIGNED #(.width(1)) u_eq_257 (
        .y(_T_387),
        .a(_T_385),
        .b(1'h0)
    );
    wire _T_389;
    EQ_UNSIGNED #(.width(1)) u_eq_258 (
        .y(_T_389),
        .a(reset),
        .b(1'h0)
    );
    wire _T_391;
    EQ_UNSIGNED #(.width(4)) u_eq_259 (
        .y(_T_391),
        .a(_value__q),
        .b(4'hA)
    );
    wire [4:0] _T_393;
    wire [3:0] _WTEMP_2;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_260 (
        .y(_WTEMP_2),
        .in(1'h1)
    );
    ADD_UNSIGNED #(.width(4)) u_add_261 (
        .y(_T_393),
        .a(_value__q),
        .b(_WTEMP_2)
    );
    wire [3:0] _T_394;
    TAIL #(.width(5), .n(1)) tail_262 (
        .y(_T_394),
        .in(_T_393)
    );
    wire _T_397;
    EQ_UNSIGNED #(.width(1)) u_eq_263 (
        .y(_T_397),
        .a(reset),
        .b(1'h0)
    );
    wire _T_400;
    EQ_UNSIGNED #(.width(1)) u_eq_264 (
        .y(_T_400),
        .a(reset),
        .b(1'h0)
    );
    wire _node_242;
    MUX_UNSIGNED #(.width(1)) u_mux_265 (
        .y(_node_242),
        .sel(_T_391),
        .a(1'h1),
        .b(__T_6__q)
    );
    wire [3:0] _node_243;
    wire [3:0] _WTEMP_3;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_266 (
        .y(_WTEMP_3),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(4)) u_mux_267 (
        .y(_node_243),
        .sel(_T_391),
        .a(_WTEMP_3),
        .b(_T_394)
    );
    assign _T_106_0 = 16'h2249;
    assign _T_106_1 = 16'h24AA;
    assign _T_106_10 = 16'h773;
    assign _T_106_2 = 16'h56B9;
    assign _T_106_3 = 16'h2DD2;
    assign _T_106_4 = 16'hC574;
    assign _T_106_5 = 16'h3A4;
    assign _T_106_6 = 16'hE213;
    assign _T_106_7 = 16'hCDEC;
    assign _T_106_8 = 16'hFDEF;
    assign _T_106_9 = 16'h773;
    assign _T_134_0 = 16'hB9CC;
    assign _T_134_1 = 16'hABCB;
    assign _T_134_10 = 16'hC9A8;
    assign _T_134_2 = 16'hB083;
    assign _T_134_3 = 16'h88AA;
    assign _T_134_4 = 16'h6A2E;
    assign _T_134_5 = 16'h652C;
    assign _T_134_6 = 16'hEE10;
    assign _T_134_7 = 16'hE781;
    assign _T_134_8 = 16'h78B3;
    assign _T_134_9 = 16'hC9A8;
    assign _T_162_0 = 16'hFA83;
    assign _T_162_1 = 16'h125;
    assign _T_162_10 = 16'hF8D1;
    assign _T_162_2 = 16'hF8B7;
    assign _T_162_3 = 16'hDABF;
    assign _T_162_4 = 16'h3613;
    assign _T_162_5 = 16'hDA92;
    assign _T_162_6 = 16'hF64A;
    assign _T_162_7 = 16'h764B;
    assign _T_162_8 = 16'h5A65;
    assign _T_162_9 = 16'hF8D1;
    assign _T_190_0 = 16'h8BCF;
    assign _T_190_1 = 16'h5BF2;
    assign _T_190_10 = 16'h1CD4;
    assign _T_190_2 = 16'h9B40;
    assign _T_190_3 = 16'h4FB6;
    assign _T_190_4 = 16'hF2BC;
    assign _T_190_5 = 16'h9E56;
    assign _T_190_6 = 16'h7A93;
    assign _T_190_7 = 16'hA820;
    assign _T_190_8 = 16'h916F;
    assign _T_190_9 = 16'h1CD4;
    assign _T_218_0 = 16'hE63A;
    assign _T_218_1 = 16'hB70C;
    assign _T_218_10 = 16'h1255;
    assign _T_218_2 = 16'h5932;
    assign _T_218_3 = 16'h9CD2;
    assign _T_218_4 = 16'hB13A;
    assign _T_218_5 = 16'hF201;
    assign _T_218_6 = 16'hFE54;
    assign _T_218_7 = 16'hAD67;
    assign _T_218_8 = 16'h8078;
    assign _T_218_9 = 16'h1255;
    assign _T_22_0 = 16'h6987;
    assign _T_22_1 = 16'h4E8F;
    assign _T_22_10 = 16'h601D;
    assign _T_22_2 = 16'hAAB6;
    assign _T_22_3 = 16'hBE94;
    assign _T_22_4 = 16'h1531;
    assign _T_22_5 = 16'hC54;
    assign _T_22_6 = 16'h64C;
    assign _T_22_7 = 16'h30CC;
    assign _T_22_8 = 16'h189C;
    assign _T_22_9 = 16'h601D;
    assign _T_246_0 = 16'h1543;
    assign _T_246_1 = 16'h7684;
    assign _T_246_10 = 16'h7BD1;
    assign _T_246_2 = 16'hDBFE;
    assign _T_246_3 = 16'h37B2;
    assign _T_246_4 = 16'hB672;
    assign _T_246_5 = 16'h64EA;
    assign _T_246_6 = 16'h2B98;
    assign _T_246_7 = 16'h7101;
    assign _T_246_8 = 16'hF822;
    assign _T_246_9 = 16'h7BD1;
    assign _T_274_0 = 16'h2F9D;
    assign _T_274_1 = 16'h4635;
    assign _T_274_10 = 16'h234;
    assign _T_274_2 = 16'hEEAF;
    assign _T_274_3 = 16'h3412;
    assign _T_274_4 = 16'hB09F;
    assign _T_274_5 = 16'h9C95;
    assign _T_274_6 = 16'h24CC;
    assign _T_274_7 = 16'h5210;
    assign _T_274_8 = 16'h90C3;
    assign _T_274_9 = 16'h234;
    assign _T_292 = 16'hFC13;
    assign _T_296 = 16'hB8EC;
    assign _T_300 = 16'hF8B7;
    assign _T_304 = 16'hDDA1;
    assign _T_308 = 16'hF2BC;
    assign _T_312 = 16'hF201;
    assign _T_316 = 16'hFE54;
    assign _T_320 = 16'hE781;
    assign _T_324 = 16'hFDEF;
    assign _T_328 = 16'hF8D1;
    PAD_UNSIGNED #(.width(1), .n(16)) u_pad_268 (
        .y(_T_332),
        .in(1'h0)
    );
    assign _T_335_0 = _T_292;
    assign _T_335_1 = _T_296;
    assign _T_335_10 = _T_332;
    assign _T_335_2 = _T_300;
    assign _T_335_3 = _T_304;
    assign _T_335_4 = _T_308;
    assign _T_335_5 = _T_312;
    assign _T_335_6 = _T_316;
    assign _T_335_7 = _T_320;
    assign _T_335_8 = _T_324;
    assign _T_335_9 = _T_328;
    assign _T_362_0 = 1'h1;
    assign _T_362_1 = 1'h1;
    assign _T_362_10 = 1'h0;
    assign _T_362_2 = 1'h1;
    assign _T_362_3 = 1'h1;
    assign _T_362_4 = 1'h1;
    assign _T_362_5 = 1'h1;
    assign _T_362_6 = 1'h1;
    assign _T_362_7 = 1'h1;
    assign _T_362_8 = 1'h1;
    assign _T_362_9 = 1'h1;
    assign _T_50_0 = 16'hFC13;
    assign _T_50_1 = 16'h1074;
    assign _T_50_10 = 16'hCD;
    assign _T_50_2 = 16'hD0E1;
    assign _T_50_3 = 16'hB81;
    assign _T_50_4 = 16'h4073;
    assign _T_50_5 = 16'hC49D;
    assign _T_50_6 = 16'h50F8;
    assign _T_50_7 = 16'h4982;
    assign _T_50_8 = 16'hB681;
    assign _T_50_9 = 16'hCD;
    MUX_UNSIGNED #(.width(1)) u_mux_269 (
        .y(_WTEMP_1),
        .sel(_T_8),
        .a(_node_242),
        .b(__T_6__q)
    );
    assign _T_78_0 = 16'h86D5;
    assign _T_78_1 = 16'hB8EC;
    assign _T_78_10 = 16'hC19;
    assign _T_78_2 = 16'h124D;
    assign _T_78_3 = 16'hDDA1;
    assign _T_78_4 = 16'h279;
    assign _T_78_5 = 16'hC878;
    assign _T_78_6 = 16'hC93A;
    assign _T_78_7 = 16'hB96B;
    assign _T_78_8 = 16'hDA52;
    assign _T_78_9 = 16'hC19;
    assign _c__clock = clock;
    assign _c__io_ins_0 = _node_21;
    assign _c__io_ins_1 = _node_65;
    assign _c__io_ins_2 = _node_109;
    assign _c__io_ins_3 = _node_175;
    assign _c__io_ins_4 = _node_43;
    assign _c__io_ins_5 = _node_87;
    assign _c__io_ins_6 = _node_153;
    assign _c__io_ins_7 = _node_197;
    assign _c__io_ins_8 = _node_219;
    assign _c__io_ins_9 = _node_131;
    assign _c__reset = reset;
    MUX_UNSIGNED #(.width(4)) u_mux_270 (
        .y(_WTEMP_0),
        .sel(_T_8),
        .a(_node_243),
        .b(_value__q)
    );
endmodule //MaxNTests
module MaxN(
    input clock,
    input reset,
    input [15:0] io_ins_0,
    input [15:0] io_ins_1,
    input [15:0] io_ins_2,
    input [15:0] io_ins_3,
    input [15:0] io_ins_4,
    input [15:0] io_ins_5,
    input [15:0] io_ins_6,
    input [15:0] io_ins_7,
    input [15:0] io_ins_8,
    input [15:0] io_ins_9,
    output [15:0] io_out
);
    wire _T_6;
    GT_UNSIGNED #(.width(16)) u_gt_1 (
        .y(_T_6),
        .a(io_ins_0),
        .b(io_ins_1)
    );
    wire [15:0] _T_7;
    MUX_UNSIGNED #(.width(16)) u_mux_2 (
        .y(_T_7),
        .sel(_T_6),
        .a(io_ins_0),
        .b(io_ins_1)
    );
    wire _T_8;
    GT_UNSIGNED #(.width(16)) u_gt_3 (
        .y(_T_8),
        .a(_T_7),
        .b(io_ins_2)
    );
    wire [15:0] _T_9;
    MUX_UNSIGNED #(.width(16)) u_mux_4 (
        .y(_T_9),
        .sel(_T_8),
        .a(_T_7),
        .b(io_ins_2)
    );
    wire _T_10;
    GT_UNSIGNED #(.width(16)) u_gt_5 (
        .y(_T_10),
        .a(_T_9),
        .b(io_ins_3)
    );
    wire [15:0] _T_11;
    MUX_UNSIGNED #(.width(16)) u_mux_6 (
        .y(_T_11),
        .sel(_T_10),
        .a(_T_9),
        .b(io_ins_3)
    );
    wire _T_12;
    GT_UNSIGNED #(.width(16)) u_gt_7 (
        .y(_T_12),
        .a(_T_11),
        .b(io_ins_4)
    );
    wire [15:0] _T_13;
    MUX_UNSIGNED #(.width(16)) u_mux_8 (
        .y(_T_13),
        .sel(_T_12),
        .a(_T_11),
        .b(io_ins_4)
    );
    wire _T_14;
    GT_UNSIGNED #(.width(16)) u_gt_9 (
        .y(_T_14),
        .a(_T_13),
        .b(io_ins_5)
    );
    wire [15:0] _T_15;
    MUX_UNSIGNED #(.width(16)) u_mux_10 (
        .y(_T_15),
        .sel(_T_14),
        .a(_T_13),
        .b(io_ins_5)
    );
    wire _T_16;
    GT_UNSIGNED #(.width(16)) u_gt_11 (
        .y(_T_16),
        .a(_T_15),
        .b(io_ins_6)
    );
    wire [15:0] _T_17;
    MUX_UNSIGNED #(.width(16)) u_mux_12 (
        .y(_T_17),
        .sel(_T_16),
        .a(_T_15),
        .b(io_ins_6)
    );
    wire _T_18;
    GT_UNSIGNED #(.width(16)) u_gt_13 (
        .y(_T_18),
        .a(_T_17),
        .b(io_ins_7)
    );
    wire [15:0] _T_19;
    MUX_UNSIGNED #(.width(16)) u_mux_14 (
        .y(_T_19),
        .sel(_T_18),
        .a(_T_17),
        .b(io_ins_7)
    );
    wire _T_20;
    GT_UNSIGNED #(.width(16)) u_gt_15 (
        .y(_T_20),
        .a(_T_19),
        .b(io_ins_8)
    );
    wire [15:0] _T_21;
    MUX_UNSIGNED #(.width(16)) u_mux_16 (
        .y(_T_21),
        .sel(_T_20),
        .a(_T_19),
        .b(io_ins_8)
    );
    wire _T_22;
    GT_UNSIGNED #(.width(16)) u_gt_17 (
        .y(_T_22),
        .a(_T_21),
        .b(io_ins_9)
    );
    wire [15:0] _T_23;
    MUX_UNSIGNED #(.width(16)) u_mux_18 (
        .y(_T_23),
        .sel(_T_22),
        .a(_T_21),
        .b(io_ins_9)
    );
    assign io_out = _T_23;
endmodule //MaxN
module GT_UNSIGNED(y, a, b);
    parameter width = 4;
    output y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a > b;
endmodule // GT_UNSIGNED
module MUX_UNSIGNED(y, sel, a, b);
    parameter width = 4;
    output [width-1:0] y;
    input sel;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = sel ? a : b;
endmodule // MUX_UNSIGNED
module DFF_POSCLK(q, d, clk);
    parameter width = 4;
    output reg [width-1:0] q;
    input [width-1:0] d;
    input clk;
    always @(posedge clk) begin
        q <= d;
    end
endmodule // DFF_POSCLK
module EQ_UNSIGNED(y, a, b);
    parameter width = 4;
    output y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a == b;
endmodule // EQ_UNSIGNED
module BITWISEOR(y, a, b);
    parameter width = 4;
    output [width-1:0] y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a | b;
endmodule // BITWISEOR
module PAD_UNSIGNED(y, in);
    parameter width = 4;
    parameter n = 4;
    output [(n > width ? n : width)-1:0] y;
    input [width-1:0] in;
    assign y = (n > width) ? {{(n - width){1'b0}}, in} : in;
endmodule // PAD_UNSIGNED
module ADD_UNSIGNED(y, a, b);
    parameter width = 4;
    output [width:0] y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a + b;
endmodule // ADD_UNSIGNED
module TAIL(y, in);
    parameter width = 4;
    parameter n = 2;
    output [width-n-1:0] y;
    input [width-1:0] in;
    assign y = in[width-n-1:0];
endmodule // TAIL
