module DutWithLogging(
  input   clock,
  input   reset
);
endmodule
