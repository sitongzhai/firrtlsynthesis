module IntervalChainedSubTester(
    input clock,
    input reset
);
    wire [4:0] intervalResult1;
    wire [4:0] intervalResult2;
    wire [10:0] uIntResult;
    wire [11:0] sIntResult;
    wire [11:0] fixedResult;
    wire [5:0] _node_0;
    ASSINT #(.width(6)) assint_1 (
        .y(_node_0),
        .in(6'h11)
    );
    wire [2:0] _node_1;
    ASSINT #(.width(3)) assint_2 (
        .y(_node_1),
        .in(3'h2)
    );
    wire [6:0] _intervalResult1_T;
    wire [5:0] _WTEMP_0;
    PAD_SIGNED #(.width(3), .n(6)) s_pad_3 (
        .y(_WTEMP_0),
        .in(_node_1)
    );
    SUB_SIGNED #(.width(6)) s_sub_4 (
        .y(_intervalResult1_T),
        .a(_node_0),
        .b(_WTEMP_0)
    );
    wire [2:0] _node_2;
    ASSINT #(.width(3)) assint_5 (
        .y(_node_2),
        .in(3'h2)
    );
    wire [7:0] _intervalResult1_T_1;
    wire [6:0] _WTEMP_1;
    PAD_SIGNED #(.width(3), .n(7)) s_pad_6 (
        .y(_WTEMP_1),
        .in(_node_2)
    );
    SUB_SIGNED #(.width(7)) s_sub_7 (
        .y(_intervalResult1_T_1),
        .a(_intervalResult1_T),
        .b(_WTEMP_1)
    );
    wire [2:0] _node_3;
    ASSINT #(.width(3)) assint_8 (
        .y(_node_3),
        .in(3'h2)
    );
    wire [8:0] _intervalResult1_T_2;
    wire [7:0] _WTEMP_2;
    PAD_SIGNED #(.width(3), .n(8)) s_pad_9 (
        .y(_WTEMP_2),
        .in(_node_3)
    );
    SUB_SIGNED #(.width(8)) s_sub_10 (
        .y(_intervalResult1_T_2),
        .a(_intervalResult1_T_1),
        .b(_WTEMP_2)
    );
    wire [2:0] _node_4;
    ASSINT #(.width(3)) assint_11 (
        .y(_node_4),
        .in(3'h2)
    );
    wire [9:0] _intervalResult1_T_3;
    wire [8:0] _WTEMP_3;
    PAD_SIGNED #(.width(3), .n(9)) s_pad_12 (
        .y(_WTEMP_3),
        .in(_node_4)
    );
    SUB_SIGNED #(.width(9)) s_sub_13 (
        .y(_intervalResult1_T_3),
        .a(_intervalResult1_T_2),
        .b(_WTEMP_3)
    );
    wire [2:0] _node_5;
    ASSINT #(.width(3)) assint_14 (
        .y(_node_5),
        .in(3'h2)
    );
    wire [10:0] _intervalResult1_T_4;
    wire [9:0] _WTEMP_4;
    PAD_SIGNED #(.width(3), .n(10)) s_pad_15 (
        .y(_WTEMP_4),
        .in(_node_5)
    );
    SUB_SIGNED #(.width(10)) s_sub_16 (
        .y(_intervalResult1_T_4),
        .a(_intervalResult1_T_3),
        .b(_WTEMP_4)
    );
    wire [2:0] _node_6;
    ASSINT #(.width(3)) assint_17 (
        .y(_node_6),
        .in(3'h2)
    );
    wire [11:0] _intervalResult1_T_5;
    wire [10:0] _WTEMP_5;
    PAD_SIGNED #(.width(3), .n(11)) s_pad_18 (
        .y(_WTEMP_5),
        .in(_node_6)
    );
    SUB_SIGNED #(.width(11)) s_sub_19 (
        .y(_intervalResult1_T_5),
        .a(_intervalResult1_T_4),
        .b(_WTEMP_5)
    );
    wire [5:0] _node_7;
    ASSINT #(.width(6)) assint_20 (
        .y(_node_7),
        .in(6'h11)
    );
    wire [2:0] _node_8;
    ASSINT #(.width(3)) assint_21 (
        .y(_node_8),
        .in(3'h2)
    );
    wire [6:0] _intervalResult2_T;
    wire [5:0] _WTEMP_6;
    PAD_SIGNED #(.width(3), .n(6)) s_pad_22 (
        .y(_WTEMP_6),
        .in(_node_8)
    );
    SUB_SIGNED #(.width(6)) s_sub_23 (
        .y(_intervalResult2_T),
        .a(_node_7),
        .b(_WTEMP_6)
    );
    wire [2:0] _node_9;
    ASSINT #(.width(3)) assint_24 (
        .y(_node_9),
        .in(3'h2)
    );
    wire [7:0] _intervalResult2_T_1;
    wire [6:0] _WTEMP_7;
    PAD_SIGNED #(.width(3), .n(7)) s_pad_25 (
        .y(_WTEMP_7),
        .in(_node_9)
    );
    SUB_SIGNED #(.width(7)) s_sub_26 (
        .y(_intervalResult2_T_1),
        .a(_intervalResult2_T),
        .b(_WTEMP_7)
    );
    wire [2:0] _node_10;
    ASSINT #(.width(3)) assint_27 (
        .y(_node_10),
        .in(3'h2)
    );
    wire [8:0] _intervalResult2_T_2;
    wire [7:0] _WTEMP_8;
    PAD_SIGNED #(.width(3), .n(8)) s_pad_28 (
        .y(_WTEMP_8),
        .in(_node_10)
    );
    SUB_SIGNED #(.width(8)) s_sub_29 (
        .y(_intervalResult2_T_2),
        .a(_intervalResult2_T_1),
        .b(_WTEMP_8)
    );
    wire [2:0] _node_11;
    ASSINT #(.width(3)) assint_30 (
        .y(_node_11),
        .in(3'h2)
    );
    wire [9:0] _intervalResult2_T_3;
    wire [8:0] _WTEMP_9;
    PAD_SIGNED #(.width(3), .n(9)) s_pad_31 (
        .y(_WTEMP_9),
        .in(_node_11)
    );
    SUB_SIGNED #(.width(9)) s_sub_32 (
        .y(_intervalResult2_T_3),
        .a(_intervalResult2_T_2),
        .b(_WTEMP_9)
    );
    wire [2:0] _node_12;
    ASSINT #(.width(3)) assint_33 (
        .y(_node_12),
        .in(3'h2)
    );
    wire [10:0] _intervalResult2_T_4;
    wire [9:0] _WTEMP_10;
    PAD_SIGNED #(.width(3), .n(10)) s_pad_34 (
        .y(_WTEMP_10),
        .in(_node_12)
    );
    SUB_SIGNED #(.width(10)) s_sub_35 (
        .y(_intervalResult2_T_4),
        .a(_intervalResult2_T_3),
        .b(_WTEMP_10)
    );
    wire [2:0] _node_13;
    ASSINT #(.width(3)) assint_36 (
        .y(_node_13),
        .in(3'h2)
    );
    wire [11:0] _intervalResult2_T_5;
    wire [10:0] _WTEMP_11;
    PAD_SIGNED #(.width(3), .n(11)) s_pad_37 (
        .y(_WTEMP_11),
        .in(_node_13)
    );
    SUB_SIGNED #(.width(11)) s_sub_38 (
        .y(_intervalResult2_T_5),
        .a(_intervalResult2_T_4),
        .b(_WTEMP_11)
    );
    wire [5:0] _uIntResult_T;
    assign _uIntResult_T = 6'hF;
    wire [5:0] _uIntResult_T_1;
    assign _uIntResult_T_1 = 6'hF;
    wire [6:0] _uIntResult_T_2;
    assign _uIntResult_T_2 = 7'hD;
    wire [6:0] _uIntResult_T_3;
    assign _uIntResult_T_3 = 7'hD;
    wire [7:0] _uIntResult_T_4;
    assign _uIntResult_T_4 = 8'hB;
    wire [7:0] _uIntResult_T_5;
    assign _uIntResult_T_5 = 8'hB;
    wire [8:0] _uIntResult_T_6;
    assign _uIntResult_T_6 = 9'h9;
    wire [8:0] _uIntResult_T_7;
    assign _uIntResult_T_7 = 9'h9;
    wire [9:0] _uIntResult_T_8;
    assign _uIntResult_T_8 = 10'h7;
    wire [9:0] _uIntResult_T_9;
    assign _uIntResult_T_9 = 10'h7;
    wire [10:0] _uIntResult_T_10;
    assign _uIntResult_T_10 = 11'h5;
    wire [10:0] _uIntResult_T_11;
    assign _uIntResult_T_11 = 11'h5;
    wire [5:0] _node_14;
    ASSINT #(.width(6)) assint_39 (
        .y(_node_14),
        .in(6'h11)
    );
    wire [2:0] _node_15;
    ASSINT #(.width(3)) assint_40 (
        .y(_node_15),
        .in(3'h2)
    );
    wire [6:0] _fixedResult_T;
    wire [5:0] _WTEMP_12;
    PAD_SIGNED #(.width(3), .n(6)) s_pad_41 (
        .y(_WTEMP_12),
        .in(_node_15)
    );
    SUB_SIGNED #(.width(6)) s_sub_42 (
        .y(_fixedResult_T),
        .a(_node_14),
        .b(_WTEMP_12)
    );
    wire [2:0] _node_16;
    ASSINT #(.width(3)) assint_43 (
        .y(_node_16),
        .in(3'h2)
    );
    wire [7:0] _fixedResult_T_1;
    wire [6:0] _WTEMP_13;
    PAD_SIGNED #(.width(3), .n(7)) s_pad_44 (
        .y(_WTEMP_13),
        .in(_node_16)
    );
    SUB_SIGNED #(.width(7)) s_sub_45 (
        .y(_fixedResult_T_1),
        .a(_fixedResult_T),
        .b(_WTEMP_13)
    );
    wire [2:0] _node_17;
    ASSINT #(.width(3)) assint_46 (
        .y(_node_17),
        .in(3'h2)
    );
    wire [8:0] _fixedResult_T_2;
    wire [7:0] _WTEMP_14;
    PAD_SIGNED #(.width(3), .n(8)) s_pad_47 (
        .y(_WTEMP_14),
        .in(_node_17)
    );
    SUB_SIGNED #(.width(8)) s_sub_48 (
        .y(_fixedResult_T_2),
        .a(_fixedResult_T_1),
        .b(_WTEMP_14)
    );
    wire [2:0] _node_18;
    ASSINT #(.width(3)) assint_49 (
        .y(_node_18),
        .in(3'h2)
    );
    wire [9:0] _fixedResult_T_3;
    wire [8:0] _WTEMP_15;
    PAD_SIGNED #(.width(3), .n(9)) s_pad_50 (
        .y(_WTEMP_15),
        .in(_node_18)
    );
    SUB_SIGNED #(.width(9)) s_sub_51 (
        .y(_fixedResult_T_3),
        .a(_fixedResult_T_2),
        .b(_WTEMP_15)
    );
    wire [2:0] _node_19;
    ASSINT #(.width(3)) assint_52 (
        .y(_node_19),
        .in(3'h2)
    );
    wire [10:0] _fixedResult_T_4;
    wire [9:0] _WTEMP_16;
    PAD_SIGNED #(.width(3), .n(10)) s_pad_53 (
        .y(_WTEMP_16),
        .in(_node_19)
    );
    SUB_SIGNED #(.width(10)) s_sub_54 (
        .y(_fixedResult_T_4),
        .a(_fixedResult_T_3),
        .b(_WTEMP_16)
    );
    wire [2:0] _node_20;
    ASSINT #(.width(3)) assint_55 (
        .y(_node_20),
        .in(3'h2)
    );
    wire [11:0] _fixedResult_T_5;
    wire [10:0] _WTEMP_17;
    PAD_SIGNED #(.width(3), .n(11)) s_pad_56 (
        .y(_WTEMP_17),
        .in(_node_20)
    );
    SUB_SIGNED #(.width(11)) s_sub_57 (
        .y(_fixedResult_T_5),
        .a(_fixedResult_T_4),
        .b(_WTEMP_17)
    );
    wire [6:0] _sIntResult_T;
    assign _sIntResult_T = 7'shF;
    wire [7:0] _sIntResult_T_1;
    assign _sIntResult_T_1 = 8'shD;
    wire [8:0] _sIntResult_T_2;
    assign _sIntResult_T_2 = 9'shB;
    wire [9:0] _sIntResult_T_3;
    assign _sIntResult_T_3 = 10'sh9;
    wire [10:0] _sIntResult_T_4;
    assign _sIntResult_T_4 = 11'sh7;
    wire [11:0] _sIntResult_T_5;
    assign _sIntResult_T_5 = 12'sh5;
    wire _T;
    wire [10:0] _WTEMP_18;
    PAD_UNSIGNED #(.width(3), .n(11)) u_pad_58 (
        .y(_WTEMP_18),
        .in(3'h5)
    );
    EQ_UNSIGNED #(.width(11)) u_eq_59 (
        .y(_T),
        .a(uIntResult),
        .b(_WTEMP_18)
    );
    wire _T_1;
    BITS #(.width(1), .high(0), .low(0)) bits_60 (
        .y(_T_1),
        .in(reset)
    );
    wire _T_2;
    BITWISEOR #(.width(1)) bitwiseor_61 (
        .y(_T_2),
        .a(_T),
        .b(_T_1)
    );
    wire _T_3;
    EQ_UNSIGNED #(.width(1)) u_eq_62 (
        .y(_T_3),
        .a(_T_2),
        .b(1'h0)
    );
    wire _T_4;
    wire [11:0] _WTEMP_19;
    PAD_SIGNED #(.width(4), .n(12)) s_pad_63 (
        .y(_WTEMP_19),
        .in(4'sh5)
    );
    EQ_SIGNED #(.width(12)) s_eq_64 (
        .y(_T_4),
        .a(sIntResult),
        .b(_WTEMP_19)
    );
    wire _T_5;
    BITS #(.width(1), .high(0), .low(0)) bits_65 (
        .y(_T_5),
        .in(reset)
    );
    wire _T_6;
    BITWISEOR #(.width(1)) bitwiseor_66 (
        .y(_T_6),
        .a(_T_4),
        .b(_T_5)
    );
    wire _T_7;
    EQ_UNSIGNED #(.width(1)) u_eq_67 (
        .y(_T_7),
        .a(_T_6),
        .b(1'h0)
    );
    wire [11:0] _T_8;
    ASUINT #(.width(12)) asuint_68 (
        .y(_T_8),
        .in(fixedResult)
    );
    wire _T_9;
    wire [11:0] _WTEMP_20;
    PAD_UNSIGNED #(.width(3), .n(12)) u_pad_69 (
        .y(_WTEMP_20),
        .in(3'h5)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_70 (
        .y(_T_9),
        .a(_T_8),
        .b(_WTEMP_20)
    );
    wire _T_10;
    BITS #(.width(1), .high(0), .low(0)) bits_71 (
        .y(_T_10),
        .in(reset)
    );
    wire _T_11;
    BITWISEOR #(.width(1)) bitwiseor_72 (
        .y(_T_11),
        .a(_T_9),
        .b(_T_10)
    );
    wire _T_12;
    EQ_UNSIGNED #(.width(1)) u_eq_73 (
        .y(_T_12),
        .a(_T_11),
        .b(1'h0)
    );
    wire [3:0] _node_21;
    ASSINT #(.width(4)) assint_74 (
        .y(_node_21),
        .in(4'h5)
    );
    wire _T_13;
    wire [4:0] _WTEMP_21;
    PAD_SIGNED #(.width(4), .n(5)) s_pad_75 (
        .y(_WTEMP_21),
        .in(_node_21)
    );
    EQ_SIGNED #(.width(5)) s_eq_76 (
        .y(_T_13),
        .a(intervalResult1),
        .b(_WTEMP_21)
    );
    wire _T_14;
    BITS #(.width(1), .high(0), .low(0)) bits_77 (
        .y(_T_14),
        .in(reset)
    );
    wire _T_15;
    BITWISEOR #(.width(1)) bitwiseor_78 (
        .y(_T_15),
        .a(_T_13),
        .b(_T_14)
    );
    wire _T_16;
    EQ_UNSIGNED #(.width(1)) u_eq_79 (
        .y(_T_16),
        .a(_T_15),
        .b(1'h0)
    );
    wire [3:0] _node_22;
    ASSINT #(.width(4)) assint_80 (
        .y(_node_22),
        .in(4'h5)
    );
    wire _T_17;
    wire [4:0] _WTEMP_22;
    PAD_SIGNED #(.width(4), .n(5)) s_pad_81 (
        .y(_WTEMP_22),
        .in(_node_22)
    );
    EQ_SIGNED #(.width(5)) s_eq_82 (
        .y(_T_17),
        .a(intervalResult2),
        .b(_WTEMP_22)
    );
    wire _T_18;
    BITS #(.width(1), .high(0), .low(0)) bits_83 (
        .y(_T_18),
        .in(reset)
    );
    wire _T_19;
    BITWISEOR #(.width(1)) bitwiseor_84 (
        .y(_T_19),
        .a(_T_17),
        .b(_T_18)
    );
    wire _T_20;
    EQ_UNSIGNED #(.width(1)) u_eq_85 (
        .y(_T_20),
        .a(_T_19),
        .b(1'h0)
    );
    wire _T_21;
    BITS #(.width(1), .high(0), .low(0)) bits_86 (
        .y(_T_21),
        .in(reset)
    );
    wire _T_22;
    EQ_UNSIGNED #(.width(1)) u_eq_87 (
        .y(_T_22),
        .a(_T_21),
        .b(1'h0)
    );
    assign fixedResult = _fixedResult_T_5;
    wire [4:0] _WTEMP_23;
    BITS #(.width(12), .high(4), .low(0)) bits_88 (
        .y(_WTEMP_23),
        .in(_intervalResult1_T_5)
    );
    ASSINT #(.width(5)) assint_89 (
        .y(intervalResult1),
        .in(_WTEMP_23)
    );
    wire [4:0] _WTEMP_24;
    BITS #(.width(12), .high(4), .low(0)) bits_90 (
        .y(_WTEMP_24),
        .in(_intervalResult2_T_5)
    );
    ASSINT #(.width(5)) assint_91 (
        .y(intervalResult2),
        .in(_WTEMP_24)
    );
    assign sIntResult = 12'sh5;
    assign uIntResult = 11'h5;
endmodule //IntervalChainedSubTester
module ASSINT(y, in);
    parameter width = 4;
    output [width-1:0] y;
    input [width-1:0] in;
    assign y = $signed(in);
endmodule // ASSINT
module PAD_SIGNED(y, in);
    parameter width = 4;
    parameter n = 4;
    output [(n > width ? n : width)-1:0] y;
    input [width-1:0] in;
    assign y = n > width ? {{(n - width){in[width-1]}}, in} : in;
endmodule // PAD_SIGNED
module SUB_SIGNED(y, a, b);
    parameter width = 4;
    output [width:0] y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = $signed(a) - $signed(b);
endmodule // SUB_SIGNED
module PAD_UNSIGNED(y, in);
    parameter width = 4;
    parameter n = 4;
    output [(n > width ? n : width)-1:0] y;
    input [width-1:0] in;
    assign y = (n > width) ? {{(n - width){1'b0}}, in} : in;
endmodule // PAD_UNSIGNED
module EQ_UNSIGNED(y, a, b);
    parameter width = 4;
    output y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a == b;
endmodule // EQ_UNSIGNED
module BITS(y, in);
    parameter width = 4;
    parameter high = 2;
    parameter low = 0;
    output [high-low:0] y;
    input [width-1:0] in;
    assign y = in[high:low];
endmodule // BITS
module BITWISEOR(y, a, b);
    parameter width = 4;
    output [width-1:0] y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a | b;
endmodule // BITWISEOR
module EQ_SIGNED(y, a, b);
    parameter width = 4;
    output y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = $signed(a) == $signed(b);
endmodule // EQ_SIGNED
module ASUINT(y, in);
    parameter width = 4;
    output [width-1:0] y;
    input [width-1:0] in;
    assign y = $unsigned(in);
endmodule // ASUINT
