module HardwareHashMaker(
  input         clock,
  input         reset,
  input  [63:0] io_x_0,
  input  [63:0] io_x_1,
  input  [63:0] io_x_2,
  input  [63:0] io_x_3,
  output [63:0] io_out
);
  wire [127:0] _T_31 = $signed(io_x_0) * 64'shcd72ce8f; // @[HardwareHashMaker.scala 71:18]
  wire [128:0] _T_32 = {{1{_T_31[127]}},_T_31}; // @[HardwareHashMaker.scala 71:13]
  wire [127:0] _T_34 = _T_32[127:0]; // @[HardwareHashMaker.scala 71:13]
  wire [127:0] _T_35 = $signed(io_x_1) * -64'she6cbb976; // @[HardwareHashMaker.scala 71:18]
  wire [127:0] _T_38 = $signed(_T_34) + $signed(_T_35); // @[HardwareHashMaker.scala 71:13]
  wire [127:0] _T_39 = $signed(io_x_2) * 64'sh214b73994; // @[HardwareHashMaker.scala 71:18]
  wire [127:0] _T_42 = $signed(_T_38) + $signed(_T_39); // @[HardwareHashMaker.scala 71:13]
  wire [127:0] _T_43 = $signed(io_x_3) * 64'shc3867b28; // @[HardwareHashMaker.scala 71:18]
  wire [127:0] _T_46 = $signed(_T_42) + $signed(_T_43); // @[HardwareHashMaker.scala 71:13]
  wire [128:0] _T_47 = {{1{_T_46[127]}},_T_46}; // @[HardwareHashMaker.scala 74:10]
  wire [127:0] _T_49 = _T_47[127:0]; // @[HardwareHashMaker.scala 74:10]
  wire [101:0] _T_50 = _T_49[127:26]; // @[HardwareHashMaker.scala 74:34]
  wire [127:0] _T_52 = $signed(io_x_0) * 64'shfc0d139b; // @[HardwareHashMaker.scala 71:18]
  wire [128:0] _T_53 = {{1{_T_52[127]}},_T_52}; // @[HardwareHashMaker.scala 71:13]
  wire [127:0] _T_55 = _T_53[127:0]; // @[HardwareHashMaker.scala 71:13]
  wire [127:0] _T_56 = $signed(io_x_1) * -64'sh1aef41b15; // @[HardwareHashMaker.scala 71:18]
  wire [127:0] _T_59 = $signed(_T_55) + $signed(_T_56); // @[HardwareHashMaker.scala 71:13]
  wire [127:0] _T_60 = $signed(io_x_2) * -64'sh6fc7ea3; // @[HardwareHashMaker.scala 71:18]
  wire [127:0] _T_63 = $signed(_T_59) + $signed(_T_60); // @[HardwareHashMaker.scala 71:13]
  wire [127:0] _T_64 = $signed(io_x_3) * 64'sh1d80be0d; // @[HardwareHashMaker.scala 71:18]
  wire [127:0] _T_67 = $signed(_T_63) + $signed(_T_64); // @[HardwareHashMaker.scala 71:13]
  wire [128:0] _T_68 = {{1{_T_67[127]}},_T_67}; // @[HardwareHashMaker.scala 74:10]
  wire [127:0] _T_70 = _T_68[127:0]; // @[HardwareHashMaker.scala 74:10]
  wire [101:0] _T_71 = _T_70[127:26]; // @[HardwareHashMaker.scala 74:34]
  wire [127:0] _T_73 = $signed(io_x_0) * -64'sh63e1fcbb; // @[HardwareHashMaker.scala 71:18]
  wire [128:0] _T_74 = {{1{_T_73[127]}},_T_73}; // @[HardwareHashMaker.scala 71:13]
  wire [127:0] _T_76 = _T_74[127:0]; // @[HardwareHashMaker.scala 71:13]
  wire [127:0] _T_77 = $signed(io_x_1) * -64'sha4b52117; // @[HardwareHashMaker.scala 71:18]
  wire [127:0] _T_80 = $signed(_T_76) + $signed(_T_77); // @[HardwareHashMaker.scala 71:13]
  wire [127:0] _T_81 = $signed(io_x_2) * 64'shd6e13f9; // @[HardwareHashMaker.scala 71:18]
  wire [127:0] _T_84 = $signed(_T_80) + $signed(_T_81); // @[HardwareHashMaker.scala 71:13]
  wire [127:0] _T_85 = $signed(io_x_3) * 64'sh8576aca2; // @[HardwareHashMaker.scala 71:18]
  wire [127:0] _T_88 = $signed(_T_84) + $signed(_T_85); // @[HardwareHashMaker.scala 71:13]
  wire [128:0] _T_89 = {{1{_T_88[127]}},_T_88}; // @[HardwareHashMaker.scala 74:10]
  wire [127:0] _T_91 = _T_89[127:0]; // @[HardwareHashMaker.scala 74:10]
  wire [101:0] _T_92 = _T_91[127:26]; // @[HardwareHashMaker.scala 74:34]
  wire [127:0] _T_94 = $signed(io_x_0) * -64'shd2ef8062; // @[HardwareHashMaker.scala 71:18]
  wire [128:0] _T_95 = {{1{_T_94[127]}},_T_94}; // @[HardwareHashMaker.scala 71:13]
  wire [127:0] _T_97 = _T_95[127:0]; // @[HardwareHashMaker.scala 71:13]
  wire [127:0] _T_98 = $signed(io_x_1) * 64'sh42be6d75; // @[HardwareHashMaker.scala 71:18]
  wire [127:0] _T_101 = $signed(_T_97) + $signed(_T_98); // @[HardwareHashMaker.scala 71:13]
  wire [127:0] _T_102 = $signed(io_x_2) * -64'sh73f7016d; // @[HardwareHashMaker.scala 71:18]
  wire [127:0] _T_105 = $signed(_T_101) + $signed(_T_102); // @[HardwareHashMaker.scala 71:13]
  wire [127:0] _T_106 = $signed(io_x_3) * 64'sh16734aab4; // @[HardwareHashMaker.scala 71:18]
  wire [127:0] _T_109 = $signed(_T_105) + $signed(_T_106); // @[HardwareHashMaker.scala 71:13]
  wire [128:0] _T_110 = {{1{_T_109[127]}},_T_109}; // @[HardwareHashMaker.scala 74:10]
  wire [127:0] _T_112 = _T_110[127:0]; // @[HardwareHashMaker.scala 74:10]
  wire [101:0] _T_113 = _T_112[127:26]; // @[HardwareHashMaker.scala 74:34]
  wire [127:0] _T_115 = $signed(io_x_0) * 64'sh4568d0ed; // @[HardwareHashMaker.scala 71:18]
  wire [128:0] _T_116 = {{1{_T_115[127]}},_T_115}; // @[HardwareHashMaker.scala 71:13]
  wire [127:0] _T_118 = _T_116[127:0]; // @[HardwareHashMaker.scala 71:13]
  wire [127:0] _T_119 = $signed(io_x_1) * -64'sh1ce4abd; // @[HardwareHashMaker.scala 71:18]
  wire [127:0] _T_122 = $signed(_T_118) + $signed(_T_119); // @[HardwareHashMaker.scala 71:13]
  wire [127:0] _T_123 = $signed(io_x_2) * 64'she7ab5f92; // @[HardwareHashMaker.scala 71:18]
  wire [127:0] _T_126 = $signed(_T_122) + $signed(_T_123); // @[HardwareHashMaker.scala 71:13]
  wire [127:0] _T_127 = $signed(io_x_3) * 64'shdb5acccd; // @[HardwareHashMaker.scala 71:18]
  wire [127:0] _T_130 = $signed(_T_126) + $signed(_T_127); // @[HardwareHashMaker.scala 71:13]
  wire [128:0] _T_131 = {{1{_T_130[127]}},_T_130}; // @[HardwareHashMaker.scala 74:10]
  wire [127:0] _T_133 = _T_131[127:0]; // @[HardwareHashMaker.scala 74:10]
  wire [101:0] _T_134 = _T_133[127:26]; // @[HardwareHashMaker.scala 74:34]
  wire [101:0] _T_137 = $signed(_T_50) + $signed(_T_71); // @[HardwareHashMaker.scala 78:39]
  wire [101:0] _T_140 = $signed(_T_137) + $signed(_T_92); // @[HardwareHashMaker.scala 78:39]
  wire [101:0] _T_143 = $signed(_T_140) + $signed(_T_113); // @[HardwareHashMaker.scala 78:39]
  wire [101:0] _T_146 = $signed(_T_143) + $signed(_T_134); // @[HardwareHashMaker.scala 78:39]
  wire [95:0] _GEN_0 = _T_146[101:6]; // @[HardwareHashMaker.scala 78:10]
  assign io_out = _GEN_0[63:0]; // @[HardwareHashMaker.scala 78:10]
endmodule
