module CoreTester(
    input clock,
    input reset
);
    wire _dut__clock;
    wire _dut__reset;
    wire _dut__io_host_fromhost_valid;
    wire [31:0] _dut__io_host_fromhost_bits;
    wire [31:0] _dut__io_host_tohost;
    wire _dut__io_icache_abort;
    wire _dut__io_icache_req_valid;
    wire [31:0] _dut__io_icache_req_bits_addr;
    wire [31:0] _dut__io_icache_req_bits_data;
    wire [3:0] _dut__io_icache_req_bits_mask;
    wire _dut__io_icache_resp_valid;
    wire [31:0] _dut__io_icache_resp_bits_data;
    wire _dut__io_dcache_abort;
    wire _dut__io_dcache_req_valid;
    wire [31:0] _dut__io_dcache_req_bits_addr;
    wire [31:0] _dut__io_dcache_req_bits_data;
    wire [3:0] _dut__io_dcache_req_bits_mask;
    wire _dut__io_dcache_resp_valid;
    wire [31:0] _dut__io_dcache_resp_bits_data;
    Core dut (
        .clock(_dut__clock),
        .reset(_dut__reset),
        .io_host_fromhost_valid(_dut__io_host_fromhost_valid),
        .io_host_fromhost_bits(_dut__io_host_fromhost_bits),
        .io_host_tohost(_dut__io_host_tohost),
        .io_icache_abort(_dut__io_icache_abort),
        .io_icache_req_valid(_dut__io_icache_req_valid),
        .io_icache_req_bits_addr(_dut__io_icache_req_bits_addr),
        .io_icache_req_bits_data(_dut__io_icache_req_bits_data),
        .io_icache_req_bits_mask(_dut__io_icache_req_bits_mask),
        .io_icache_resp_valid(_dut__io_icache_resp_valid),
        .io_icache_resp_bits_data(_dut__io_icache_resp_bits_data),
        .io_dcache_abort(_dut__io_dcache_abort),
        .io_dcache_req_valid(_dut__io_dcache_req_valid),
        .io_dcache_req_bits_addr(_dut__io_dcache_req_bits_addr),
        .io_dcache_req_bits_data(_dut__io_dcache_req_bits_data),
        .io_dcache_req_bits_mask(_dut__io_dcache_req_bits_mask),
        .io_dcache_resp_valid(_dut__io_dcache_resp_valid),
        .io_dcache_resp_bits_data(_dut__io_dcache_resp_bits_data)
    );
    wire [31:0] imem__T_385_data;
    wire imem__T_385_clk;
    wire imem__T_385_en;
    wire [19:0] imem__T_385_addr;
    wire imem__T_402_clk;
    wire imem__T_402_en;
    wire imem__T_402_mask;
    wire [19:0] imem__T_402_addr;
    wire [31:0] imem__T_402_data;
    RAMMEM #(.depth(1048576), .addrbits(20), .width(32), .isSyncRead(0)) imem (
        .read_data(imem__T_385_data),
        .read_clk(imem__T_385_clk),
        .read_en(imem__T_385_en),
        .read_addr(imem__T_385_addr),
        .write_clk(imem__T_402_clk),
        .write_en(imem__T_402_en),
        .write_mask(imem__T_402_mask),
        .write_addr(imem__T_402_addr),
        .write_data(imem__T_402_data)
    );
    wire [31:0] dmem__T_349_data;
    wire dmem__T_349_clk;
    wire dmem__T_349_en;
    wire [19:0] dmem__T_349_addr;
    wire [31:0] dmem__T_358_data;
    wire dmem__T_358_clk;
    wire dmem__T_358_en;
    wire [19:0] dmem__T_358_addr;
    wire [31:0] dmem__T_367_data;
    wire dmem__T_367_clk;
    wire dmem__T_367_en;
    wire [19:0] dmem__T_367_addr;
    wire [31:0] dmem__T_376_data;
    wire dmem__T_376_clk;
    wire dmem__T_376_en;
    wire [19:0] dmem__T_376_addr;
    wire [31:0] dmem__T_388_data;
    wire dmem__T_388_clk;
    wire dmem__T_388_en;
    wire [19:0] dmem__T_388_addr;
    wire dmem__T_403_clk;
    wire dmem__T_403_en;
    wire dmem__T_403_mask;
    wire [19:0] dmem__T_403_addr;
    wire [31:0] dmem__T_403_data;
    wire dmem__T_408_clk;
    wire dmem__T_408_en;
    wire dmem__T_408_mask;
    wire [19:0] dmem__T_408_addr;
    wire [31:0] dmem__T_408_data;
    wire [159:0] dmem_read_datas;
    wire [4:0] dmem_read_clks;
    wire [4:0] dmem_read_ens;
    wire [99:0] dmem_read_addrs;
    wire [1:0] dmem_write_clks;
    wire [1:0] dmem_write_ens;
    wire [1:0] dmem_write_masks;
    wire [39:0] dmem_write_addrs;
    wire [63:0] dmem_write_datas;
    BITS #(.width(160), .high(31), .low(0)) bits_1878 (
        .y(dmem__T_349_data),
        .in(dmem_read_datas)
    );
    BITS #(.width(160), .high(63), .low(32)) bits_1879 (
        .y(dmem__T_358_data),
        .in(dmem_read_datas)
    );
    BITS #(.width(160), .high(95), .low(64)) bits_1880 (
        .y(dmem__T_367_data),
        .in(dmem_read_datas)
    );
    BITS #(.width(160), .high(127), .low(96)) bits_1881 (
        .y(dmem__T_376_data),
        .in(dmem_read_datas)
    );
    BITS #(.width(160), .high(159), .low(128)) bits_1882 (
        .y(dmem__T_388_data),
        .in(dmem_read_datas)
    );
    wire [1:0] _WTEMP_182;
    CAT #(.width_a(1), .width_b(1)) cat_1883 (
        .y(_WTEMP_182),
        .a(dmem__T_388_clk),
        .b(dmem__T_376_clk)
    );
    wire [2:0] _WTEMP_183;
    CAT #(.width_a(2), .width_b(1)) cat_1884 (
        .y(_WTEMP_183),
        .a(_WTEMP_182),
        .b(dmem__T_367_clk)
    );
    wire [3:0] _WTEMP_184;
    CAT #(.width_a(3), .width_b(1)) cat_1885 (
        .y(_WTEMP_184),
        .a(_WTEMP_183),
        .b(dmem__T_358_clk)
    );
    CAT #(.width_a(4), .width_b(1)) cat_1886 (
        .y(dmem_read_clks),
        .a(_WTEMP_184),
        .b(dmem__T_349_clk)
    );
    wire [1:0] _WTEMP_185;
    CAT #(.width_a(1), .width_b(1)) cat_1887 (
        .y(_WTEMP_185),
        .a(dmem__T_388_en),
        .b(dmem__T_376_en)
    );
    wire [2:0] _WTEMP_186;
    CAT #(.width_a(2), .width_b(1)) cat_1888 (
        .y(_WTEMP_186),
        .a(_WTEMP_185),
        .b(dmem__T_367_en)
    );
    wire [3:0] _WTEMP_187;
    CAT #(.width_a(3), .width_b(1)) cat_1889 (
        .y(_WTEMP_187),
        .a(_WTEMP_186),
        .b(dmem__T_358_en)
    );
    CAT #(.width_a(4), .width_b(1)) cat_1890 (
        .y(dmem_read_ens),
        .a(_WTEMP_187),
        .b(dmem__T_349_en)
    );
    wire [39:0] _WTEMP_188;
    CAT #(.width_a(20), .width_b(20)) cat_1891 (
        .y(_WTEMP_188),
        .a(dmem__T_388_addr),
        .b(dmem__T_376_addr)
    );
    wire [59:0] _WTEMP_189;
    CAT #(.width_a(40), .width_b(20)) cat_1892 (
        .y(_WTEMP_189),
        .a(_WTEMP_188),
        .b(dmem__T_367_addr)
    );
    wire [79:0] _WTEMP_190;
    CAT #(.width_a(60), .width_b(20)) cat_1893 (
        .y(_WTEMP_190),
        .a(_WTEMP_189),
        .b(dmem__T_358_addr)
    );
    CAT #(.width_a(80), .width_b(20)) cat_1894 (
        .y(dmem_read_addrs),
        .a(_WTEMP_190),
        .b(dmem__T_349_addr)
    );
    CAT #(.width_a(32), .width_b(32)) cat_1895 (
        .y(dmem_write_datas),
        .a(dmem__T_408_data),
        .b(dmem__T_403_data)
    );
    CAT #(.width_a(1), .width_b(1)) cat_1896 (
        .y(dmem_write_clks),
        .a(dmem__T_408_clk),
        .b(dmem__T_403_clk)
    );
    CAT #(.width_a(1), .width_b(1)) cat_1897 (
        .y(dmem_write_ens),
        .a(dmem__T_408_en),
        .b(dmem__T_403_en)
    );
    CAT #(.width_a(20), .width_b(20)) cat_1898 (
        .y(dmem_write_addrs),
        .a(dmem__T_408_addr),
        .b(dmem__T_403_addr)
    );
    CAT #(.width_a(1), .width_b(1)) cat_1899 (
        .y(dmem_write_masks),
        .a(dmem__T_408_mask),
        .b(dmem__T_403_mask)
    );
    MRMWMEM #(.depth(1048576), .addrbits(20), .width(32), .readernum(5), .writernum(2), .isSyncRead(0)) dmem (
        .read_datas(dmem_read_datas),
        .read_clks(dmem_read_clks),
        .read_ens(dmem_read_ens),
        .read_addrs(dmem_read_addrs),
        .write_clks(dmem_write_clks),
        .write_ens(dmem_write_ens),
        .write_masks(dmem_write_masks),
        .write_addrs(dmem_write_addrs),
        .write_datas(dmem_write_datas)
    );
    wire _state__q;
    wire _state__d;
    DFF_POSCLK #(.width(1)) state (
        .q(_state__q),
        .d(_state__d),
        .clk(clock)
    );
    wire [31:0] _cycle__q;
    wire [31:0] _cycle__d;
    DFF_POSCLK #(.width(32)) cycle (
        .q(_cycle__q),
        .d(_cycle__d),
        .clk(clock)
    );
    wire [7:0] _cntr__q;
    wire [7:0] _cntr__d;
    DFF_POSCLK #(.width(8)) cntr (
        .q(_cntr__q),
        .d(_cntr__d),
        .clk(clock)
    );
    wire [31:0] __T_386__q;
    wire [31:0] __T_386__d;
    DFF_POSCLK #(.width(32)) _T_386 (
        .q(__T_386__q),
        .d(__T_386__d),
        .clk(clock)
    );
    wire [31:0] __T_389__q;
    wire [31:0] __T_389__d;
    DFF_POSCLK #(.width(32)) _T_389 (
        .q(__T_389__q),
        .d(__T_389__d),
        .clk(clock)
    );
    wire [63:0] _T_164;
    assign _T_164 = 64'h10101464C457F;
    wire [63:0] _T_165;
    assign _T_165 = 64'hF3000200000000;
    wire [95:0] _T_166;
    assign _T_166 = 96'hF300020000000000000000;
    wire [159:0] _T_167;
    assign _T_167 = 160'hF30002000000000000000000010101464C457F;
    wire [63:0] _T_168;
    assign _T_168 = 64'h10000000001;
    wire [63:0] _T_169;
    assign _T_169 = 64'h454;
    wire [95:0] _T_170;
    assign _T_170 = 96'h45400000034;
    wire [159:0] _T_171;
    assign _T_171 = 160'h454000000340000010000000001;
    wire [319:0] _T_172;
    assign _T_172 = 320'h45400000034000001000000000100F30002000000000000000000010101464C457F;
    wire [63:0] _T_173;
    assign _T_173 = 64'h28000100200034;
    wire [63:0] _T_174;
    assign _T_174 = 64'h1;
    wire [95:0] _T_175;
    assign _T_175 = 96'h100020005;
    wire [159:0] _T_176;
    assign _T_176 = 160'h1000200050028000100200034;
    wire [63:0] _T_177;
    assign _T_177 = 64'h0;
    wire [63:0] _T_178;
    assign _T_178 = 64'h500000260;
    wire [95:0] _T_179;
    assign _T_179 = 96'h50000026000000260;
    wire [159:0] _T_180;
    assign _T_180 = 160'h500000260000002600000000000000000;
    wire [319:0] _T_181;
    assign _T_181 = 320'h5000002600000026000000000000000000000000000000001000200050028000100200034;
    wire [639:0] _T_182;
    assign _T_182 = 640'h5000002600000026000000000000000000000000000000001000200050028000100200034000000000000045400000034000001000000000100F30002000000000000000000010101464C457F;
    wire [63:0] _T_183;
    assign _T_183 = 64'h2000;
    wire [63:0] _T_184;
    assign _T_184 = 64'h0;
    wire [95:0] _T_185;
    assign _T_185 = 96'h0;
    wire [159:0] _T_186;
    assign _T_186 = 160'h2000;
    wire [63:0] _T_187;
    assign _T_187 = 64'h0;
    wire [63:0] _T_188;
    assign _T_188 = 64'h0;
    wire [95:0] _T_189;
    assign _T_189 = 96'h0;
    wire [159:0] _T_190;
    assign _T_190 = 160'h0;
    wire [319:0] _T_191;
    assign _T_191 = 320'h2000;
    wire [63:0] _T_192;
    assign _T_192 = 64'h0;
    wire [63:0] _T_193;
    assign _T_193 = 64'h0;
    wire [95:0] _T_194;
    assign _T_194 = 96'h0;
    wire [159:0] _T_195;
    assign _T_195 = 160'h0;
    wire [63:0] _T_196;
    assign _T_196 = 64'h0;
    wire [63:0] _T_197;
    assign _T_197 = 64'h0;
    wire [95:0] _T_198;
    assign _T_198 = 96'h0;
    wire [159:0] _T_199;
    assign _T_199 = 160'h0;
    wire [319:0] _T_200;
    assign _T_200 = 320'h0;
    wire [639:0] _T_201;
    assign _T_201 = 640'h2000;
    wire [1279:0] _T_202;
    assign _T_202 = 1280'h200000000005000002600000026000000000000000000000000000000001000200050028000100200034000000000000045400000034000001000000000100F30002000000000000000000010101464C457F;
    wire [63:0] _T_203;
    assign _T_203 = 64'h0;
    wire [63:0] _T_204;
    assign _T_204 = 64'h0;
    wire [95:0] _T_205;
    assign _T_205 = 96'h0;
    wire [159:0] _T_206;
    assign _T_206 = 160'h0;
    wire [63:0] _T_207;
    assign _T_207 = 64'h0;
    wire [63:0] _T_208;
    assign _T_208 = 64'h0;
    wire [95:0] _T_209;
    assign _T_209 = 96'h0;
    wire [159:0] _T_210;
    assign _T_210 = 160'h0;
    wire [319:0] _T_211;
    assign _T_211 = 320'h0;
    wire [63:0] _T_212;
    assign _T_212 = 64'h0;
    wire [63:0] _T_213;
    assign _T_213 = 64'h0;
    wire [95:0] _T_214;
    assign _T_214 = 96'h0;
    wire [159:0] _T_215;
    assign _T_215 = 160'h0;
    wire [63:0] _T_216;
    assign _T_216 = 64'h0;
    wire [63:0] _T_217;
    assign _T_217 = 64'h0;
    wire [95:0] _T_218;
    assign _T_218 = 96'h0;
    wire [159:0] _T_219;
    assign _T_219 = 160'h0;
    wire [319:0] _T_220;
    assign _T_220 = 320'h0;
    wire [639:0] _T_221;
    assign _T_221 = 640'h0;
    wire [63:0] _T_222;
    assign _T_222 = 64'h0;
    wire [63:0] _T_223;
    assign _T_223 = 64'hF1700000000;
    wire [95:0] _T_224;
    assign _T_224 = 96'hF170000000000000000;
    wire [159:0] _T_225;
    assign _T_225 = 160'hF1700000000000000000000000000000000;
    wire [63:0] _T_226;
    assign _T_226 = 64'h34102FF3158F0F13;
    wire [63:0] _T_227;
    assign _T_227 = 64'hEF0F0F1300000F17;
    wire [95:0] _T_228;
    assign _T_228 = 96'hEF0F0F1300000F1707FF0C63;
    wire [159:0] _T_229;
    assign _T_229 = 160'hEF0F0F1300000F1707FF0C6334102FF3158F0F13;
    wire [319:0] _T_230;
    assign _T_230 = 320'hEF0F0F1300000F1707FF0C6334102FF3158F0F1300000F1700000000000000000000000000000000;
    wire [63:0] _T_231;
    assign _T_231 = 64'hF17020F1863;
    wire [63:0] _T_232;
    assign _T_232 = 64'hED9FF06F000F0463;
    wire [95:0] _T_233;
    assign _T_233 = 96'hED9FF06F000F0463EE4F0F13;
    wire [159:0] _T_234;
    assign _T_234 = 160'hED9FF06F000F0463EE4F0F1300000F17020F1863;
    wire [63:0] _T_235;
    assign _T_235 = 64'h130540006F;
    wire [63:0] _T_236;
    assign _T_236 = 64'h1300000013;
    wire [95:0] _T_237;
    assign _T_237 = 96'h130000001300000013;
    wire [159:0] _T_238;
    assign _T_238 = 160'h130000001300000013000000130540006F;
    wire [319:0] _T_239;
    assign _T_239 = 320'h130000001300000013000000130540006FED9FF06F000F0463EE4F0F1300000F17020F1863;
    wire [639:0] _T_240;
    assign _T_240 = 640'h130000001300000013000000130540006FED9FF06F000F0463EE4F0F1300000F17020F1863EF0F0F1300000F1707FF0C6334102FF3158F0F1300000F1700000000000000000000000000000000;
    wire [1279:0] _T_241;
    assign _T_241 = 1280'h130000001300000013000000130540006FED9FF06F000F0463EE4F0F1300000F17020F1863EF0F0F1300000F1707FF0C6334102FF3158F0F1300000F17000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [2559:0] _T_242;
    assign _T_242 = 2560'h130000001300000013000000130540006FED9FF06F000F0463EE4F0F1300000F17020F1863EF0F0F1300000F1707FF0C6334102FF3158F0F1300000F17000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000200000000005000002600000026000000000000000000000000000000001000200050028000100200034000000000000045400000034000001000000000100F30002000000000000000000010101464C457F;
    wire [63:0] _T_243;
    assign _T_243 = 64'hFA0F5EE334202F73;
    wire [63:0] _T_244;
    assign _T_244 = 64'h1300000013;
    wire [95:0] _T_245;
    assign _T_245 = 96'h130000001330500073;
    wire [159:0] _T_246;
    assign _T_246 = 160'h130000001330500073FA0F5EE334202F73;
    wire [63:0] _T_247;
    assign _T_247 = 64'h1300000013;
    wire [63:0] _T_248;
    assign _T_248 = 64'h1300000013;
    wire [95:0] _T_249;
    assign _T_249 = 96'h130000001300000013;
    wire [159:0] _T_250;
    assign _T_250 = 160'h1300000013000000130000001300000013;
    wire [319:0] _T_251;
    assign _T_251 = 320'h1300000013000000130000001300000013000000130000001330500073FA0F5EE334202F73;
    wire [63:0] _T_252;
    assign _T_252 = 64'h1300000013;
    wire [63:0] _T_253;
    assign _T_253 = 64'h1300000013;
    wire [95:0] _T_254;
    assign _T_254 = 96'h130000001300000013;
    wire [159:0] _T_255;
    assign _T_255 = 160'h1300000013000000130000001300000013;
    wire [63:0] _T_256;
    assign _T_256 = 64'h539E6E1300000013;
    wire [63:0] _T_257;
    assign _T_257 = 64'h13FFDFF06F;
    wire [95:0] _T_258;
    assign _T_258 = 96'h13FFDFF06F780E1073;
    wire [159:0] _T_259;
    assign _T_259 = 160'h13FFDFF06F780E1073539E6E1300000013;
    wire [319:0] _T_260;
    assign _T_260 = 320'h13FFDFF06F780E1073539E6E13000000130000001300000013000000130000001300000013;
    wire [639:0] _T_261;
    assign _T_261 = 640'h13FFDFF06F780E1073539E6E130000001300000013000000130000001300000013000000130000001300000013000000130000001300000013000000130000001330500073FA0F5EE334202F73;
    wire [63:0] _T_262;
    assign _T_262 = 64'h1300000013;
    wire [63:0] _T_263;
    assign _T_263 = 64'h1300000013;
    wire [95:0] _T_264;
    assign _T_264 = 96'h130000001300000013;
    wire [159:0] _T_265;
    assign _T_265 = 160'h1300000013000000130000001300000013;
    wire [63:0] _T_266;
    assign _T_266 = 64'h1300000013;
    wire [63:0] _T_267;
    assign _T_267 = 64'h1300000013;
    wire [95:0] _T_268;
    assign _T_268 = 96'h130000001300000013;
    wire [159:0] _T_269;
    assign _T_269 = 160'h1300000013000000130000001300000013;
    wire [319:0] _T_270;
    assign _T_270 = 320'h13000000130000001300000013000000130000001300000013000000130000001300000013;
    wire [63:0] _T_271;
    assign _T_271 = 64'h1300000013;
    wire [63:0] _T_272;
    assign _T_272 = 64'h34102FF3098F0F13;
    wire [95:0] _T_273;
    assign _T_273 = 96'h34102FF3098F0F1300000F17;
    wire [159:0] _T_274;
    assign _T_274 = 160'h34102FF3098F0F1300000F170000001300000013;
    wire [63:0] _T_275;
    assign _T_275 = 64'hF17FBFF0CE3;
    wire [63:0] _T_276;
    assign _T_276 = 64'hE25FF06F000F0463;
    wire [95:0] _T_277;
    assign _T_277 = 96'hE25FF06F000F0463E30F0F13;
    wire [159:0] _T_278;
    assign _T_278 = 160'hE25FF06F000F0463E30F0F1300000F17FBFF0CE3;
    wire [319:0] _T_279;
    assign _T_279 = 320'hE25FF06F000F0463E30F0F1300000F17FBFF0CE334102FF3098F0F1300000F170000001300000013;
    wire [639:0] _T_280;
    assign _T_280 = 640'hE25FF06F000F0463E30F0F1300000F17FBFF0CE334102FF3098F0F1300000F17000000130000001300000013000000130000001300000013000000130000001300000013000000130000001300000013;
    wire [1279:0] _T_281;
    assign _T_281 = 1280'hE25FF06F000F0463E30F0F1300000F17FBFF0CE334102FF3098F0F1300000F1700000013000000130000001300000013000000130000001300000013000000130000001300000013000000130000001300000013FFDFF06F780E1073539E6E130000001300000013000000130000001300000013000000130000001300000013000000130000001300000013000000130000001330500073FA0F5EE334202F73;
    wire [63:0] _T_282;
    assign _T_282 = 64'h13FA1FF06F;
    wire [63:0] _T_283;
    assign _T_283 = 64'h1300000013;
    wire [95:0] _T_284;
    assign _T_284 = 96'h130000001300000013;
    wire [159:0] _T_285;
    assign _T_285 = 160'h13000000130000001300000013FA1FF06F;
    wire [63:0] _T_286;
    assign _T_286 = 64'h1300000013;
    wire [63:0] _T_287;
    assign _T_287 = 64'h51063F1002573;
    wire [95:0] _T_288;
    assign _T_288 = 96'h51063F100257300000013;
    wire [159:0] _T_289;
    assign _T_289 = 160'h51063F1002573000000130000001300000013;
    wire [319:0] _T_290;
    assign _T_290 = 320'h51063F100257300000013000000130000001300000013000000130000001300000013FA1FF06F;
    wire [63:0] _T_291;
    assign _T_291 = 64'h55863F0002573;
    wire [63:0] _T_292;
    assign _T_292 = 64'h400006F00100E13;
    wire [95:0] _T_293;
    assign _T_293 = 96'h400006F00100E130FF0000F;
    wire [159:0] _T_294;
    assign _T_294 = 160'h400006F00100E130FF0000F00055863F0002573;
    wire [63:0] _T_295;
    assign _T_295 = 64'h29700000E13;
    wire [63:0] _T_296;
    assign _T_296 = 64'h1012907300028463;
    wire [95:0] _T_297;
    assign _T_297 = 96'h1012907300028463DE028293;
    wire [159:0] _T_298;
    assign _T_298 = 160'h1012907300028463DE0282930000029700000E13;
    wire [319:0] _T_299;
    assign _T_299 = 320'h1012907300028463DE0282930000029700000E130400006F00100E130FF0000F00055863F0002573;
    wire [639:0] _T_300;
    assign _T_300 = 640'h1012907300028463DE0282930000029700000E130400006F00100E130FF0000F00055863F000257300051063F100257300000013000000130000001300000013000000130000001300000013FA1FF06F;
    wire [63:0] _T_301;
    assign _T_301 = 64'h3002B0731F800293;
    wire [63:0] _T_302;
    assign _T_302 = 64'h3412907301428293;
    wire [95:0] _T_303;
    assign _T_303 = 96'h341290730142829300000297;
    wire [159:0] _T_304;
    assign _T_304 = 160'h3412907301428293000002973002B0731F800293;
    wire [63:0] _T_305;
    assign _T_305 = 64'h10000073F1002573;
    wire [63:0] _T_306;
    assign _T_306 = 64'h40006F00100E13;
    wire [95:0] _T_307;
    assign _T_307 = 96'h40006F00100E130FF0000F;
    wire [159:0] _T_308;
    assign _T_308 = 160'h40006F00100E130FF0000F10000073F1002573;
    wire [319:0] _T_309;
    assign _T_309 = 320'h40006F00100E130FF0000F10000073F10025733412907301428293000002973002B0731F800293;
    wire [63:0] _T_310;
    assign _T_310 = 64'hFFDFF06F00000073;
    wire [63:0] _T_311;
    assign _T_311 = 64'h0;
    wire [95:0] _T_312;
    assign _T_312 = 96'h0;
    wire [159:0] _T_313;
    assign _T_313 = 160'hFFDFF06F00000073;
    wire [63:0] _T_314;
    assign _T_314 = 64'h0;
    wire [63:0] _T_315;
    assign _T_315 = 64'h0;
    wire [95:0] _T_316;
    assign _T_316 = 96'h0;
    wire [159:0] _T_317;
    assign _T_317 = 160'h0;
    wire [319:0] _T_318;
    assign _T_318 = 320'hFFDFF06F00000073;
    wire [639:0] _T_319;
    assign _T_319 = 640'hFFDFF06F000000730040006F00100E130FF0000F10000073F10025733412907301428293000002973002B0731F800293;
    wire [1279:0] _T_320;
    assign _T_320 = 1280'hFFDFF06F000000730040006F00100E130FF0000F10000073F10025733412907301428293000002973002B0731F8002931012907300028463DE0282930000029700000E130400006F00100E130FF0000F00055863F000257300051063F100257300000013000000130000001300000013000000130000001300000013FA1FF06F;
    wire [2559:0] _T_321;
    assign _T_321 = 2560'hFFDFF06F000000730040006F00100E130FF0000F10000073F10025733412907301428293000002973002B0731F8002931012907300028463DE0282930000029700000E130400006F00100E130FF0000F00055863F000257300051063F100257300000013000000130000001300000013000000130000001300000013FA1FF06FE25FF06F000F0463E30F0F1300000F17FBFF0CE334102FF3098F0F1300000F1700000013000000130000001300000013000000130000001300000013000000130000001300000013000000130000001300000013FFDFF06F780E1073539E6E130000001300000013000000130000001300000013000000130000001300000013000000130000001300000013000000130000001330500073FA0F5EE334202F73;
    wire [5119:0] _T_322;
    assign _T_322 = 5120'hFFDFF06F000000730040006F00100E130FF0000F10000073F10025733412907301428293000002973002B0731F8002931012907300028463DE0282930000029700000E130400006F00100E130FF0000F00055863F000257300051063F100257300000013000000130000001300000013000000130000001300000013FA1FF06FE25FF06F000F0463E30F0F1300000F17FBFF0CE334102FF3098F0F1300000F1700000013000000130000001300000013000000130000001300000013000000130000001300000013000000130000001300000013FFDFF06F780E1073539E6E130000001300000013000000130000001300000013000000130000001300000013000000130000001300000013000000130000001330500073FA0F5EE334202F73000000130000001300000013000000130540006FED9FF06F000F0463EE4F0F1300000F17020F1863EF0F0F1300000F1707FF0C6334102FF3158F0F1300000F17000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000200000000005000002600000026000000000000000000000000000000001000200050028000100200034000000000000045400000034000001000000000100F30002000000000000000000010101464C457F;
    wire _T_336;
    EQ_UNSIGNED #(.width(1)) u_eq_1900 (
        .y(_T_336),
        .a(_state__q),
        .b(1'h0)
    );
    wire _T_339;
    EQ_UNSIGNED #(.width(8)) u_eq_1901 (
        .y(_T_339),
        .a(_cntr__q),
        .b(8'hFF)
    );
    wire [8:0] _T_341;
    wire [7:0] _WTEMP_191;
    PAD_UNSIGNED #(.width(1), .n(8)) u_pad_1902 (
        .y(_WTEMP_191),
        .in(1'h1)
    );
    ADD_UNSIGNED #(.width(8)) u_add_1903 (
        .y(_T_341),
        .a(_cntr__q),
        .b(_WTEMP_191)
    );
    wire [7:0] _T_342;
    TAIL #(.width(9), .n(1)) tail_1904 (
        .y(_T_342),
        .in(_T_341)
    );
    wire [7:0] _GEN_0;
    MUX_UNSIGNED #(.width(8)) u_mux_1905 (
        .y(_GEN_0),
        .sel(_T_336),
        .a(_T_342),
        .b(_cntr__q)
    );
    wire done;
    BITWISEAND #(.width(1)) bitwiseand_1906 (
        .y(done),
        .a(_T_336),
        .b(_T_339)
    );
    wire [31:0] iaddr;
    DIV_UNSIGNED #(.width_num(32), .width_den(3)) u_div_1907 (
        .y(iaddr),
        .num(_dut__io_icache_req_bits_addr),
        .den(3'h4)
    );
    wire [31:0] daddr;
    DIV_UNSIGNED #(.width_num(32), .width_den(3)) u_div_1908 (
        .y(daddr),
        .num(_dut__io_dcache_req_bits_addr),
        .den(3'h4)
    );
    wire _T_346;
    BITS #(.width(4), .high(0), .low(0)) bits_1909 (
        .y(_T_346),
        .in(_dut__io_dcache_req_bits_mask)
    );
    wire _T_347;
    BITWISEAND #(.width(1)) bitwiseand_1910 (
        .y(_T_347),
        .a(_dut__io_dcache_req_valid),
        .b(_T_346)
    );
    wire [19:0] _T_348;
    BITS #(.width(32), .high(19), .low(0)) bits_1911 (
        .y(_T_348),
        .in(daddr)
    );
    wire [31:0] _T_350;
    MUX_UNSIGNED #(.width(32)) u_mux_1912 (
        .y(_T_350),
        .sel(_T_347),
        .a(_dut__io_dcache_req_bits_data),
        .b(dmem__T_349_data)
    );
    wire [7:0] _T_351;
    BITS #(.width(32), .high(7), .low(0)) bits_1913 (
        .y(_T_351),
        .in(_T_350)
    );
    wire [8:0] _T_353;
    DSHL_UNSIGNED #(.width_in(8), .width_n(1)) u_dshl_1914 (
        .y(_T_353),
        .in(_T_351),
        .n(1'h0)
    );
    wire [31:0] _T_354;
    wire [31:0] _WTEMP_192;
    PAD_UNSIGNED #(.width(9), .n(32)) u_pad_1915 (
        .y(_WTEMP_192),
        .in(_T_353)
    );
    BITWISEOR #(.width(32)) bitwiseor_1916 (
        .y(_T_354),
        .a(32'h0),
        .b(_WTEMP_192)
    );
    wire _T_355;
    BITS #(.width(4), .high(1), .low(1)) bits_1917 (
        .y(_T_355),
        .in(_dut__io_dcache_req_bits_mask)
    );
    wire _T_356;
    BITWISEAND #(.width(1)) bitwiseand_1918 (
        .y(_T_356),
        .a(_dut__io_dcache_req_valid),
        .b(_T_355)
    );
    wire [19:0] _T_357;
    BITS #(.width(32), .high(19), .low(0)) bits_1919 (
        .y(_T_357),
        .in(daddr)
    );
    wire [31:0] _T_359;
    MUX_UNSIGNED #(.width(32)) u_mux_1920 (
        .y(_T_359),
        .sel(_T_356),
        .a(_dut__io_dcache_req_bits_data),
        .b(dmem__T_358_data)
    );
    wire [7:0] _T_360;
    BITS #(.width(32), .high(15), .low(8)) bits_1921 (
        .y(_T_360),
        .in(_T_359)
    );
    wire [22:0] _T_362;
    DSHL_UNSIGNED #(.width_in(8), .width_n(4)) u_dshl_1922 (
        .y(_T_362),
        .in(_T_360),
        .n(4'h8)
    );
    wire [31:0] _T_363;
    wire [31:0] _WTEMP_193;
    PAD_UNSIGNED #(.width(23), .n(32)) u_pad_1923 (
        .y(_WTEMP_193),
        .in(_T_362)
    );
    BITWISEOR #(.width(32)) bitwiseor_1924 (
        .y(_T_363),
        .a(_T_354),
        .b(_WTEMP_193)
    );
    wire _T_364;
    BITS #(.width(4), .high(2), .low(2)) bits_1925 (
        .y(_T_364),
        .in(_dut__io_dcache_req_bits_mask)
    );
    wire _T_365;
    BITWISEAND #(.width(1)) bitwiseand_1926 (
        .y(_T_365),
        .a(_dut__io_dcache_req_valid),
        .b(_T_364)
    );
    wire [19:0] _T_366;
    BITS #(.width(32), .high(19), .low(0)) bits_1927 (
        .y(_T_366),
        .in(daddr)
    );
    wire [31:0] _T_368;
    MUX_UNSIGNED #(.width(32)) u_mux_1928 (
        .y(_T_368),
        .sel(_T_365),
        .a(_dut__io_dcache_req_bits_data),
        .b(dmem__T_367_data)
    );
    wire [7:0] _T_369;
    BITS #(.width(32), .high(23), .low(16)) bits_1929 (
        .y(_T_369),
        .in(_T_368)
    );
    wire [38:0] _T_371;
    DSHL_UNSIGNED #(.width_in(8), .width_n(5)) u_dshl_1930 (
        .y(_T_371),
        .in(_T_369),
        .n(5'h10)
    );
    wire [38:0] _T_372;
    wire [38:0] _WTEMP_194;
    PAD_UNSIGNED #(.width(32), .n(39)) u_pad_1931 (
        .y(_WTEMP_194),
        .in(_T_363)
    );
    BITWISEOR #(.width(39)) bitwiseor_1932 (
        .y(_T_372),
        .a(_WTEMP_194),
        .b(_T_371)
    );
    wire _T_373;
    BITS #(.width(4), .high(3), .low(3)) bits_1933 (
        .y(_T_373),
        .in(_dut__io_dcache_req_bits_mask)
    );
    wire _T_374;
    BITWISEAND #(.width(1)) bitwiseand_1934 (
        .y(_T_374),
        .a(_dut__io_dcache_req_valid),
        .b(_T_373)
    );
    wire [19:0] _T_375;
    BITS #(.width(32), .high(19), .low(0)) bits_1935 (
        .y(_T_375),
        .in(daddr)
    );
    wire [31:0] _T_377;
    MUX_UNSIGNED #(.width(32)) u_mux_1936 (
        .y(_T_377),
        .sel(_T_374),
        .a(_dut__io_dcache_req_bits_data),
        .b(dmem__T_376_data)
    );
    wire [7:0] _T_378;
    BITS #(.width(32), .high(31), .low(24)) bits_1937 (
        .y(_T_378),
        .in(_T_377)
    );
    wire [38:0] _T_380;
    DSHL_UNSIGNED #(.width_in(8), .width_n(5)) u_dshl_1938 (
        .y(_T_380),
        .in(_T_378),
        .n(5'h18)
    );
    wire [38:0] write;
    BITWISEOR #(.width(39)) bitwiseor_1939 (
        .y(write),
        .a(_T_372),
        .b(_T_380)
    );
    wire _T_381;
    EQ_UNSIGNED #(.width(1)) u_eq_1940 (
        .y(_T_381),
        .a(_state__q),
        .b(1'h0)
    );
    wire _T_382;
    EQ_UNSIGNED #(.width(1)) u_eq_1941 (
        .y(_T_382),
        .a(_state__q),
        .b(1'h1)
    );
    wire _T_383;
    EQ_UNSIGNED #(.width(1)) u_eq_1942 (
        .y(_T_383),
        .a(_state__q),
        .b(1'h1)
    );
    wire [19:0] _T_384;
    BITS #(.width(32), .high(19), .low(0)) bits_1943 (
        .y(_T_384),
        .in(iaddr)
    );
    wire [19:0] _T_387;
    BITS #(.width(32), .high(19), .low(0)) bits_1944 (
        .y(_T_387),
        .in(daddr)
    );
    wire [7:0] _T_392;
    DSHR_UNSIGNED #(.width_in(8), .width_n(4)) u_dshr_1945 (
        .y(_T_392),
        .in(_cntr__q),
        .n(4'h8)
    );
    wire [7:0] _T_395;
    BITS #(.width(8), .high(7), .low(0)) bits_1946 (
        .y(_T_395),
        .in(_cntr__q)
    );
    wire [13:0] _T_397;
    MUL2_UNSIGNED #(.width_a(8), .width_b(6)) u_mul2_1947 (
        .y(_T_397),
        .a(_T_395),
        .b(6'h20)
    );
    wire [5119:0] _hex_0;
    assign _hex_0 = 5120'hFFDFF06F000000730040006F00100E130FF0000F10000073F10025733412907301428293000002973002B0731F8002931012907300028463DE0282930000029700000E130400006F00100E130FF0000F00055863F000257300051063F100257300000013000000130000001300000013000000130000001300000013FA1FF06FE25FF06F000F0463E30F0F1300000F17FBFF0CE334102FF3098F0F1300000F1700000013000000130000001300000013000000130000001300000013000000130000001300000013000000130000001300000013FFDFF06F780E1073539E6E130000001300000013000000130000001300000013000000130000001300000013000000130000001300000013000000130000001330500073FA0F5EE334202F73000000130000001300000013000000130540006FED9FF06F000F0463EE4F0F1300000F17020F1863EF0F0F1300000F1707FF0C6334102FF3158F0F1300000F17000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000200000000005000002600000026000000000000000000000000000000001000200050028000100200034000000000000045400000034000001000000000100F30002000000000000000000010101464C457F;
    wire [5119:0] _T_398;
    DSHR_UNSIGNED #(.width_in(5120), .width_n(14)) u_dshr_1948 (
        .y(_T_398),
        .in(_hex_0),
        .n(_T_397)
    );
    wire _T_400;
    EQ_UNSIGNED #(.width(1)) u_eq_1949 (
        .y(_T_400),
        .a(reset),
        .b(1'h0)
    );
    wire _T_401;
    EQ_UNSIGNED #(.width(1)) u_eq_1950 (
        .y(_T_401),
        .a(1'h0),
        .b(_state__q)
    );
    wire _GEN_1;
    MUX_UNSIGNED #(.width(1)) u_mux_1951 (
        .y(_GEN_1),
        .sel(done),
        .a(1'h1),
        .b(_state__q)
    );
    wire [7:0] _GEN_2;
    assign _GEN_2 = _cntr__q;
    wire _GEN_3;
    assign _GEN_3 = clock;
    wire _GEN_4;
    MUX_UNSIGNED #(.width(1)) u_mux_1952 (
        .y(_GEN_4),
        .sel(_T_401),
        .a(1'h1),
        .b(1'h0)
    );
    wire [31:0] chunk;
    BITS #(.width(5120), .high(31), .low(0)) bits_1953 (
        .y(chunk),
        .in(_T_398)
    );
    wire [31:0] _GEN_5;
    assign _GEN_5 = chunk;
    wire _GEN_6;
    MUX_UNSIGNED #(.width(1)) u_mux_1954 (
        .y(_GEN_6),
        .sel(_T_401),
        .a(_GEN_1),
        .b(_state__q)
    );
    wire _T_404;
    EQ_UNSIGNED #(.width(1)) u_eq_1955 (
        .y(_T_404),
        .a(1'h1),
        .b(_state__q)
    );
    wire _T_406;
    wire [3:0] _WTEMP_195;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1956 (
        .y(_WTEMP_195),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_1957 (
        .y(_T_406),
        .a(_dut__io_dcache_req_bits_mask),
        .b(_WTEMP_195)
    );
    wire [19:0] _T_407;
    BITS #(.width(32), .high(19), .low(0)) bits_1958 (
        .y(_T_407),
        .in(daddr)
    );
    wire [19:0] _GEN_7;
    assign _GEN_7 = _T_407;
    wire _GEN_8;
    assign _GEN_8 = clock;
    wire _GEN_9;
    MUX_UNSIGNED #(.width(1)) u_mux_1959 (
        .y(_GEN_9),
        .sel(_T_406),
        .a(1'h1),
        .b(1'h0)
    );
    wire [38:0] _GEN_10;
    assign _GEN_10 = write;
    wire _T_410;
    EQ_UNSIGNED #(.width(1)) u_eq_1960 (
        .y(_T_410),
        .a(_T_406),
        .b(1'h0)
    );
    wire [19:0] _GEN_11;
    assign _GEN_11 = _GEN_7;
    wire _GEN_12;
    assign _GEN_12 = _GEN_8;
    wire _GEN_13;
    MUX_UNSIGNED #(.width(1)) u_mux_1961 (
        .y(_GEN_13),
        .sel(_dut__io_dcache_req_valid),
        .a(_GEN_9),
        .b(1'h0)
    );
    wire [38:0] _GEN_14;
    assign _GEN_14 = _GEN_10;
    wire [32:0] _T_412;
    wire [31:0] _WTEMP_196;
    PAD_UNSIGNED #(.width(1), .n(32)) u_pad_1962 (
        .y(_WTEMP_196),
        .in(1'h1)
    );
    ADD_UNSIGNED #(.width(32)) u_add_1963 (
        .y(_T_412),
        .a(_cycle__q),
        .b(_WTEMP_196)
    );
    wire [31:0] _T_413;
    TAIL #(.width(33), .n(1)) tail_1964 (
        .y(_T_413),
        .in(_T_412)
    );
    wire _T_415;
    wire [31:0] _WTEMP_197;
    PAD_UNSIGNED #(.width(14), .n(32)) u_pad_1965 (
        .y(_WTEMP_197),
        .in(14'h3A98)
    );
    LT_UNSIGNED #(.width(32)) u_lt_1966 (
        .y(_T_415),
        .a(_cycle__q),
        .b(_WTEMP_197)
    );
    wire _T_416;
    BITWISEOR #(.width(1)) bitwiseor_1967 (
        .y(_T_416),
        .a(_T_415),
        .b(reset)
    );
    wire _T_418;
    EQ_UNSIGNED #(.width(1)) u_eq_1968 (
        .y(_T_418),
        .a(_T_416),
        .b(1'h0)
    );
    wire _T_420;
    wire [31:0] _WTEMP_198;
    PAD_UNSIGNED #(.width(1), .n(32)) u_pad_1969 (
        .y(_WTEMP_198),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(32)) u_neq_1970 (
        .y(_T_420),
        .a(_dut__io_host_tohost),
        .b(_WTEMP_198)
    );
    wire _T_422;
    EQ_UNSIGNED #(.width(1)) u_eq_1971 (
        .y(_T_422),
        .a(reset),
        .b(1'h0)
    );
    wire [31:0] _T_424;
    DSHR_UNSIGNED #(.width_in(32), .width_n(1)) u_dshr_1972 (
        .y(_T_424),
        .in(_dut__io_host_tohost),
        .n(1'h1)
    );
    wire _T_426;
    wire [31:0] _WTEMP_199;
    PAD_UNSIGNED #(.width(1), .n(32)) u_pad_1973 (
        .y(_WTEMP_199),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(32)) u_eq_1974 (
        .y(_T_426),
        .a(_T_424),
        .b(_WTEMP_199)
    );
    wire _T_427;
    BITWISEOR #(.width(1)) bitwiseor_1975 (
        .y(_T_427),
        .a(_T_426),
        .b(reset)
    );
    wire _T_429;
    EQ_UNSIGNED #(.width(1)) u_eq_1976 (
        .y(_T_429),
        .a(_T_427),
        .b(1'h0)
    );
    wire _T_431;
    EQ_UNSIGNED #(.width(1)) u_eq_1977 (
        .y(_T_431),
        .a(reset),
        .b(1'h0)
    );
    wire _T_433;
    EQ_UNSIGNED #(.width(1)) u_eq_1978 (
        .y(_T_433),
        .a(reset),
        .b(1'h0)
    );
    wire [19:0] _GEN_15;
    assign _GEN_15 = _GEN_11;
    wire _GEN_16;
    assign _GEN_16 = _GEN_12;
    wire _GEN_17;
    MUX_UNSIGNED #(.width(1)) u_mux_1979 (
        .y(_GEN_17),
        .sel(_T_404),
        .a(_GEN_13),
        .b(1'h0)
    );
    wire [38:0] _GEN_18;
    assign _GEN_18 = _GEN_14;
    wire [31:0] _GEN_19;
    MUX_UNSIGNED #(.width(32)) u_mux_1980 (
        .y(_GEN_19),
        .sel(_T_404),
        .a(_T_413),
        .b(_cycle__q)
    );
    assign __T_386__d = imem__T_385_data;
    assign __T_389__d = dmem__T_388_data;
    MUX_UNSIGNED #(.width(8)) u_mux_1981 (
        .y(_cntr__d),
        .sel(reset),
        .a(8'h0),
        .b(_GEN_0)
    );
    MUX_UNSIGNED #(.width(32)) u_mux_1982 (
        .y(_cycle__d),
        .sel(reset),
        .a(32'h0),
        .b(_GEN_19)
    );
    assign dmem__T_349_addr = _T_348;
    assign dmem__T_349_clk = clock;
    assign dmem__T_349_en = 1'h1;
    assign dmem__T_358_addr = _T_357;
    assign dmem__T_358_clk = clock;
    assign dmem__T_358_en = 1'h1;
    assign dmem__T_367_addr = _T_366;
    assign dmem__T_367_clk = clock;
    assign dmem__T_367_en = 1'h1;
    assign dmem__T_376_addr = _T_375;
    assign dmem__T_376_clk = clock;
    assign dmem__T_376_en = 1'h1;
    assign dmem__T_388_addr = _T_387;
    assign dmem__T_388_clk = clock;
    assign dmem__T_388_en = 1'h1;
    PAD_UNSIGNED #(.width(8), .n(20)) u_pad_1983 (
        .y(dmem__T_403_addr),
        .in(_GEN_2)
    );
    assign dmem__T_403_clk = _GEN_3;
    assign dmem__T_403_data = _GEN_5;
    assign dmem__T_403_en = _GEN_4;
    assign dmem__T_403_mask = _GEN_4;
    assign dmem__T_408_addr = _GEN_15;
    assign dmem__T_408_clk = _GEN_16;
    BITS #(.width(39), .high(31), .low(0)) bits_1984 (
        .y(dmem__T_408_data),
        .in(_GEN_18)
    );
    assign dmem__T_408_en = _GEN_17;
    assign dmem__T_408_mask = _GEN_17;
    assign _dut__clock = clock;
    assign _dut__io_dcache_resp_bits_data = __T_389__q;
    assign _dut__io_dcache_resp_valid = _T_383;
    PAD_UNSIGNED #(.width(1), .n(32)) u_pad_1985 (
        .y(_dut__io_host_fromhost_bits),
        .in(1'h0)
    );
    assign _dut__io_host_fromhost_valid = 1'h0;
    assign _dut__io_icache_resp_bits_data = __T_386__q;
    assign _dut__io_icache_resp_valid = _T_382;
    assign _dut__reset = _T_381;
    assign imem__T_385_addr = _T_384;
    assign imem__T_385_clk = clock;
    assign imem__T_385_en = 1'h1;
    PAD_UNSIGNED #(.width(8), .n(20)) u_pad_1986 (
        .y(imem__T_402_addr),
        .in(_GEN_2)
    );
    assign imem__T_402_clk = _GEN_3;
    assign imem__T_402_data = _GEN_5;
    assign imem__T_402_en = _GEN_4;
    assign imem__T_402_mask = _GEN_4;
    MUX_UNSIGNED #(.width(1)) u_mux_1987 (
        .y(_state__d),
        .sel(reset),
        .a(1'h0),
        .b(_GEN_6)
    );
endmodule //CoreTester
module Core(
    input clock,
    input reset,
    input io_host_fromhost_valid,
    input [31:0] io_host_fromhost_bits,
    output [31:0] io_host_tohost,
    output io_icache_abort,
    output io_icache_req_valid,
    output [31:0] io_icache_req_bits_addr,
    output [31:0] io_icache_req_bits_data,
    output [3:0] io_icache_req_bits_mask,
    input io_icache_resp_valid,
    input [31:0] io_icache_resp_bits_data,
    output io_dcache_abort,
    output io_dcache_req_valid,
    output [31:0] io_dcache_req_bits_addr,
    output [31:0] io_dcache_req_bits_data,
    output [3:0] io_dcache_req_bits_mask,
    input io_dcache_resp_valid,
    input [31:0] io_dcache_resp_bits_data
);
    wire _dpath__clock;
    wire _dpath__reset;
    wire _dpath__io_host_fromhost_valid;
    wire [31:0] _dpath__io_host_fromhost_bits;
    wire [31:0] _dpath__io_host_tohost;
    wire _dpath__io_icache_abort;
    wire _dpath__io_icache_req_valid;
    wire [31:0] _dpath__io_icache_req_bits_addr;
    wire [31:0] _dpath__io_icache_req_bits_data;
    wire [3:0] _dpath__io_icache_req_bits_mask;
    wire _dpath__io_icache_resp_valid;
    wire [31:0] _dpath__io_icache_resp_bits_data;
    wire _dpath__io_dcache_abort;
    wire _dpath__io_dcache_req_valid;
    wire [31:0] _dpath__io_dcache_req_bits_addr;
    wire [31:0] _dpath__io_dcache_req_bits_data;
    wire [3:0] _dpath__io_dcache_req_bits_mask;
    wire _dpath__io_dcache_resp_valid;
    wire [31:0] _dpath__io_dcache_resp_bits_data;
    wire [31:0] _dpath__io_ctrl_inst;
    wire [1:0] _dpath__io_ctrl_pc_sel;
    wire _dpath__io_ctrl_inst_kill;
    wire _dpath__io_ctrl_A_sel;
    wire _dpath__io_ctrl_B_sel;
    wire [2:0] _dpath__io_ctrl_imm_sel;
    wire [3:0] _dpath__io_ctrl_alu_op;
    wire [2:0] _dpath__io_ctrl_br_type;
    wire [1:0] _dpath__io_ctrl_st_type;
    wire [2:0] _dpath__io_ctrl_ld_type;
    wire [1:0] _dpath__io_ctrl_wb_sel;
    wire _dpath__io_ctrl_wb_en;
    wire [2:0] _dpath__io_ctrl_csr_cmd;
    wire _dpath__io_ctrl_illegal;
    Datapath dpath (
        .clock(_dpath__clock),
        .reset(_dpath__reset),
        .io_host_fromhost_valid(_dpath__io_host_fromhost_valid),
        .io_host_fromhost_bits(_dpath__io_host_fromhost_bits),
        .io_host_tohost(_dpath__io_host_tohost),
        .io_icache_abort(_dpath__io_icache_abort),
        .io_icache_req_valid(_dpath__io_icache_req_valid),
        .io_icache_req_bits_addr(_dpath__io_icache_req_bits_addr),
        .io_icache_req_bits_data(_dpath__io_icache_req_bits_data),
        .io_icache_req_bits_mask(_dpath__io_icache_req_bits_mask),
        .io_icache_resp_valid(_dpath__io_icache_resp_valid),
        .io_icache_resp_bits_data(_dpath__io_icache_resp_bits_data),
        .io_dcache_abort(_dpath__io_dcache_abort),
        .io_dcache_req_valid(_dpath__io_dcache_req_valid),
        .io_dcache_req_bits_addr(_dpath__io_dcache_req_bits_addr),
        .io_dcache_req_bits_data(_dpath__io_dcache_req_bits_data),
        .io_dcache_req_bits_mask(_dpath__io_dcache_req_bits_mask),
        .io_dcache_resp_valid(_dpath__io_dcache_resp_valid),
        .io_dcache_resp_bits_data(_dpath__io_dcache_resp_bits_data),
        .io_ctrl_inst(_dpath__io_ctrl_inst),
        .io_ctrl_pc_sel(_dpath__io_ctrl_pc_sel),
        .io_ctrl_inst_kill(_dpath__io_ctrl_inst_kill),
        .io_ctrl_A_sel(_dpath__io_ctrl_A_sel),
        .io_ctrl_B_sel(_dpath__io_ctrl_B_sel),
        .io_ctrl_imm_sel(_dpath__io_ctrl_imm_sel),
        .io_ctrl_alu_op(_dpath__io_ctrl_alu_op),
        .io_ctrl_br_type(_dpath__io_ctrl_br_type),
        .io_ctrl_st_type(_dpath__io_ctrl_st_type),
        .io_ctrl_ld_type(_dpath__io_ctrl_ld_type),
        .io_ctrl_wb_sel(_dpath__io_ctrl_wb_sel),
        .io_ctrl_wb_en(_dpath__io_ctrl_wb_en),
        .io_ctrl_csr_cmd(_dpath__io_ctrl_csr_cmd),
        .io_ctrl_illegal(_dpath__io_ctrl_illegal)
    );
    wire _ctrl__clock;
    wire _ctrl__reset;
    wire [31:0] _ctrl__io_inst;
    wire [1:0] _ctrl__io_pc_sel;
    wire _ctrl__io_inst_kill;
    wire _ctrl__io_A_sel;
    wire _ctrl__io_B_sel;
    wire [2:0] _ctrl__io_imm_sel;
    wire [3:0] _ctrl__io_alu_op;
    wire [2:0] _ctrl__io_br_type;
    wire [1:0] _ctrl__io_st_type;
    wire [2:0] _ctrl__io_ld_type;
    wire [1:0] _ctrl__io_wb_sel;
    wire _ctrl__io_wb_en;
    wire [2:0] _ctrl__io_csr_cmd;
    wire _ctrl__io_illegal;
    Control ctrl (
        .clock(_ctrl__clock),
        .reset(_ctrl__reset),
        .io_inst(_ctrl__io_inst),
        .io_pc_sel(_ctrl__io_pc_sel),
        .io_inst_kill(_ctrl__io_inst_kill),
        .io_A_sel(_ctrl__io_A_sel),
        .io_B_sel(_ctrl__io_B_sel),
        .io_imm_sel(_ctrl__io_imm_sel),
        .io_alu_op(_ctrl__io_alu_op),
        .io_br_type(_ctrl__io_br_type),
        .io_st_type(_ctrl__io_st_type),
        .io_ld_type(_ctrl__io_ld_type),
        .io_wb_sel(_ctrl__io_wb_sel),
        .io_wb_en(_ctrl__io_wb_en),
        .io_csr_cmd(_ctrl__io_csr_cmd),
        .io_illegal(_ctrl__io_illegal)
    );
    assign _ctrl__clock = clock;
    assign _ctrl__io_inst = _dpath__io_ctrl_inst;
    assign _ctrl__reset = reset;
    assign _dpath__clock = clock;
    assign _dpath__io_ctrl_A_sel = _ctrl__io_A_sel;
    assign _dpath__io_ctrl_B_sel = _ctrl__io_B_sel;
    assign _dpath__io_ctrl_alu_op = _ctrl__io_alu_op;
    assign _dpath__io_ctrl_br_type = _ctrl__io_br_type;
    assign _dpath__io_ctrl_csr_cmd = _ctrl__io_csr_cmd;
    assign _dpath__io_ctrl_illegal = _ctrl__io_illegal;
    assign _dpath__io_ctrl_imm_sel = _ctrl__io_imm_sel;
    assign _dpath__io_ctrl_inst_kill = _ctrl__io_inst_kill;
    assign _dpath__io_ctrl_ld_type = _ctrl__io_ld_type;
    assign _dpath__io_ctrl_pc_sel = _ctrl__io_pc_sel;
    assign _dpath__io_ctrl_st_type = _ctrl__io_st_type;
    assign _dpath__io_ctrl_wb_en = _ctrl__io_wb_en;
    assign _dpath__io_ctrl_wb_sel = _ctrl__io_wb_sel;
    assign _dpath__io_dcache_resp_bits_data = io_dcache_resp_bits_data;
    assign _dpath__io_dcache_resp_valid = io_dcache_resp_valid;
    assign _dpath__io_host_fromhost_bits = io_host_fromhost_bits;
    assign _dpath__io_host_fromhost_valid = io_host_fromhost_valid;
    assign _dpath__io_icache_resp_bits_data = io_icache_resp_bits_data;
    assign _dpath__io_icache_resp_valid = io_icache_resp_valid;
    assign _dpath__reset = reset;
    assign io_dcache_abort = _dpath__io_dcache_abort;
    assign io_dcache_req_bits_addr = _dpath__io_dcache_req_bits_addr;
    assign io_dcache_req_bits_data = _dpath__io_dcache_req_bits_data;
    assign io_dcache_req_bits_mask = _dpath__io_dcache_req_bits_mask;
    assign io_dcache_req_valid = _dpath__io_dcache_req_valid;
    assign io_host_tohost = _dpath__io_host_tohost;
    assign io_icache_abort = _dpath__io_icache_abort;
    assign io_icache_req_bits_addr = _dpath__io_icache_req_bits_addr;
    assign io_icache_req_bits_data = _dpath__io_icache_req_bits_data;
    assign io_icache_req_bits_mask = _dpath__io_icache_req_bits_mask;
    assign io_icache_req_valid = _dpath__io_icache_req_valid;
endmodule //Core
module Datapath(
    input clock,
    input reset,
    input io_host_fromhost_valid,
    input [31:0] io_host_fromhost_bits,
    output [31:0] io_host_tohost,
    output io_icache_abort,
    output io_icache_req_valid,
    output [31:0] io_icache_req_bits_addr,
    output [31:0] io_icache_req_bits_data,
    output [3:0] io_icache_req_bits_mask,
    input io_icache_resp_valid,
    input [31:0] io_icache_resp_bits_data,
    output io_dcache_abort,
    output io_dcache_req_valid,
    output [31:0] io_dcache_req_bits_addr,
    output [31:0] io_dcache_req_bits_data,
    output [3:0] io_dcache_req_bits_mask,
    input io_dcache_resp_valid,
    input [31:0] io_dcache_resp_bits_data,
    output [31:0] io_ctrl_inst,
    input [1:0] io_ctrl_pc_sel,
    input io_ctrl_inst_kill,
    input io_ctrl_A_sel,
    input io_ctrl_B_sel,
    input [2:0] io_ctrl_imm_sel,
    input [3:0] io_ctrl_alu_op,
    input [2:0] io_ctrl_br_type,
    input [1:0] io_ctrl_st_type,
    input [2:0] io_ctrl_ld_type,
    input [1:0] io_ctrl_wb_sel,
    input io_ctrl_wb_en,
    input [2:0] io_ctrl_csr_cmd,
    input io_ctrl_illegal
);
    wire _csr__clock;
    wire _csr__reset;
    wire _csr__io_stall;
    wire [2:0] _csr__io_cmd;
    wire [31:0] _csr__io_in;
    wire [31:0] _csr__io_out;
    wire [31:0] _csr__io_pc;
    wire [31:0] _csr__io_addr;
    wire [31:0] _csr__io_inst;
    wire _csr__io_illegal;
    wire [1:0] _csr__io_st_type;
    wire [2:0] _csr__io_ld_type;
    wire _csr__io_pc_check;
    wire _csr__io_expt;
    wire [31:0] _csr__io_evec;
    wire [31:0] _csr__io_epc;
    wire _csr__io_host_fromhost_valid;
    wire [31:0] _csr__io_host_fromhost_bits;
    wire [31:0] _csr__io_host_tohost;
    CSR csr (
        .clock(_csr__clock),
        .reset(_csr__reset),
        .io_stall(_csr__io_stall),
        .io_cmd(_csr__io_cmd),
        .io_in(_csr__io_in),
        .io_out(_csr__io_out),
        .io_pc(_csr__io_pc),
        .io_addr(_csr__io_addr),
        .io_inst(_csr__io_inst),
        .io_illegal(_csr__io_illegal),
        .io_st_type(_csr__io_st_type),
        .io_ld_type(_csr__io_ld_type),
        .io_pc_check(_csr__io_pc_check),
        .io_expt(_csr__io_expt),
        .io_evec(_csr__io_evec),
        .io_epc(_csr__io_epc),
        .io_host_fromhost_valid(_csr__io_host_fromhost_valid),
        .io_host_fromhost_bits(_csr__io_host_fromhost_bits),
        .io_host_tohost(_csr__io_host_tohost)
    );
    wire _regFile__clock;
    wire _regFile__reset;
    wire [4:0] _regFile__io_raddr1;
    wire [4:0] _regFile__io_raddr2;
    wire [31:0] _regFile__io_rdata1;
    wire [31:0] _regFile__io_rdata2;
    wire _regFile__io_wen;
    wire [4:0] _regFile__io_waddr;
    wire [31:0] _regFile__io_wdata;
    RegFile regFile (
        .clock(_regFile__clock),
        .reset(_regFile__reset),
        .io_raddr1(_regFile__io_raddr1),
        .io_raddr2(_regFile__io_raddr2),
        .io_rdata1(_regFile__io_rdata1),
        .io_rdata2(_regFile__io_rdata2),
        .io_wen(_regFile__io_wen),
        .io_waddr(_regFile__io_waddr),
        .io_wdata(_regFile__io_wdata)
    );
    wire _alu__clock;
    wire _alu__reset;
    wire [31:0] _alu__io_A;
    wire [31:0] _alu__io_B;
    wire [3:0] _alu__io_alu_op;
    wire [31:0] _alu__io_out;
    wire [31:0] _alu__io_sum;
    ALUArea alu (
        .clock(_alu__clock),
        .reset(_alu__reset),
        .io_A(_alu__io_A),
        .io_B(_alu__io_B),
        .io_alu_op(_alu__io_alu_op),
        .io_out(_alu__io_out),
        .io_sum(_alu__io_sum)
    );
    wire _immGen__clock;
    wire _immGen__reset;
    wire [31:0] _immGen__io_inst;
    wire [2:0] _immGen__io_sel;
    wire [31:0] _immGen__io_out;
    ImmGenWire immGen (
        .clock(_immGen__clock),
        .reset(_immGen__reset),
        .io_inst(_immGen__io_inst),
        .io_sel(_immGen__io_sel),
        .io_out(_immGen__io_out)
    );
    wire _brCond__clock;
    wire _brCond__reset;
    wire [31:0] _brCond__io_rs1;
    wire [31:0] _brCond__io_rs2;
    wire [2:0] _brCond__io_br_type;
    wire _brCond__io_taken;
    BrCondArea brCond (
        .clock(_brCond__clock),
        .reset(_brCond__reset),
        .io_rs1(_brCond__io_rs1),
        .io_rs2(_brCond__io_rs2),
        .io_br_type(_brCond__io_br_type),
        .io_taken(_brCond__io_taken)
    );
    wire [31:0] _fe_inst__q;
    wire [31:0] _fe_inst__d;
    DFF_POSCLK #(.width(32)) fe_inst (
        .q(_fe_inst__q),
        .d(_fe_inst__d),
        .clk(clock)
    );
    wire [32:0] _fe_pc__q;
    wire [32:0] _fe_pc__d;
    DFF_POSCLK #(.width(33)) fe_pc (
        .q(_fe_pc__q),
        .d(_fe_pc__d),
        .clk(clock)
    );
    wire [31:0] _ew_inst__q;
    wire [31:0] _ew_inst__d;
    DFF_POSCLK #(.width(32)) ew_inst (
        .q(_ew_inst__q),
        .d(_ew_inst__d),
        .clk(clock)
    );
    wire [32:0] _ew_pc__q;
    wire [32:0] _ew_pc__d;
    DFF_POSCLK #(.width(33)) ew_pc (
        .q(_ew_pc__q),
        .d(_ew_pc__d),
        .clk(clock)
    );
    wire [31:0] _ew_alu__q;
    wire [31:0] _ew_alu__d;
    DFF_POSCLK #(.width(32)) ew_alu (
        .q(_ew_alu__q),
        .d(_ew_alu__d),
        .clk(clock)
    );
    wire [31:0] _csr_in__q;
    wire [31:0] _csr_in__d;
    DFF_POSCLK #(.width(32)) csr_in (
        .q(_csr_in__q),
        .d(_csr_in__d),
        .clk(clock)
    );
    wire [1:0] _st_type__q;
    wire [1:0] _st_type__d;
    DFF_POSCLK #(.width(2)) st_type (
        .q(_st_type__q),
        .d(_st_type__d),
        .clk(clock)
    );
    wire [2:0] _ld_type__q;
    wire [2:0] _ld_type__d;
    DFF_POSCLK #(.width(3)) ld_type (
        .q(_ld_type__q),
        .d(_ld_type__d),
        .clk(clock)
    );
    wire [1:0] _wb_sel__q;
    wire [1:0] _wb_sel__d;
    DFF_POSCLK #(.width(2)) wb_sel (
        .q(_wb_sel__q),
        .d(_wb_sel__d),
        .clk(clock)
    );
    wire _wb_en__q;
    wire _wb_en__d;
    DFF_POSCLK #(.width(1)) wb_en (
        .q(_wb_en__q),
        .d(_wb_en__d),
        .clk(clock)
    );
    wire [2:0] _csr_cmd__q;
    wire [2:0] _csr_cmd__d;
    DFF_POSCLK #(.width(3)) csr_cmd (
        .q(_csr_cmd__q),
        .d(_csr_cmd__d),
        .clk(clock)
    );
    wire _illegal__q;
    wire _illegal__d;
    DFF_POSCLK #(.width(1)) illegal (
        .q(_illegal__q),
        .d(_illegal__d),
        .clk(clock)
    );
    wire _pc_check__q;
    wire _pc_check__d;
    DFF_POSCLK #(.width(1)) pc_check (
        .q(_pc_check__q),
        .d(_pc_check__d),
        .clk(clock)
    );
    wire _started__q;
    wire _started__d;
    DFF_POSCLK #(.width(1)) started (
        .q(_started__q),
        .d(_started__d),
        .clk(clock)
    );
    wire [32:0] _pc__q;
    wire [32:0] _pc__d;
    DFF_POSCLK #(.width(33)) pc (
        .q(_pc__q),
        .d(_pc__d),
        .clk(clock)
    );
    wire _T_240;
    EQ_UNSIGNED #(.width(1)) u_eq_1030 (
        .y(_T_240),
        .a(io_icache_resp_valid),
        .b(1'h0)
    );
    wire _T_242;
    EQ_UNSIGNED #(.width(1)) u_eq_1031 (
        .y(_T_242),
        .a(io_dcache_resp_valid),
        .b(1'h0)
    );
    wire stall;
    BITWISEOR #(.width(1)) bitwiseor_1032 (
        .y(stall),
        .a(_T_240),
        .b(_T_242)
    );
    wire [32:0] _T_245;
    assign _T_245 = 33'h1FC;
    wire [31:0] _T_246;
    assign _T_246 = 32'h1FC;
    wire _T_247;
    EQ_UNSIGNED #(.width(2)) u_eq_1033 (
        .y(_T_247),
        .a(io_ctrl_pc_sel),
        .b(2'h3)
    );
    wire _T_248;
    EQ_UNSIGNED #(.width(2)) u_eq_1034 (
        .y(_T_248),
        .a(io_ctrl_pc_sel),
        .b(2'h1)
    );
    wire _T_249;
    BITWISEOR #(.width(1)) bitwiseor_1035 (
        .y(_T_249),
        .a(_T_248),
        .b(_brCond__io_taken)
    );
    wire [31:0] _T_251;
    DSHR_UNSIGNED #(.width_in(32), .width_n(1)) u_dshr_1036 (
        .y(_T_251),
        .in(_alu__io_sum),
        .n(1'h1)
    );
    wire [32:0] _T_253;
    DSHL_UNSIGNED #(.width_in(32), .width_n(1)) u_dshl_1037 (
        .y(_T_253),
        .in(_T_251),
        .n(1'h1)
    );
    wire _T_254;
    EQ_UNSIGNED #(.width(2)) u_eq_1038 (
        .y(_T_254),
        .a(io_ctrl_pc_sel),
        .b(2'h2)
    );
    wire [33:0] _T_256;
    wire [32:0] _WTEMP_79;
    PAD_UNSIGNED #(.width(3), .n(33)) u_pad_1039 (
        .y(_WTEMP_79),
        .in(3'h4)
    );
    ADD_UNSIGNED #(.width(33)) u_add_1040 (
        .y(_T_256),
        .a(_pc__q),
        .b(_WTEMP_79)
    );
    wire [32:0] _T_257;
    TAIL #(.width(34), .n(1)) tail_1041 (
        .y(_T_257),
        .in(_T_256)
    );
    wire [32:0] _T_258;
    MUX_UNSIGNED #(.width(33)) u_mux_1042 (
        .y(_T_258),
        .sel(_T_254),
        .a(_pc__q),
        .b(_T_257)
    );
    wire [32:0] _T_259;
    MUX_UNSIGNED #(.width(33)) u_mux_1043 (
        .y(_T_259),
        .sel(_T_249),
        .a(_T_253),
        .b(_T_258)
    );
    wire [32:0] _T_260;
    wire [32:0] _WTEMP_80;
    PAD_UNSIGNED #(.width(32), .n(33)) u_pad_1044 (
        .y(_WTEMP_80),
        .in(_csr__io_epc)
    );
    MUX_UNSIGNED #(.width(33)) u_mux_1045 (
        .y(_T_260),
        .sel(_T_247),
        .a(_WTEMP_80),
        .b(_T_259)
    );
    wire [32:0] _T_261;
    wire [32:0] _WTEMP_81;
    PAD_UNSIGNED #(.width(32), .n(33)) u_pad_1046 (
        .y(_WTEMP_81),
        .in(_csr__io_evec)
    );
    MUX_UNSIGNED #(.width(33)) u_mux_1047 (
        .y(_T_261),
        .sel(_csr__io_expt),
        .a(_WTEMP_81),
        .b(_T_260)
    );
    wire [32:0] npc;
    MUX_UNSIGNED #(.width(33)) u_mux_1048 (
        .y(npc),
        .sel(stall),
        .a(_pc__q),
        .b(_T_261)
    );
    wire _T_262;
    BITWISEOR #(.width(1)) bitwiseor_1049 (
        .y(_T_262),
        .a(_started__q),
        .b(io_ctrl_inst_kill)
    );
    wire _T_263;
    BITWISEOR #(.width(1)) bitwiseor_1050 (
        .y(_T_263),
        .a(_T_262),
        .b(_brCond__io_taken)
    );
    wire _T_264;
    BITWISEOR #(.width(1)) bitwiseor_1051 (
        .y(_T_264),
        .a(_T_263),
        .b(_csr__io_expt)
    );
    wire [31:0] inst;
    MUX_UNSIGNED #(.width(32)) u_mux_1052 (
        .y(inst),
        .sel(_T_264),
        .a(32'h13),
        .b(io_icache_resp_bits_data)
    );
    wire _T_269;
    EQ_UNSIGNED #(.width(1)) u_eq_1053 (
        .y(_T_269),
        .a(stall),
        .b(1'h0)
    );
    wire _T_272;
    EQ_UNSIGNED #(.width(1)) u_eq_1054 (
        .y(_T_272),
        .a(stall),
        .b(1'h0)
    );
    wire [32:0] _GEN_0;
    MUX_UNSIGNED #(.width(33)) u_mux_1055 (
        .y(_GEN_0),
        .sel(_T_272),
        .a(_pc__q),
        .b(_fe_pc__q)
    );
    wire [31:0] _GEN_1;
    MUX_UNSIGNED #(.width(32)) u_mux_1056 (
        .y(_GEN_1),
        .sel(_T_272),
        .a(inst),
        .b(_fe_inst__q)
    );
    wire [4:0] rd_addr;
    BITS #(.width(32), .high(11), .low(7)) bits_1057 (
        .y(rd_addr),
        .in(_fe_inst__q)
    );
    wire [4:0] rs1_addr;
    BITS #(.width(32), .high(19), .low(15)) bits_1058 (
        .y(rs1_addr),
        .in(_fe_inst__q)
    );
    wire [4:0] rs2_addr;
    BITS #(.width(32), .high(24), .low(20)) bits_1059 (
        .y(rs2_addr),
        .in(_fe_inst__q)
    );
    wire [4:0] wb_rd_addr;
    BITS #(.width(32), .high(11), .low(7)) bits_1060 (
        .y(wb_rd_addr),
        .in(_ew_inst__q)
    );
    wire _T_274;
    wire [4:0] _WTEMP_82;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_1061 (
        .y(_WTEMP_82),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(5)) u_neq_1062 (
        .y(_T_274),
        .a(rs1_addr),
        .b(_WTEMP_82)
    );
    wire _T_275;
    BITWISEAND #(.width(1)) bitwiseand_1063 (
        .y(_T_275),
        .a(_wb_en__q),
        .b(_T_274)
    );
    wire _T_276;
    EQ_UNSIGNED #(.width(5)) u_eq_1064 (
        .y(_T_276),
        .a(rs1_addr),
        .b(wb_rd_addr)
    );
    wire rs1hazard;
    BITWISEAND #(.width(1)) bitwiseand_1065 (
        .y(rs1hazard),
        .a(_T_275),
        .b(_T_276)
    );
    wire _T_278;
    wire [4:0] _WTEMP_83;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_1066 (
        .y(_WTEMP_83),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(5)) u_neq_1067 (
        .y(_T_278),
        .a(rs2_addr),
        .b(_WTEMP_83)
    );
    wire _T_279;
    BITWISEAND #(.width(1)) bitwiseand_1068 (
        .y(_T_279),
        .a(_wb_en__q),
        .b(_T_278)
    );
    wire _T_280;
    EQ_UNSIGNED #(.width(5)) u_eq_1069 (
        .y(_T_280),
        .a(rs2_addr),
        .b(wb_rd_addr)
    );
    wire rs2hazard;
    BITWISEAND #(.width(1)) bitwiseand_1070 (
        .y(rs2hazard),
        .a(_T_279),
        .b(_T_280)
    );
    wire _T_281;
    EQ_UNSIGNED #(.width(2)) u_eq_1071 (
        .y(_T_281),
        .a(_wb_sel__q),
        .b(2'h0)
    );
    wire _T_282;
    BITWISEAND #(.width(1)) bitwiseand_1072 (
        .y(_T_282),
        .a(_T_281),
        .b(rs1hazard)
    );
    wire [31:0] rs1;
    MUX_UNSIGNED #(.width(32)) u_mux_1073 (
        .y(rs1),
        .sel(_T_282),
        .a(_ew_alu__q),
        .b(_regFile__io_rdata1)
    );
    wire _T_283;
    EQ_UNSIGNED #(.width(2)) u_eq_1074 (
        .y(_T_283),
        .a(_wb_sel__q),
        .b(2'h0)
    );
    wire _T_284;
    BITWISEAND #(.width(1)) bitwiseand_1075 (
        .y(_T_284),
        .a(_T_283),
        .b(rs2hazard)
    );
    wire [31:0] rs2;
    MUX_UNSIGNED #(.width(32)) u_mux_1076 (
        .y(rs2),
        .sel(_T_284),
        .a(_ew_alu__q),
        .b(_regFile__io_rdata2)
    );
    wire _T_285;
    EQ_UNSIGNED #(.width(1)) u_eq_1077 (
        .y(_T_285),
        .a(io_ctrl_A_sel),
        .b(1'h1)
    );
    wire [32:0] _T_286;
    wire [32:0] _WTEMP_84;
    PAD_UNSIGNED #(.width(32), .n(33)) u_pad_1078 (
        .y(_WTEMP_84),
        .in(rs1)
    );
    MUX_UNSIGNED #(.width(33)) u_mux_1079 (
        .y(_T_286),
        .sel(_T_285),
        .a(_WTEMP_84),
        .b(_fe_pc__q)
    );
    wire _T_287;
    EQ_UNSIGNED #(.width(1)) u_eq_1080 (
        .y(_T_287),
        .a(io_ctrl_B_sel),
        .b(1'h1)
    );
    wire [31:0] _T_288;
    MUX_UNSIGNED #(.width(32)) u_mux_1081 (
        .y(_T_288),
        .sel(_T_287),
        .a(rs2),
        .b(_immGen__io_out)
    );
    wire [31:0] _T_289;
    MUX_UNSIGNED #(.width(32)) u_mux_1082 (
        .y(_T_289),
        .sel(stall),
        .a(_ew_alu__q),
        .b(_alu__io_sum)
    );
    wire [31:0] _T_291;
    DSHR_UNSIGNED #(.width_in(32), .width_n(2)) u_dshr_1083 (
        .y(_T_291),
        .in(_T_289),
        .n(2'h2)
    );
    wire [34:0] daddr;
    DSHL_UNSIGNED #(.width_in(32), .width_n(2)) u_dshl_1084 (
        .y(daddr),
        .in(_T_291),
        .n(2'h2)
    );
    wire _T_293;
    BITS #(.width(32), .high(1), .low(1)) bits_1085 (
        .y(_T_293),
        .in(_alu__io_sum)
    );
    wire [7:0] _T_295;
    DSHL_UNSIGNED #(.width_in(1), .width_n(3)) u_dshl_1086 (
        .y(_T_295),
        .in(_T_293),
        .n(3'h4)
    );
    wire _T_296;
    BITS #(.width(32), .high(0), .low(0)) bits_1087 (
        .y(_T_296),
        .in(_alu__io_sum)
    );
    wire [3:0] _T_298;
    DSHL_UNSIGNED #(.width_in(1), .width_n(2)) u_dshl_1088 (
        .y(_T_298),
        .in(_T_296),
        .n(2'h3)
    );
    wire [7:0] woffset;
    wire [7:0] _WTEMP_85;
    PAD_UNSIGNED #(.width(4), .n(8)) u_pad_1089 (
        .y(_WTEMP_85),
        .in(_T_298)
    );
    BITWISEOR #(.width(8)) bitwiseor_1090 (
        .y(woffset),
        .a(_T_295),
        .b(_WTEMP_85)
    );
    wire _T_300;
    EQ_UNSIGNED #(.width(1)) u_eq_1091 (
        .y(_T_300),
        .a(stall),
        .b(1'h0)
    );
    wire _T_302;
    wire [1:0] _WTEMP_86;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_1092 (
        .y(_WTEMP_86),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(2)) u_neq_1093 (
        .y(_T_302),
        .a(io_ctrl_st_type),
        .b(_WTEMP_86)
    );
    wire _T_304;
    wire [2:0] _WTEMP_87;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_1094 (
        .y(_WTEMP_87),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(3)) u_neq_1095 (
        .y(_T_304),
        .a(io_ctrl_ld_type),
        .b(_WTEMP_87)
    );
    wire _T_305;
    BITWISEOR #(.width(1)) bitwiseor_1096 (
        .y(_T_305),
        .a(_T_302),
        .b(_T_304)
    );
    wire _T_306;
    BITWISEAND #(.width(1)) bitwiseand_1097 (
        .y(_T_306),
        .a(_T_300),
        .b(_T_305)
    );
    wire [286:0] _T_307;
    DSHL_UNSIGNED #(.width_in(32), .width_n(8)) u_dshl_1098 (
        .y(_T_307),
        .in(rs2),
        .n(woffset)
    );
    wire [1:0] _T_308;
    MUX_UNSIGNED #(.width(2)) u_mux_1099 (
        .y(_T_308),
        .sel(stall),
        .a(_st_type__q),
        .b(io_ctrl_st_type)
    );
    wire [1:0] _T_312;
    BITS #(.width(32), .high(1), .low(0)) bits_1100 (
        .y(_T_312),
        .in(_alu__io_sum)
    );
    wire [4:0] _T_313;
    DSHL_UNSIGNED #(.width_in(2), .width_n(2)) u_dshl_1101 (
        .y(_T_313),
        .in(2'h3),
        .n(_T_312)
    );
    wire [1:0] _T_315;
    BITS #(.width(32), .high(1), .low(0)) bits_1102 (
        .y(_T_315),
        .in(_alu__io_sum)
    );
    wire [3:0] _T_316;
    DSHL_UNSIGNED #(.width_in(1), .width_n(2)) u_dshl_1103 (
        .y(_T_316),
        .in(1'h1),
        .n(_T_315)
    );
    wire _T_317;
    EQ_UNSIGNED #(.width(2)) u_eq_1104 (
        .y(_T_317),
        .a(2'h3),
        .b(_T_308)
    );
    wire [3:0] _T_318;
    wire [3:0] _WTEMP_88;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1105 (
        .y(_WTEMP_88),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(4)) u_mux_1106 (
        .y(_T_318),
        .sel(_T_317),
        .a(_T_316),
        .b(_WTEMP_88)
    );
    wire _T_319;
    EQ_UNSIGNED #(.width(2)) u_eq_1107 (
        .y(_T_319),
        .a(2'h2),
        .b(_T_308)
    );
    wire [4:0] _T_320;
    wire [4:0] _WTEMP_89;
    PAD_UNSIGNED #(.width(4), .n(5)) u_pad_1108 (
        .y(_WTEMP_89),
        .in(_T_318)
    );
    MUX_UNSIGNED #(.width(5)) u_mux_1109 (
        .y(_T_320),
        .sel(_T_319),
        .a(_T_313),
        .b(_WTEMP_89)
    );
    wire _T_321;
    EQ_UNSIGNED #(.width(2)) u_eq_1110 (
        .y(_T_321),
        .a(2'h1),
        .b(_T_308)
    );
    wire [4:0] _T_322;
    wire [4:0] _WTEMP_90;
    PAD_UNSIGNED #(.width(4), .n(5)) u_pad_1111 (
        .y(_WTEMP_90),
        .in(4'hF)
    );
    MUX_UNSIGNED #(.width(5)) u_mux_1112 (
        .y(_T_322),
        .sel(_T_321),
        .a(_WTEMP_90),
        .b(_T_320)
    );
    wire _T_324;
    EQ_UNSIGNED #(.width(1)) u_eq_1113 (
        .y(_T_324),
        .a(stall),
        .b(1'h0)
    );
    wire _T_325;
    BITWISEAND #(.width(1)) bitwiseand_1114 (
        .y(_T_325),
        .a(_T_324),
        .b(_csr__io_expt)
    );
    wire _T_326;
    BITWISEOR #(.width(1)) bitwiseor_1115 (
        .y(_T_326),
        .a(reset),
        .b(_T_325)
    );
    wire [1:0] _GEN_2;
    wire [1:0] _WTEMP_91;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_1116 (
        .y(_WTEMP_91),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_1117 (
        .y(_GEN_2),
        .sel(_T_326),
        .a(_WTEMP_91),
        .b(_st_type__q)
    );
    wire [2:0] _GEN_3;
    wire [2:0] _WTEMP_92;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_1118 (
        .y(_WTEMP_92),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(3)) u_mux_1119 (
        .y(_GEN_3),
        .sel(_T_326),
        .a(_WTEMP_92),
        .b(_ld_type__q)
    );
    wire _GEN_4;
    MUX_UNSIGNED #(.width(1)) u_mux_1120 (
        .y(_GEN_4),
        .sel(_T_326),
        .a(1'h0),
        .b(_wb_en__q)
    );
    wire [2:0] _GEN_5;
    wire [2:0] _WTEMP_93;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_1121 (
        .y(_WTEMP_93),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(3)) u_mux_1122 (
        .y(_GEN_5),
        .sel(_T_326),
        .a(_WTEMP_93),
        .b(_csr_cmd__q)
    );
    wire _GEN_6;
    MUX_UNSIGNED #(.width(1)) u_mux_1123 (
        .y(_GEN_6),
        .sel(_T_326),
        .a(1'h0),
        .b(_illegal__q)
    );
    wire _GEN_7;
    MUX_UNSIGNED #(.width(1)) u_mux_1124 (
        .y(_GEN_7),
        .sel(_T_326),
        .a(1'h0),
        .b(_pc_check__q)
    );
    wire _T_334;
    EQ_UNSIGNED #(.width(1)) u_eq_1125 (
        .y(_T_334),
        .a(stall),
        .b(1'h0)
    );
    wire _T_336;
    EQ_UNSIGNED #(.width(1)) u_eq_1126 (
        .y(_T_336),
        .a(_csr__io_expt),
        .b(1'h0)
    );
    wire _T_337;
    BITWISEAND #(.width(1)) bitwiseand_1127 (
        .y(_T_337),
        .a(_T_334),
        .b(_T_336)
    );
    wire _T_339;
    EQ_UNSIGNED #(.width(1)) u_eq_1128 (
        .y(_T_339),
        .a(_T_326),
        .b(1'h0)
    );
    wire _T_340;
    BITWISEAND #(.width(1)) bitwiseand_1129 (
        .y(_T_340),
        .a(_T_339),
        .b(_T_337)
    );
    wire _T_341;
    EQ_UNSIGNED #(.width(3)) u_eq_1130 (
        .y(_T_341),
        .a(io_ctrl_imm_sel),
        .b(3'h6)
    );
    wire [31:0] _T_342;
    MUX_UNSIGNED #(.width(32)) u_mux_1131 (
        .y(_T_342),
        .sel(_T_341),
        .a(_immGen__io_out),
        .b(rs1)
    );
    wire _T_343;
    EQ_UNSIGNED #(.width(2)) u_eq_1132 (
        .y(_T_343),
        .a(io_ctrl_pc_sel),
        .b(2'h1)
    );
    wire [32:0] _GEN_8;
    MUX_UNSIGNED #(.width(33)) u_mux_1133 (
        .y(_GEN_8),
        .sel(_T_340),
        .a(_fe_pc__q),
        .b(_ew_pc__q)
    );
    wire [31:0] _GEN_9;
    MUX_UNSIGNED #(.width(32)) u_mux_1134 (
        .y(_GEN_9),
        .sel(_T_340),
        .a(_fe_inst__q),
        .b(_ew_inst__q)
    );
    wire [31:0] _GEN_10;
    MUX_UNSIGNED #(.width(32)) u_mux_1135 (
        .y(_GEN_10),
        .sel(_T_340),
        .a(_alu__io_out),
        .b(_ew_alu__q)
    );
    wire [31:0] _GEN_11;
    MUX_UNSIGNED #(.width(32)) u_mux_1136 (
        .y(_GEN_11),
        .sel(_T_340),
        .a(_T_342),
        .b(_csr_in__q)
    );
    wire [1:0] _GEN_12;
    MUX_UNSIGNED #(.width(2)) u_mux_1137 (
        .y(_GEN_12),
        .sel(_T_340),
        .a(io_ctrl_st_type),
        .b(_GEN_2)
    );
    wire [2:0] _GEN_13;
    MUX_UNSIGNED #(.width(3)) u_mux_1138 (
        .y(_GEN_13),
        .sel(_T_340),
        .a(io_ctrl_ld_type),
        .b(_GEN_3)
    );
    wire [1:0] _GEN_14;
    MUX_UNSIGNED #(.width(2)) u_mux_1139 (
        .y(_GEN_14),
        .sel(_T_340),
        .a(io_ctrl_wb_sel),
        .b(_wb_sel__q)
    );
    wire _GEN_15;
    MUX_UNSIGNED #(.width(1)) u_mux_1140 (
        .y(_GEN_15),
        .sel(_T_340),
        .a(io_ctrl_wb_en),
        .b(_GEN_4)
    );
    wire [2:0] _GEN_16;
    MUX_UNSIGNED #(.width(3)) u_mux_1141 (
        .y(_GEN_16),
        .sel(_T_340),
        .a(io_ctrl_csr_cmd),
        .b(_GEN_5)
    );
    wire _GEN_17;
    MUX_UNSIGNED #(.width(1)) u_mux_1142 (
        .y(_GEN_17),
        .sel(_T_340),
        .a(io_ctrl_illegal),
        .b(_GEN_6)
    );
    wire _GEN_18;
    MUX_UNSIGNED #(.width(1)) u_mux_1143 (
        .y(_GEN_18),
        .sel(_T_340),
        .a(_T_343),
        .b(_GEN_7)
    );
    wire _T_344;
    BITS #(.width(32), .high(1), .low(1)) bits_1144 (
        .y(_T_344),
        .in(_ew_alu__q)
    );
    wire [7:0] _T_346;
    DSHL_UNSIGNED #(.width_in(1), .width_n(3)) u_dshl_1145 (
        .y(_T_346),
        .in(_T_344),
        .n(3'h4)
    );
    wire _T_347;
    BITS #(.width(32), .high(0), .low(0)) bits_1146 (
        .y(_T_347),
        .in(_ew_alu__q)
    );
    wire [3:0] _T_349;
    DSHL_UNSIGNED #(.width_in(1), .width_n(2)) u_dshl_1147 (
        .y(_T_349),
        .in(_T_347),
        .n(2'h3)
    );
    wire [7:0] loffset;
    wire [7:0] _WTEMP_94;
    PAD_UNSIGNED #(.width(4), .n(8)) u_pad_1148 (
        .y(_WTEMP_94),
        .in(_T_349)
    );
    BITWISEOR #(.width(8)) bitwiseor_1149 (
        .y(loffset),
        .a(_T_346),
        .b(_WTEMP_94)
    );
    wire [31:0] lshift;
    DSHR_UNSIGNED #(.width_in(32), .width_n(8)) u_dshr_1150 (
        .y(lshift),
        .in(io_dcache_resp_bits_data),
        .n(loffset)
    );
    wire [32:0] _T_350;
    CVT_UNSIGNED #(.width(32)) u_cvt_1151 (
        .y(_T_350),
        .in(io_dcache_resp_bits_data)
    );
    wire [15:0] _T_351;
    BITS #(.width(32), .high(15), .low(0)) bits_1152 (
        .y(_T_351),
        .in(lshift)
    );
    wire [15:0] _T_352;
    ASSINT #(.width(16)) assint_1153 (
        .y(_T_352),
        .in(_T_351)
    );
    wire [7:0] _T_353;
    BITS #(.width(32), .high(7), .low(0)) bits_1154 (
        .y(_T_353),
        .in(lshift)
    );
    wire [7:0] _T_354;
    ASSINT #(.width(8)) assint_1155 (
        .y(_T_354),
        .in(_T_353)
    );
    wire [15:0] _T_355;
    BITS #(.width(32), .high(15), .low(0)) bits_1156 (
        .y(_T_355),
        .in(lshift)
    );
    wire [16:0] _T_356;
    CVT_UNSIGNED #(.width(16)) u_cvt_1157 (
        .y(_T_356),
        .in(_T_355)
    );
    wire [7:0] _T_357;
    BITS #(.width(32), .high(7), .low(0)) bits_1158 (
        .y(_T_357),
        .in(lshift)
    );
    wire [8:0] _T_358;
    CVT_UNSIGNED #(.width(8)) u_cvt_1159 (
        .y(_T_358),
        .in(_T_357)
    );
    wire _T_359;
    EQ_UNSIGNED #(.width(3)) u_eq_1160 (
        .y(_T_359),
        .a(3'h5),
        .b(_ld_type__q)
    );
    wire [32:0] _T_360;
    wire [32:0] _WTEMP_95;
    PAD_SIGNED #(.width(9), .n(33)) s_pad_1161 (
        .y(_WTEMP_95),
        .in(_T_358)
    );
    MUX_SIGNED #(.width(33)) s_mux_1162 (
        .y(_T_360),
        .sel(_T_359),
        .a(_WTEMP_95),
        .b(_T_350)
    );
    wire _T_361;
    EQ_UNSIGNED #(.width(3)) u_eq_1163 (
        .y(_T_361),
        .a(3'h4),
        .b(_ld_type__q)
    );
    wire [32:0] _T_362;
    wire [32:0] _WTEMP_96;
    PAD_SIGNED #(.width(17), .n(33)) s_pad_1164 (
        .y(_WTEMP_96),
        .in(_T_356)
    );
    MUX_SIGNED #(.width(33)) s_mux_1165 (
        .y(_T_362),
        .sel(_T_361),
        .a(_WTEMP_96),
        .b(_T_360)
    );
    wire _T_363;
    EQ_UNSIGNED #(.width(3)) u_eq_1166 (
        .y(_T_363),
        .a(3'h3),
        .b(_ld_type__q)
    );
    wire [32:0] _T_364;
    wire [32:0] _WTEMP_97;
    PAD_SIGNED #(.width(8), .n(33)) s_pad_1167 (
        .y(_WTEMP_97),
        .in(_T_354)
    );
    MUX_SIGNED #(.width(33)) s_mux_1168 (
        .y(_T_364),
        .sel(_T_363),
        .a(_WTEMP_97),
        .b(_T_362)
    );
    wire _T_365;
    EQ_UNSIGNED #(.width(3)) u_eq_1169 (
        .y(_T_365),
        .a(3'h2),
        .b(_ld_type__q)
    );
    wire [32:0] load;
    wire [32:0] _WTEMP_98;
    PAD_SIGNED #(.width(16), .n(33)) s_pad_1170 (
        .y(_WTEMP_98),
        .in(_T_352)
    );
    MUX_SIGNED #(.width(33)) s_mux_1171 (
        .y(load),
        .sel(_T_365),
        .a(_WTEMP_98),
        .b(_T_364)
    );
    wire [32:0] _T_366;
    CVT_UNSIGNED #(.width(32)) u_cvt_1172 (
        .y(_T_366),
        .in(_ew_alu__q)
    );
    wire [33:0] _T_368;
    wire [32:0] _WTEMP_99;
    PAD_UNSIGNED #(.width(3), .n(33)) u_pad_1173 (
        .y(_WTEMP_99),
        .in(3'h4)
    );
    ADD_UNSIGNED #(.width(33)) u_add_1174 (
        .y(_T_368),
        .a(_ew_pc__q),
        .b(_WTEMP_99)
    );
    wire [32:0] _T_369;
    TAIL #(.width(34), .n(1)) tail_1175 (
        .y(_T_369),
        .in(_T_368)
    );
    wire [33:0] _T_370;
    CVT_UNSIGNED #(.width(33)) u_cvt_1176 (
        .y(_T_370),
        .in(_T_369)
    );
    wire [32:0] _T_371;
    CVT_UNSIGNED #(.width(32)) u_cvt_1177 (
        .y(_T_371),
        .in(_csr__io_out)
    );
    wire _T_372;
    EQ_UNSIGNED #(.width(2)) u_eq_1178 (
        .y(_T_372),
        .a(2'h3),
        .b(_wb_sel__q)
    );
    wire [32:0] _T_373;
    MUX_SIGNED #(.width(33)) s_mux_1179 (
        .y(_T_373),
        .sel(_T_372),
        .a(_T_371),
        .b(_T_366)
    );
    wire _T_374;
    EQ_UNSIGNED #(.width(2)) u_eq_1180 (
        .y(_T_374),
        .a(2'h2),
        .b(_wb_sel__q)
    );
    wire [33:0] _T_375;
    wire [33:0] _WTEMP_100;
    PAD_SIGNED #(.width(33), .n(34)) s_pad_1181 (
        .y(_WTEMP_100),
        .in(_T_373)
    );
    MUX_SIGNED #(.width(34)) s_mux_1182 (
        .y(_T_375),
        .sel(_T_374),
        .a(_T_370),
        .b(_WTEMP_100)
    );
    wire _T_376;
    EQ_UNSIGNED #(.width(2)) u_eq_1183 (
        .y(_T_376),
        .a(2'h1),
        .b(_wb_sel__q)
    );
    wire [33:0] _T_377;
    wire [33:0] _WTEMP_101;
    PAD_SIGNED #(.width(33), .n(34)) s_pad_1184 (
        .y(_WTEMP_101),
        .in(load)
    );
    MUX_SIGNED #(.width(34)) s_mux_1185 (
        .y(_T_377),
        .sel(_T_376),
        .a(_WTEMP_101),
        .b(_T_375)
    );
    wire [33:0] regWrite;
    ASUINT #(.width(34)) asuint_1186 (
        .y(regWrite),
        .in(_T_377)
    );
    wire _T_379;
    EQ_UNSIGNED #(.width(1)) u_eq_1187 (
        .y(_T_379),
        .a(stall),
        .b(1'h0)
    );
    wire _T_380;
    BITWISEAND #(.width(1)) bitwiseand_1188 (
        .y(_T_380),
        .a(_wb_en__q),
        .b(_T_379)
    );
    wire _T_382;
    EQ_UNSIGNED #(.width(1)) u_eq_1189 (
        .y(_T_382),
        .a(_csr__io_expt),
        .b(1'h0)
    );
    wire _T_383;
    BITWISEAND #(.width(1)) bitwiseand_1190 (
        .y(_T_383),
        .a(_T_380),
        .b(_T_382)
    );
    assign _alu__clock = clock;
    BITS #(.width(33), .high(31), .low(0)) bits_1191 (
        .y(_alu__io_A),
        .in(_T_286)
    );
    assign _alu__io_B = _T_288;
    assign _alu__io_alu_op = io_ctrl_alu_op;
    assign _alu__reset = reset;
    assign _brCond__clock = clock;
    assign _brCond__io_br_type = io_ctrl_br_type;
    assign _brCond__io_rs1 = rs1;
    assign _brCond__io_rs2 = rs2;
    assign _brCond__reset = reset;
    assign _csr__clock = clock;
    assign _csr__io_addr = _ew_alu__q;
    assign _csr__io_cmd = _csr_cmd__q;
    assign _csr__io_host_fromhost_bits = io_host_fromhost_bits;
    assign _csr__io_host_fromhost_valid = io_host_fromhost_valid;
    assign _csr__io_illegal = _illegal__q;
    assign _csr__io_in = _csr_in__q;
    assign _csr__io_inst = _ew_inst__q;
    assign _csr__io_ld_type = _ld_type__q;
    BITS #(.width(33), .high(31), .low(0)) bits_1192 (
        .y(_csr__io_pc),
        .in(_ew_pc__q)
    );
    assign _csr__io_pc_check = _pc_check__q;
    assign _csr__io_st_type = _st_type__q;
    assign _csr__io_stall = stall;
    assign _csr__reset = reset;
    assign _csr_cmd__d = _GEN_16;
    assign _csr_in__d = _GEN_11;
    assign _ew_alu__d = _GEN_10;
    MUX_UNSIGNED #(.width(32)) u_mux_1193 (
        .y(_ew_inst__d),
        .sel(reset),
        .a(32'h13),
        .b(_GEN_9)
    );
    assign _ew_pc__d = _GEN_8;
    MUX_UNSIGNED #(.width(32)) u_mux_1194 (
        .y(_fe_inst__d),
        .sel(reset),
        .a(32'h13),
        .b(_GEN_1)
    );
    assign _fe_pc__d = _GEN_0;
    assign _illegal__d = _GEN_17;
    assign _immGen__clock = clock;
    assign _immGen__io_inst = _fe_inst__q;
    assign _immGen__io_sel = io_ctrl_imm_sel;
    assign _immGen__reset = reset;
    assign io_ctrl_inst = _fe_inst__q;
    assign io_dcache_abort = _csr__io_expt;
    BITS #(.width(35), .high(31), .low(0)) bits_1195 (
        .y(io_dcache_req_bits_addr),
        .in(daddr)
    );
    BITS #(.width(287), .high(31), .low(0)) bits_1196 (
        .y(io_dcache_req_bits_data),
        .in(_T_307)
    );
    BITS #(.width(5), .high(3), .low(0)) bits_1197 (
        .y(io_dcache_req_bits_mask),
        .in(_T_322)
    );
    assign io_dcache_req_valid = _T_306;
    assign io_host_tohost = _csr__io_host_tohost;
    assign io_icache_abort = 1'h0;
    BITS #(.width(33), .high(31), .low(0)) bits_1198 (
        .y(io_icache_req_bits_addr),
        .in(npc)
    );
    PAD_UNSIGNED #(.width(1), .n(32)) u_pad_1199 (
        .y(io_icache_req_bits_data),
        .in(1'h0)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1200 (
        .y(io_icache_req_bits_mask),
        .in(1'h0)
    );
    assign io_icache_req_valid = _T_269;
    assign _ld_type__d = _GEN_13;
    wire [32:0] _WTEMP_102;
    PAD_UNSIGNED #(.width(32), .n(33)) u_pad_1201 (
        .y(_WTEMP_102),
        .in(_T_246)
    );
    MUX_UNSIGNED #(.width(33)) u_mux_1202 (
        .y(_pc__d),
        .sel(reset),
        .a(_WTEMP_102),
        .b(npc)
    );
    assign _pc_check__d = _GEN_18;
    assign _regFile__clock = clock;
    assign _regFile__io_raddr1 = rs1_addr;
    assign _regFile__io_raddr2 = rs2_addr;
    assign _regFile__io_waddr = wb_rd_addr;
    BITS #(.width(34), .high(31), .low(0)) bits_1203 (
        .y(_regFile__io_wdata),
        .in(regWrite)
    );
    assign _regFile__io_wen = _T_383;
    assign _regFile__reset = reset;
    assign _st_type__d = _GEN_12;
    assign _started__d = reset;
    assign _wb_en__d = _GEN_15;
    assign _wb_sel__d = _GEN_14;
endmodule //Datapath
module CSR(
    input clock,
    input reset,
    input io_stall,
    input [2:0] io_cmd,
    input [31:0] io_in,
    output [31:0] io_out,
    input [31:0] io_pc,
    input [31:0] io_addr,
    input [31:0] io_inst,
    input io_illegal,
    input [1:0] io_st_type,
    input [2:0] io_ld_type,
    input io_pc_check,
    output io_expt,
    output [31:0] io_evec,
    output [31:0] io_epc,
    input io_host_fromhost_valid,
    input [31:0] io_host_fromhost_bits,
    output [31:0] io_host_tohost
);
    wire [31:0] _time___q;
    wire [31:0] _time___d;
    DFF_POSCLK #(.width(32)) time_ (
        .q(_time___q),
        .d(_time___d),
        .clk(clock)
    );
    wire [31:0] _timeh__q;
    wire [31:0] _timeh__d;
    DFF_POSCLK #(.width(32)) timeh (
        .q(_timeh__q),
        .d(_timeh__d),
        .clk(clock)
    );
    wire [31:0] _cycle__q;
    wire [31:0] _cycle__d;
    DFF_POSCLK #(.width(32)) cycle (
        .q(_cycle__q),
        .d(_cycle__d),
        .clk(clock)
    );
    wire [31:0] _cycleh__q;
    wire [31:0] _cycleh__d;
    DFF_POSCLK #(.width(32)) cycleh (
        .q(_cycleh__q),
        .d(_cycleh__d),
        .clk(clock)
    );
    wire [31:0] _instret__q;
    wire [31:0] _instret__d;
    DFF_POSCLK #(.width(32)) instret (
        .q(_instret__q),
        .d(_instret__d),
        .clk(clock)
    );
    wire [31:0] _instreth__q;
    wire [31:0] _instreth__d;
    DFF_POSCLK #(.width(32)) instreth (
        .q(_instreth__q),
        .d(_instreth__d),
        .clk(clock)
    );
    wire [1:0] _PRV__q;
    wire [1:0] _PRV__d;
    DFF_POSCLK #(.width(2)) PRV (
        .q(_PRV__q),
        .d(_PRV__d),
        .clk(clock)
    );
    wire [1:0] _PRV1__q;
    wire [1:0] _PRV1__d;
    DFF_POSCLK #(.width(2)) PRV1 (
        .q(_PRV1__q),
        .d(_PRV1__d),
        .clk(clock)
    );
    wire _IE__q;
    wire _IE__d;
    DFF_POSCLK #(.width(1)) IE (
        .q(_IE__q),
        .d(_IE__d),
        .clk(clock)
    );
    wire _IE1__q;
    wire _IE1__d;
    DFF_POSCLK #(.width(1)) IE1 (
        .q(_IE1__q),
        .d(_IE1__d),
        .clk(clock)
    );
    wire _MTIP__q;
    wire _MTIP__d;
    DFF_POSCLK #(.width(1)) MTIP (
        .q(_MTIP__q),
        .d(_MTIP__d),
        .clk(clock)
    );
    wire _MTIE__q;
    wire _MTIE__d;
    DFF_POSCLK #(.width(1)) MTIE (
        .q(_MTIE__q),
        .d(_MTIE__d),
        .clk(clock)
    );
    wire _MSIP__q;
    wire _MSIP__d;
    DFF_POSCLK #(.width(1)) MSIP (
        .q(_MSIP__q),
        .d(_MSIP__d),
        .clk(clock)
    );
    wire _MSIE__q;
    wire _MSIE__d;
    DFF_POSCLK #(.width(1)) MSIE (
        .q(_MSIE__q),
        .d(_MSIE__d),
        .clk(clock)
    );
    wire [31:0] _mtimecmp__q;
    wire [31:0] _mtimecmp__d;
    DFF_POSCLK #(.width(32)) mtimecmp (
        .q(_mtimecmp__q),
        .d(_mtimecmp__d),
        .clk(clock)
    );
    wire [31:0] _mscratch__q;
    wire [31:0] _mscratch__d;
    DFF_POSCLK #(.width(32)) mscratch (
        .q(_mscratch__q),
        .d(_mscratch__d),
        .clk(clock)
    );
    wire [31:0] _mepc__q;
    wire [31:0] _mepc__d;
    DFF_POSCLK #(.width(32)) mepc (
        .q(_mepc__q),
        .d(_mepc__d),
        .clk(clock)
    );
    wire [31:0] _mcause__q;
    wire [31:0] _mcause__d;
    DFF_POSCLK #(.width(32)) mcause (
        .q(_mcause__q),
        .d(_mcause__d),
        .clk(clock)
    );
    wire [31:0] _mbadaddr__q;
    wire [31:0] _mbadaddr__d;
    DFF_POSCLK #(.width(32)) mbadaddr (
        .q(_mbadaddr__q),
        .d(_mbadaddr__d),
        .clk(clock)
    );
    wire [31:0] _mtohost__q;
    wire [31:0] _mtohost__d;
    DFF_POSCLK #(.width(32)) mtohost (
        .q(_mtohost__q),
        .d(_mtohost__d),
        .clk(clock)
    );
    wire [31:0] _mfromhost__q;
    wire [31:0] _mfromhost__d;
    DFF_POSCLK #(.width(32)) mfromhost (
        .q(_mfromhost__q),
        .d(_mfromhost__d),
        .clk(clock)
    );
    wire [11:0] csr_addr;
    BITS #(.width(32), .high(31), .low(20)) bits_1 (
        .y(csr_addr),
        .in(io_inst)
    );
    wire [4:0] rs1_addr;
    BITS #(.width(32), .high(19), .low(15)) bits_2 (
        .y(rs1_addr),
        .in(io_inst)
    );
    wire [5:0] _T_53;
    assign _T_53 = 6'h0;
    wire [31:0] mcpuid;
    assign mcpuid = 32'h100100;
    wire [2:0] _T_93;
    CAT #(.width_a(1), .width_b(2)) cat_3 (
        .y(_T_93),
        .a(_IE1__q),
        .b(_PRV__q)
    );
    wire [3:0] _T_94;
    CAT #(.width_a(3), .width_b(1)) cat_4 (
        .y(_T_94),
        .a(_T_93),
        .b(_IE__q)
    );
    wire [2:0] _T_95;
    CAT #(.width_a(1), .width_b(2)) cat_5 (
        .y(_T_95),
        .a(1'h0),
        .b(_PRV1__q)
    );
    wire [2:0] _T_96;
    assign _T_96 = 3'h0;
    wire [5:0] _T_97;
    CAT #(.width_a(3), .width_b(3)) cat_6 (
        .y(_T_97),
        .a(_T_96),
        .b(_T_95)
    );
    wire [9:0] _T_98;
    CAT #(.width_a(6), .width_b(4)) cat_7 (
        .y(_T_98),
        .a(_T_97),
        .b(_T_94)
    );
    wire [3:0] _T_99;
    assign _T_99 = 4'h0;
    wire [5:0] _T_100;
    assign _T_100 = 6'h0;
    wire [5:0] _T_101;
    assign _T_101 = 6'h0;
    wire [9:0] _T_102;
    assign _T_102 = 10'h0;
    wire [15:0] _T_103;
    assign _T_103 = 16'h0;
    wire [21:0] _T_104;
    assign _T_104 = 22'h0;
    wire [31:0] mstatus;
    CAT #(.width_a(22), .width_b(10)) cat_8 (
        .y(mstatus),
        .a(_T_104),
        .b(_T_98)
    );
    wire [1:0] _T_112;
    assign _T_112 = 2'h0;
    wire [1:0] _T_113;
    CAT #(.width_a(1), .width_b(1)) cat_9 (
        .y(_T_113),
        .a(_MSIP__q),
        .b(1'h0)
    );
    wire [3:0] _T_114;
    CAT #(.width_a(2), .width_b(2)) cat_10 (
        .y(_T_114),
        .a(_T_113),
        .b(_T_112)
    );
    wire [1:0] _T_115;
    assign _T_115 = 2'h0;
    wire [24:0] _T_116;
    CAT #(.width_a(24), .width_b(1)) cat_11 (
        .y(_T_116),
        .a(24'h0),
        .b(_MTIP__q)
    );
    wire [25:0] _T_117;
    CAT #(.width_a(25), .width_b(1)) cat_12 (
        .y(_T_117),
        .a(_T_116),
        .b(1'h0)
    );
    wire [27:0] _T_118;
    CAT #(.width_a(26), .width_b(2)) cat_13 (
        .y(_T_118),
        .a(_T_117),
        .b(_T_115)
    );
    wire [31:0] mip;
    CAT #(.width_a(28), .width_b(4)) cat_14 (
        .y(mip),
        .a(_T_118),
        .b(_T_114)
    );
    wire [1:0] _T_122;
    assign _T_122 = 2'h0;
    wire [1:0] _T_123;
    CAT #(.width_a(1), .width_b(1)) cat_15 (
        .y(_T_123),
        .a(_MSIE__q),
        .b(1'h0)
    );
    wire [3:0] _T_124;
    CAT #(.width_a(2), .width_b(2)) cat_16 (
        .y(_T_124),
        .a(_T_123),
        .b(_T_122)
    );
    wire [1:0] _T_125;
    assign _T_125 = 2'h0;
    wire [24:0] _T_126;
    CAT #(.width_a(24), .width_b(1)) cat_17 (
        .y(_T_126),
        .a(24'h0),
        .b(_MTIE__q)
    );
    wire [25:0] _T_127;
    CAT #(.width_a(25), .width_b(1)) cat_18 (
        .y(_T_127),
        .a(_T_126),
        .b(1'h0)
    );
    wire [27:0] _T_128;
    CAT #(.width_a(26), .width_b(2)) cat_19 (
        .y(_T_128),
        .a(_T_127),
        .b(_T_125)
    );
    wire [31:0] mie;
    CAT #(.width_a(28), .width_b(4)) cat_20 (
        .y(mie),
        .a(_T_128),
        .b(_T_124)
    );
    wire [31:0] _GEN_0;
    MUX_UNSIGNED #(.width(32)) u_mux_21 (
        .y(_GEN_0),
        .sel(io_host_fromhost_valid),
        .a(io_host_fromhost_bits),
        .b(_mfromhost__q)
    );
    wire [11:0] _T_139;
    BITWISEAND #(.width(12)) bitwiseand_22 (
        .y(_T_139),
        .a(csr_addr),
        .b(12'hFFF)
    );
    wire _T_140;
    EQ_UNSIGNED #(.width(12)) u_eq_23 (
        .y(_T_140),
        .a(12'hC00),
        .b(_T_139)
    );
    wire [11:0] _T_143;
    BITWISEAND #(.width(12)) bitwiseand_24 (
        .y(_T_143),
        .a(csr_addr),
        .b(12'hFFF)
    );
    wire _T_144;
    EQ_UNSIGNED #(.width(12)) u_eq_25 (
        .y(_T_144),
        .a(12'hC01),
        .b(_T_143)
    );
    wire [11:0] _T_147;
    BITWISEAND #(.width(12)) bitwiseand_26 (
        .y(_T_147),
        .a(csr_addr),
        .b(12'hFFF)
    );
    wire _T_148;
    EQ_UNSIGNED #(.width(12)) u_eq_27 (
        .y(_T_148),
        .a(12'hC02),
        .b(_T_147)
    );
    wire [11:0] _T_151;
    BITWISEAND #(.width(12)) bitwiseand_28 (
        .y(_T_151),
        .a(csr_addr),
        .b(12'hFFF)
    );
    wire _T_152;
    EQ_UNSIGNED #(.width(12)) u_eq_29 (
        .y(_T_152),
        .a(12'hC80),
        .b(_T_151)
    );
    wire [11:0] _T_155;
    BITWISEAND #(.width(12)) bitwiseand_30 (
        .y(_T_155),
        .a(csr_addr),
        .b(12'hFFF)
    );
    wire _T_156;
    EQ_UNSIGNED #(.width(12)) u_eq_31 (
        .y(_T_156),
        .a(12'hC81),
        .b(_T_155)
    );
    wire [11:0] _T_159;
    BITWISEAND #(.width(12)) bitwiseand_32 (
        .y(_T_159),
        .a(csr_addr),
        .b(12'hFFF)
    );
    wire _T_160;
    EQ_UNSIGNED #(.width(12)) u_eq_33 (
        .y(_T_160),
        .a(12'hC82),
        .b(_T_159)
    );
    wire [11:0] _T_163;
    BITWISEAND #(.width(12)) bitwiseand_34 (
        .y(_T_163),
        .a(csr_addr),
        .b(12'hFFF)
    );
    wire _T_164;
    EQ_UNSIGNED #(.width(12)) u_eq_35 (
        .y(_T_164),
        .a(12'h900),
        .b(_T_163)
    );
    wire [11:0] _T_167;
    BITWISEAND #(.width(12)) bitwiseand_36 (
        .y(_T_167),
        .a(csr_addr),
        .b(12'hFFF)
    );
    wire _T_168;
    EQ_UNSIGNED #(.width(12)) u_eq_37 (
        .y(_T_168),
        .a(12'h901),
        .b(_T_167)
    );
    wire [11:0] _T_171;
    BITWISEAND #(.width(12)) bitwiseand_38 (
        .y(_T_171),
        .a(csr_addr),
        .b(12'hFFF)
    );
    wire _T_172;
    EQ_UNSIGNED #(.width(12)) u_eq_39 (
        .y(_T_172),
        .a(12'h902),
        .b(_T_171)
    );
    wire [11:0] _T_175;
    BITWISEAND #(.width(12)) bitwiseand_40 (
        .y(_T_175),
        .a(csr_addr),
        .b(12'hFFF)
    );
    wire _T_176;
    EQ_UNSIGNED #(.width(12)) u_eq_41 (
        .y(_T_176),
        .a(12'h980),
        .b(_T_175)
    );
    wire [11:0] _T_179;
    BITWISEAND #(.width(12)) bitwiseand_42 (
        .y(_T_179),
        .a(csr_addr),
        .b(12'hFFF)
    );
    wire _T_180;
    EQ_UNSIGNED #(.width(12)) u_eq_43 (
        .y(_T_180),
        .a(12'h981),
        .b(_T_179)
    );
    wire [11:0] _T_183;
    BITWISEAND #(.width(12)) bitwiseand_44 (
        .y(_T_183),
        .a(csr_addr),
        .b(12'hFFF)
    );
    wire _T_184;
    EQ_UNSIGNED #(.width(12)) u_eq_45 (
        .y(_T_184),
        .a(12'h982),
        .b(_T_183)
    );
    wire [11:0] _T_187;
    BITWISEAND #(.width(12)) bitwiseand_46 (
        .y(_T_187),
        .a(csr_addr),
        .b(12'hFFF)
    );
    wire _T_188;
    EQ_UNSIGNED #(.width(12)) u_eq_47 (
        .y(_T_188),
        .a(12'hF00),
        .b(_T_187)
    );
    wire [11:0] _T_191;
    BITWISEAND #(.width(12)) bitwiseand_48 (
        .y(_T_191),
        .a(csr_addr),
        .b(12'hFFF)
    );
    wire _T_192;
    EQ_UNSIGNED #(.width(12)) u_eq_49 (
        .y(_T_192),
        .a(12'hF01),
        .b(_T_191)
    );
    wire [11:0] _T_195;
    BITWISEAND #(.width(12)) bitwiseand_50 (
        .y(_T_195),
        .a(csr_addr),
        .b(12'hFFF)
    );
    wire _T_196;
    EQ_UNSIGNED #(.width(12)) u_eq_51 (
        .y(_T_196),
        .a(12'hF10),
        .b(_T_195)
    );
    wire [11:0] _T_199;
    BITWISEAND #(.width(12)) bitwiseand_52 (
        .y(_T_199),
        .a(csr_addr),
        .b(12'hFFF)
    );
    wire _T_200;
    wire [11:0] _WTEMP_0;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_53 (
        .y(_WTEMP_0),
        .in(10'h301)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_54 (
        .y(_T_200),
        .a(_WTEMP_0),
        .b(_T_199)
    );
    wire [11:0] _T_203;
    BITWISEAND #(.width(12)) bitwiseand_55 (
        .y(_T_203),
        .a(csr_addr),
        .b(12'hFFF)
    );
    wire _T_204;
    wire [11:0] _WTEMP_1;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_56 (
        .y(_WTEMP_1),
        .in(10'h302)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_57 (
        .y(_T_204),
        .a(_WTEMP_1),
        .b(_T_203)
    );
    wire [11:0] _T_207;
    BITWISEAND #(.width(12)) bitwiseand_58 (
        .y(_T_207),
        .a(csr_addr),
        .b(12'hFFF)
    );
    wire _T_208;
    wire [11:0] _WTEMP_2;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_59 (
        .y(_WTEMP_2),
        .in(10'h304)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_60 (
        .y(_T_208),
        .a(_WTEMP_2),
        .b(_T_207)
    );
    wire [11:0] _T_211;
    BITWISEAND #(.width(12)) bitwiseand_61 (
        .y(_T_211),
        .a(csr_addr),
        .b(12'hFFF)
    );
    wire _T_212;
    wire [11:0] _WTEMP_3;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_62 (
        .y(_WTEMP_3),
        .in(10'h321)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_63 (
        .y(_T_212),
        .a(_WTEMP_3),
        .b(_T_211)
    );
    wire [11:0] _T_215;
    BITWISEAND #(.width(12)) bitwiseand_64 (
        .y(_T_215),
        .a(csr_addr),
        .b(12'hFFF)
    );
    wire _T_216;
    wire [11:0] _WTEMP_4;
    PAD_UNSIGNED #(.width(11), .n(12)) u_pad_65 (
        .y(_WTEMP_4),
        .in(11'h701)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_66 (
        .y(_T_216),
        .a(_WTEMP_4),
        .b(_T_215)
    );
    wire [11:0] _T_219;
    BITWISEAND #(.width(12)) bitwiseand_67 (
        .y(_T_219),
        .a(csr_addr),
        .b(12'hFFF)
    );
    wire _T_220;
    wire [11:0] _WTEMP_5;
    PAD_UNSIGNED #(.width(11), .n(12)) u_pad_68 (
        .y(_WTEMP_5),
        .in(11'h741)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_69 (
        .y(_T_220),
        .a(_WTEMP_5),
        .b(_T_219)
    );
    wire [11:0] _T_223;
    BITWISEAND #(.width(12)) bitwiseand_70 (
        .y(_T_223),
        .a(csr_addr),
        .b(12'hFFF)
    );
    wire _T_224;
    wire [11:0] _WTEMP_6;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_71 (
        .y(_WTEMP_6),
        .in(10'h340)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_72 (
        .y(_T_224),
        .a(_WTEMP_6),
        .b(_T_223)
    );
    wire [11:0] _T_227;
    BITWISEAND #(.width(12)) bitwiseand_73 (
        .y(_T_227),
        .a(csr_addr),
        .b(12'hFFF)
    );
    wire _T_228;
    wire [11:0] _WTEMP_7;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_74 (
        .y(_WTEMP_7),
        .in(10'h341)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_75 (
        .y(_T_228),
        .a(_WTEMP_7),
        .b(_T_227)
    );
    wire [11:0] _T_231;
    BITWISEAND #(.width(12)) bitwiseand_76 (
        .y(_T_231),
        .a(csr_addr),
        .b(12'hFFF)
    );
    wire _T_232;
    wire [11:0] _WTEMP_8;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_77 (
        .y(_WTEMP_8),
        .in(10'h342)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_78 (
        .y(_T_232),
        .a(_WTEMP_8),
        .b(_T_231)
    );
    wire [11:0] _T_235;
    BITWISEAND #(.width(12)) bitwiseand_79 (
        .y(_T_235),
        .a(csr_addr),
        .b(12'hFFF)
    );
    wire _T_236;
    wire [11:0] _WTEMP_9;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_80 (
        .y(_WTEMP_9),
        .in(10'h343)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_81 (
        .y(_T_236),
        .a(_WTEMP_9),
        .b(_T_235)
    );
    wire [11:0] _T_239;
    BITWISEAND #(.width(12)) bitwiseand_82 (
        .y(_T_239),
        .a(csr_addr),
        .b(12'hFFF)
    );
    wire _T_240;
    wire [11:0] _WTEMP_10;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_83 (
        .y(_WTEMP_10),
        .in(10'h344)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_84 (
        .y(_T_240),
        .a(_WTEMP_10),
        .b(_T_239)
    );
    wire [11:0] _T_243;
    BITWISEAND #(.width(12)) bitwiseand_85 (
        .y(_T_243),
        .a(csr_addr),
        .b(12'hFFF)
    );
    wire _T_244;
    wire [11:0] _WTEMP_11;
    PAD_UNSIGNED #(.width(11), .n(12)) u_pad_86 (
        .y(_WTEMP_11),
        .in(11'h780)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_87 (
        .y(_T_244),
        .a(_WTEMP_11),
        .b(_T_243)
    );
    wire [11:0] _T_247;
    BITWISEAND #(.width(12)) bitwiseand_88 (
        .y(_T_247),
        .a(csr_addr),
        .b(12'hFFF)
    );
    wire _T_248;
    wire [11:0] _WTEMP_12;
    PAD_UNSIGNED #(.width(11), .n(12)) u_pad_89 (
        .y(_WTEMP_12),
        .in(11'h781)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_90 (
        .y(_T_248),
        .a(_WTEMP_12),
        .b(_T_247)
    );
    wire [11:0] _T_251;
    BITWISEAND #(.width(12)) bitwiseand_91 (
        .y(_T_251),
        .a(csr_addr),
        .b(12'hFFF)
    );
    wire _T_252;
    wire [11:0] _WTEMP_13;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_92 (
        .y(_WTEMP_13),
        .in(10'h300)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_93 (
        .y(_T_252),
        .a(_WTEMP_13),
        .b(_T_251)
    );
    wire [31:0] _T_253;
    wire [31:0] _WTEMP_14;
    PAD_UNSIGNED #(.width(1), .n(32)) u_pad_94 (
        .y(_WTEMP_14),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(32)) u_mux_95 (
        .y(_T_253),
        .sel(_T_252),
        .a(mstatus),
        .b(_WTEMP_14)
    );
    wire [31:0] _T_254;
    MUX_UNSIGNED #(.width(32)) u_mux_96 (
        .y(_T_254),
        .sel(_T_248),
        .a(_mfromhost__q),
        .b(_T_253)
    );
    wire [31:0] _T_255;
    MUX_UNSIGNED #(.width(32)) u_mux_97 (
        .y(_T_255),
        .sel(_T_244),
        .a(_mtohost__q),
        .b(_T_254)
    );
    wire [31:0] _T_256;
    MUX_UNSIGNED #(.width(32)) u_mux_98 (
        .y(_T_256),
        .sel(_T_240),
        .a(mip),
        .b(_T_255)
    );
    wire [31:0] _T_257;
    MUX_UNSIGNED #(.width(32)) u_mux_99 (
        .y(_T_257),
        .sel(_T_236),
        .a(_mbadaddr__q),
        .b(_T_256)
    );
    wire [31:0] _T_258;
    MUX_UNSIGNED #(.width(32)) u_mux_100 (
        .y(_T_258),
        .sel(_T_232),
        .a(_mcause__q),
        .b(_T_257)
    );
    wire [31:0] _T_259;
    MUX_UNSIGNED #(.width(32)) u_mux_101 (
        .y(_T_259),
        .sel(_T_228),
        .a(_mepc__q),
        .b(_T_258)
    );
    wire [31:0] _T_260;
    MUX_UNSIGNED #(.width(32)) u_mux_102 (
        .y(_T_260),
        .sel(_T_224),
        .a(_mscratch__q),
        .b(_T_259)
    );
    wire [31:0] _T_261;
    MUX_UNSIGNED #(.width(32)) u_mux_103 (
        .y(_T_261),
        .sel(_T_220),
        .a(_timeh__q),
        .b(_T_260)
    );
    wire [31:0] _T_262;
    MUX_UNSIGNED #(.width(32)) u_mux_104 (
        .y(_T_262),
        .sel(_T_216),
        .a(_time___q),
        .b(_T_261)
    );
    wire [31:0] _T_263;
    MUX_UNSIGNED #(.width(32)) u_mux_105 (
        .y(_T_263),
        .sel(_T_212),
        .a(_mtimecmp__q),
        .b(_T_262)
    );
    wire [31:0] _T_264;
    MUX_UNSIGNED #(.width(32)) u_mux_106 (
        .y(_T_264),
        .sel(_T_208),
        .a(mie),
        .b(_T_263)
    );
    wire [31:0] _T_265;
    MUX_UNSIGNED #(.width(32)) u_mux_107 (
        .y(_T_265),
        .sel(_T_204),
        .a(32'h0),
        .b(_T_264)
    );
    wire [31:0] _T_266;
    MUX_UNSIGNED #(.width(32)) u_mux_108 (
        .y(_T_266),
        .sel(_T_200),
        .a(32'h100),
        .b(_T_265)
    );
    wire [31:0] _T_267;
    MUX_UNSIGNED #(.width(32)) u_mux_109 (
        .y(_T_267),
        .sel(_T_196),
        .a(32'h0),
        .b(_T_266)
    );
    wire [31:0] _T_268;
    MUX_UNSIGNED #(.width(32)) u_mux_110 (
        .y(_T_268),
        .sel(_T_192),
        .a(32'h0),
        .b(_T_267)
    );
    wire [31:0] _T_269;
    MUX_UNSIGNED #(.width(32)) u_mux_111 (
        .y(_T_269),
        .sel(_T_188),
        .a(mcpuid),
        .b(_T_268)
    );
    wire [31:0] _T_270;
    MUX_UNSIGNED #(.width(32)) u_mux_112 (
        .y(_T_270),
        .sel(_T_184),
        .a(_instreth__q),
        .b(_T_269)
    );
    wire [31:0] _T_271;
    MUX_UNSIGNED #(.width(32)) u_mux_113 (
        .y(_T_271),
        .sel(_T_180),
        .a(_timeh__q),
        .b(_T_270)
    );
    wire [31:0] _T_272;
    MUX_UNSIGNED #(.width(32)) u_mux_114 (
        .y(_T_272),
        .sel(_T_176),
        .a(_cycleh__q),
        .b(_T_271)
    );
    wire [31:0] _T_273;
    MUX_UNSIGNED #(.width(32)) u_mux_115 (
        .y(_T_273),
        .sel(_T_172),
        .a(_instret__q),
        .b(_T_272)
    );
    wire [31:0] _T_274;
    MUX_UNSIGNED #(.width(32)) u_mux_116 (
        .y(_T_274),
        .sel(_T_168),
        .a(_time___q),
        .b(_T_273)
    );
    wire [31:0] _T_275;
    MUX_UNSIGNED #(.width(32)) u_mux_117 (
        .y(_T_275),
        .sel(_T_164),
        .a(_cycle__q),
        .b(_T_274)
    );
    wire [31:0] _T_276;
    MUX_UNSIGNED #(.width(32)) u_mux_118 (
        .y(_T_276),
        .sel(_T_160),
        .a(_instreth__q),
        .b(_T_275)
    );
    wire [31:0] _T_277;
    MUX_UNSIGNED #(.width(32)) u_mux_119 (
        .y(_T_277),
        .sel(_T_156),
        .a(_timeh__q),
        .b(_T_276)
    );
    wire [31:0] _T_278;
    MUX_UNSIGNED #(.width(32)) u_mux_120 (
        .y(_T_278),
        .sel(_T_152),
        .a(_cycleh__q),
        .b(_T_277)
    );
    wire [31:0] _T_279;
    MUX_UNSIGNED #(.width(32)) u_mux_121 (
        .y(_T_279),
        .sel(_T_148),
        .a(_instret__q),
        .b(_T_278)
    );
    wire [31:0] _T_280;
    MUX_UNSIGNED #(.width(32)) u_mux_122 (
        .y(_T_280),
        .sel(_T_144),
        .a(_time___q),
        .b(_T_279)
    );
    wire [31:0] _T_281;
    MUX_UNSIGNED #(.width(32)) u_mux_123 (
        .y(_T_281),
        .sel(_T_140),
        .a(_cycle__q),
        .b(_T_280)
    );
    wire [1:0] _T_282;
    BITS #(.width(12), .high(9), .low(8)) bits_124 (
        .y(_T_282),
        .in(csr_addr)
    );
    wire privValid;
    LEQ_UNSIGNED #(.width(2)) u_leq_125 (
        .y(privValid),
        .a(_T_282),
        .b(_PRV__q)
    );
    wire privInst;
    EQ_UNSIGNED #(.width(3)) u_eq_126 (
        .y(privInst),
        .a(io_cmd),
        .b(3'h4)
    );
    wire _T_283;
    BITS #(.width(12), .high(0), .low(0)) bits_127 (
        .y(_T_283),
        .in(csr_addr)
    );
    wire _T_285;
    EQ_UNSIGNED #(.width(1)) u_eq_128 (
        .y(_T_285),
        .a(_T_283),
        .b(1'h0)
    );
    wire _T_286;
    BITWISEAND #(.width(1)) bitwiseand_129 (
        .y(_T_286),
        .a(privInst),
        .b(_T_285)
    );
    wire _T_287;
    BITS #(.width(12), .high(8), .low(8)) bits_130 (
        .y(_T_287),
        .in(csr_addr)
    );
    wire _T_289;
    EQ_UNSIGNED #(.width(1)) u_eq_131 (
        .y(_T_289),
        .a(_T_287),
        .b(1'h0)
    );
    wire isEcall;
    BITWISEAND #(.width(1)) bitwiseand_132 (
        .y(isEcall),
        .a(_T_286),
        .b(_T_289)
    );
    wire _T_290;
    BITS #(.width(12), .high(0), .low(0)) bits_133 (
        .y(_T_290),
        .in(csr_addr)
    );
    wire _T_291;
    BITWISEAND #(.width(1)) bitwiseand_134 (
        .y(_T_291),
        .a(privInst),
        .b(_T_290)
    );
    wire _T_292;
    BITS #(.width(12), .high(8), .low(8)) bits_135 (
        .y(_T_292),
        .in(csr_addr)
    );
    wire _T_294;
    EQ_UNSIGNED #(.width(1)) u_eq_136 (
        .y(_T_294),
        .a(_T_292),
        .b(1'h0)
    );
    wire isEbreak;
    BITWISEAND #(.width(1)) bitwiseand_137 (
        .y(isEbreak),
        .a(_T_291),
        .b(_T_294)
    );
    wire _T_295;
    BITS #(.width(12), .high(0), .low(0)) bits_138 (
        .y(_T_295),
        .in(csr_addr)
    );
    wire _T_297;
    EQ_UNSIGNED #(.width(1)) u_eq_139 (
        .y(_T_297),
        .a(_T_295),
        .b(1'h0)
    );
    wire _T_298;
    BITWISEAND #(.width(1)) bitwiseand_140 (
        .y(_T_298),
        .a(privInst),
        .b(_T_297)
    );
    wire _T_299;
    BITS #(.width(12), .high(8), .low(8)) bits_141 (
        .y(_T_299),
        .in(csr_addr)
    );
    wire isEret;
    BITWISEAND #(.width(1)) bitwiseand_142 (
        .y(isEret),
        .a(_T_298),
        .b(_T_299)
    );
    wire [11:0] _T_302;
    BITWISEAND #(.width(12)) bitwiseand_143 (
        .y(_T_302),
        .a(csr_addr),
        .b(12'hFFF)
    );
    wire _T_303;
    EQ_UNSIGNED #(.width(12)) u_eq_144 (
        .y(_T_303),
        .a(12'hC00),
        .b(_T_302)
    );
    wire [11:0] _T_306;
    BITWISEAND #(.width(12)) bitwiseand_145 (
        .y(_T_306),
        .a(csr_addr),
        .b(12'hFFF)
    );
    wire _T_307;
    EQ_UNSIGNED #(.width(12)) u_eq_146 (
        .y(_T_307),
        .a(12'hC01),
        .b(_T_306)
    );
    wire [11:0] _T_310;
    BITWISEAND #(.width(12)) bitwiseand_147 (
        .y(_T_310),
        .a(csr_addr),
        .b(12'hFFF)
    );
    wire _T_311;
    EQ_UNSIGNED #(.width(12)) u_eq_148 (
        .y(_T_311),
        .a(12'hC02),
        .b(_T_310)
    );
    wire [11:0] _T_314;
    BITWISEAND #(.width(12)) bitwiseand_149 (
        .y(_T_314),
        .a(csr_addr),
        .b(12'hFFF)
    );
    wire _T_315;
    EQ_UNSIGNED #(.width(12)) u_eq_150 (
        .y(_T_315),
        .a(12'hC80),
        .b(_T_314)
    );
    wire [11:0] _T_318;
    BITWISEAND #(.width(12)) bitwiseand_151 (
        .y(_T_318),
        .a(csr_addr),
        .b(12'hFFF)
    );
    wire _T_319;
    EQ_UNSIGNED #(.width(12)) u_eq_152 (
        .y(_T_319),
        .a(12'hC81),
        .b(_T_318)
    );
    wire [11:0] _T_322;
    BITWISEAND #(.width(12)) bitwiseand_153 (
        .y(_T_322),
        .a(csr_addr),
        .b(12'hFFF)
    );
    wire _T_323;
    EQ_UNSIGNED #(.width(12)) u_eq_154 (
        .y(_T_323),
        .a(12'hC82),
        .b(_T_322)
    );
    wire [11:0] _T_326;
    BITWISEAND #(.width(12)) bitwiseand_155 (
        .y(_T_326),
        .a(csr_addr),
        .b(12'hFFF)
    );
    wire _T_327;
    EQ_UNSIGNED #(.width(12)) u_eq_156 (
        .y(_T_327),
        .a(12'h900),
        .b(_T_326)
    );
    wire [11:0] _T_330;
    BITWISEAND #(.width(12)) bitwiseand_157 (
        .y(_T_330),
        .a(csr_addr),
        .b(12'hFFF)
    );
    wire _T_331;
    EQ_UNSIGNED #(.width(12)) u_eq_158 (
        .y(_T_331),
        .a(12'h901),
        .b(_T_330)
    );
    wire [11:0] _T_334;
    BITWISEAND #(.width(12)) bitwiseand_159 (
        .y(_T_334),
        .a(csr_addr),
        .b(12'hFFF)
    );
    wire _T_335;
    EQ_UNSIGNED #(.width(12)) u_eq_160 (
        .y(_T_335),
        .a(12'h902),
        .b(_T_334)
    );
    wire [11:0] _T_338;
    BITWISEAND #(.width(12)) bitwiseand_161 (
        .y(_T_338),
        .a(csr_addr),
        .b(12'hFFF)
    );
    wire _T_339;
    EQ_UNSIGNED #(.width(12)) u_eq_162 (
        .y(_T_339),
        .a(12'h980),
        .b(_T_338)
    );
    wire [11:0] _T_342;
    BITWISEAND #(.width(12)) bitwiseand_163 (
        .y(_T_342),
        .a(csr_addr),
        .b(12'hFFF)
    );
    wire _T_343;
    EQ_UNSIGNED #(.width(12)) u_eq_164 (
        .y(_T_343),
        .a(12'h981),
        .b(_T_342)
    );
    wire [11:0] _T_346;
    BITWISEAND #(.width(12)) bitwiseand_165 (
        .y(_T_346),
        .a(csr_addr),
        .b(12'hFFF)
    );
    wire _T_347;
    EQ_UNSIGNED #(.width(12)) u_eq_166 (
        .y(_T_347),
        .a(12'h982),
        .b(_T_346)
    );
    wire [11:0] _T_350;
    BITWISEAND #(.width(12)) bitwiseand_167 (
        .y(_T_350),
        .a(csr_addr),
        .b(12'hFFF)
    );
    wire _T_351;
    EQ_UNSIGNED #(.width(12)) u_eq_168 (
        .y(_T_351),
        .a(12'hF00),
        .b(_T_350)
    );
    wire [11:0] _T_354;
    BITWISEAND #(.width(12)) bitwiseand_169 (
        .y(_T_354),
        .a(csr_addr),
        .b(12'hFFF)
    );
    wire _T_355;
    EQ_UNSIGNED #(.width(12)) u_eq_170 (
        .y(_T_355),
        .a(12'hF01),
        .b(_T_354)
    );
    wire [11:0] _T_358;
    BITWISEAND #(.width(12)) bitwiseand_171 (
        .y(_T_358),
        .a(csr_addr),
        .b(12'hFFF)
    );
    wire _T_359;
    EQ_UNSIGNED #(.width(12)) u_eq_172 (
        .y(_T_359),
        .a(12'hF10),
        .b(_T_358)
    );
    wire [11:0] _T_362;
    BITWISEAND #(.width(12)) bitwiseand_173 (
        .y(_T_362),
        .a(csr_addr),
        .b(12'hFFF)
    );
    wire _T_363;
    wire [11:0] _WTEMP_15;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_174 (
        .y(_WTEMP_15),
        .in(10'h301)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_175 (
        .y(_T_363),
        .a(_WTEMP_15),
        .b(_T_362)
    );
    wire [11:0] _T_366;
    BITWISEAND #(.width(12)) bitwiseand_176 (
        .y(_T_366),
        .a(csr_addr),
        .b(12'hFFF)
    );
    wire _T_367;
    wire [11:0] _WTEMP_16;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_177 (
        .y(_WTEMP_16),
        .in(10'h302)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_178 (
        .y(_T_367),
        .a(_WTEMP_16),
        .b(_T_366)
    );
    wire [11:0] _T_370;
    BITWISEAND #(.width(12)) bitwiseand_179 (
        .y(_T_370),
        .a(csr_addr),
        .b(12'hFFF)
    );
    wire _T_371;
    wire [11:0] _WTEMP_17;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_180 (
        .y(_WTEMP_17),
        .in(10'h304)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_181 (
        .y(_T_371),
        .a(_WTEMP_17),
        .b(_T_370)
    );
    wire [11:0] _T_374;
    BITWISEAND #(.width(12)) bitwiseand_182 (
        .y(_T_374),
        .a(csr_addr),
        .b(12'hFFF)
    );
    wire _T_375;
    wire [11:0] _WTEMP_18;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_183 (
        .y(_WTEMP_18),
        .in(10'h321)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_184 (
        .y(_T_375),
        .a(_WTEMP_18),
        .b(_T_374)
    );
    wire [11:0] _T_378;
    BITWISEAND #(.width(12)) bitwiseand_185 (
        .y(_T_378),
        .a(csr_addr),
        .b(12'hFFF)
    );
    wire _T_379;
    wire [11:0] _WTEMP_19;
    PAD_UNSIGNED #(.width(11), .n(12)) u_pad_186 (
        .y(_WTEMP_19),
        .in(11'h701)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_187 (
        .y(_T_379),
        .a(_WTEMP_19),
        .b(_T_378)
    );
    wire [11:0] _T_382;
    BITWISEAND #(.width(12)) bitwiseand_188 (
        .y(_T_382),
        .a(csr_addr),
        .b(12'hFFF)
    );
    wire _T_383;
    wire [11:0] _WTEMP_20;
    PAD_UNSIGNED #(.width(11), .n(12)) u_pad_189 (
        .y(_WTEMP_20),
        .in(11'h741)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_190 (
        .y(_T_383),
        .a(_WTEMP_20),
        .b(_T_382)
    );
    wire [11:0] _T_386;
    BITWISEAND #(.width(12)) bitwiseand_191 (
        .y(_T_386),
        .a(csr_addr),
        .b(12'hFFF)
    );
    wire _T_387;
    wire [11:0] _WTEMP_21;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_192 (
        .y(_WTEMP_21),
        .in(10'h340)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_193 (
        .y(_T_387),
        .a(_WTEMP_21),
        .b(_T_386)
    );
    wire [11:0] _T_390;
    BITWISEAND #(.width(12)) bitwiseand_194 (
        .y(_T_390),
        .a(csr_addr),
        .b(12'hFFF)
    );
    wire _T_391;
    wire [11:0] _WTEMP_22;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_195 (
        .y(_WTEMP_22),
        .in(10'h341)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_196 (
        .y(_T_391),
        .a(_WTEMP_22),
        .b(_T_390)
    );
    wire [11:0] _T_394;
    BITWISEAND #(.width(12)) bitwiseand_197 (
        .y(_T_394),
        .a(csr_addr),
        .b(12'hFFF)
    );
    wire _T_395;
    wire [11:0] _WTEMP_23;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_198 (
        .y(_WTEMP_23),
        .in(10'h342)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_199 (
        .y(_T_395),
        .a(_WTEMP_23),
        .b(_T_394)
    );
    wire [11:0] _T_398;
    BITWISEAND #(.width(12)) bitwiseand_200 (
        .y(_T_398),
        .a(csr_addr),
        .b(12'hFFF)
    );
    wire _T_399;
    wire [11:0] _WTEMP_24;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_201 (
        .y(_WTEMP_24),
        .in(10'h343)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_202 (
        .y(_T_399),
        .a(_WTEMP_24),
        .b(_T_398)
    );
    wire [11:0] _T_402;
    BITWISEAND #(.width(12)) bitwiseand_203 (
        .y(_T_402),
        .a(csr_addr),
        .b(12'hFFF)
    );
    wire _T_403;
    wire [11:0] _WTEMP_25;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_204 (
        .y(_WTEMP_25),
        .in(10'h344)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_205 (
        .y(_T_403),
        .a(_WTEMP_25),
        .b(_T_402)
    );
    wire [11:0] _T_406;
    BITWISEAND #(.width(12)) bitwiseand_206 (
        .y(_T_406),
        .a(csr_addr),
        .b(12'hFFF)
    );
    wire _T_407;
    wire [11:0] _WTEMP_26;
    PAD_UNSIGNED #(.width(11), .n(12)) u_pad_207 (
        .y(_WTEMP_26),
        .in(11'h780)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_208 (
        .y(_T_407),
        .a(_WTEMP_26),
        .b(_T_406)
    );
    wire [11:0] _T_410;
    BITWISEAND #(.width(12)) bitwiseand_209 (
        .y(_T_410),
        .a(csr_addr),
        .b(12'hFFF)
    );
    wire _T_411;
    wire [11:0] _WTEMP_27;
    PAD_UNSIGNED #(.width(11), .n(12)) u_pad_210 (
        .y(_WTEMP_27),
        .in(11'h781)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_211 (
        .y(_T_411),
        .a(_WTEMP_27),
        .b(_T_410)
    );
    wire [11:0] _T_414;
    BITWISEAND #(.width(12)) bitwiseand_212 (
        .y(_T_414),
        .a(csr_addr),
        .b(12'hFFF)
    );
    wire _T_415;
    wire [11:0] _WTEMP_28;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_213 (
        .y(_WTEMP_28),
        .in(10'h300)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_214 (
        .y(_T_415),
        .a(_WTEMP_28),
        .b(_T_414)
    );
    wire _T_416;
    BITWISEOR #(.width(1)) bitwiseor_215 (
        .y(_T_416),
        .a(_T_303),
        .b(_T_307)
    );
    wire _T_417;
    BITWISEOR #(.width(1)) bitwiseor_216 (
        .y(_T_417),
        .a(_T_416),
        .b(_T_311)
    );
    wire _T_418;
    BITWISEOR #(.width(1)) bitwiseor_217 (
        .y(_T_418),
        .a(_T_417),
        .b(_T_315)
    );
    wire _T_419;
    BITWISEOR #(.width(1)) bitwiseor_218 (
        .y(_T_419),
        .a(_T_418),
        .b(_T_319)
    );
    wire _T_420;
    BITWISEOR #(.width(1)) bitwiseor_219 (
        .y(_T_420),
        .a(_T_419),
        .b(_T_323)
    );
    wire _T_421;
    BITWISEOR #(.width(1)) bitwiseor_220 (
        .y(_T_421),
        .a(_T_420),
        .b(_T_327)
    );
    wire _T_422;
    BITWISEOR #(.width(1)) bitwiseor_221 (
        .y(_T_422),
        .a(_T_421),
        .b(_T_331)
    );
    wire _T_423;
    BITWISEOR #(.width(1)) bitwiseor_222 (
        .y(_T_423),
        .a(_T_422),
        .b(_T_335)
    );
    wire _T_424;
    BITWISEOR #(.width(1)) bitwiseor_223 (
        .y(_T_424),
        .a(_T_423),
        .b(_T_339)
    );
    wire _T_425;
    BITWISEOR #(.width(1)) bitwiseor_224 (
        .y(_T_425),
        .a(_T_424),
        .b(_T_343)
    );
    wire _T_426;
    BITWISEOR #(.width(1)) bitwiseor_225 (
        .y(_T_426),
        .a(_T_425),
        .b(_T_347)
    );
    wire _T_427;
    BITWISEOR #(.width(1)) bitwiseor_226 (
        .y(_T_427),
        .a(_T_426),
        .b(_T_351)
    );
    wire _T_428;
    BITWISEOR #(.width(1)) bitwiseor_227 (
        .y(_T_428),
        .a(_T_427),
        .b(_T_355)
    );
    wire _T_429;
    BITWISEOR #(.width(1)) bitwiseor_228 (
        .y(_T_429),
        .a(_T_428),
        .b(_T_359)
    );
    wire _T_430;
    BITWISEOR #(.width(1)) bitwiseor_229 (
        .y(_T_430),
        .a(_T_429),
        .b(_T_363)
    );
    wire _T_431;
    BITWISEOR #(.width(1)) bitwiseor_230 (
        .y(_T_431),
        .a(_T_430),
        .b(_T_367)
    );
    wire _T_432;
    BITWISEOR #(.width(1)) bitwiseor_231 (
        .y(_T_432),
        .a(_T_431),
        .b(_T_371)
    );
    wire _T_433;
    BITWISEOR #(.width(1)) bitwiseor_232 (
        .y(_T_433),
        .a(_T_432),
        .b(_T_375)
    );
    wire _T_434;
    BITWISEOR #(.width(1)) bitwiseor_233 (
        .y(_T_434),
        .a(_T_433),
        .b(_T_379)
    );
    wire _T_435;
    BITWISEOR #(.width(1)) bitwiseor_234 (
        .y(_T_435),
        .a(_T_434),
        .b(_T_383)
    );
    wire _T_436;
    BITWISEOR #(.width(1)) bitwiseor_235 (
        .y(_T_436),
        .a(_T_435),
        .b(_T_387)
    );
    wire _T_437;
    BITWISEOR #(.width(1)) bitwiseor_236 (
        .y(_T_437),
        .a(_T_436),
        .b(_T_391)
    );
    wire _T_438;
    BITWISEOR #(.width(1)) bitwiseor_237 (
        .y(_T_438),
        .a(_T_437),
        .b(_T_395)
    );
    wire _T_439;
    BITWISEOR #(.width(1)) bitwiseor_238 (
        .y(_T_439),
        .a(_T_438),
        .b(_T_399)
    );
    wire _T_440;
    BITWISEOR #(.width(1)) bitwiseor_239 (
        .y(_T_440),
        .a(_T_439),
        .b(_T_403)
    );
    wire _T_441;
    BITWISEOR #(.width(1)) bitwiseor_240 (
        .y(_T_441),
        .a(_T_440),
        .b(_T_407)
    );
    wire _T_442;
    BITWISEOR #(.width(1)) bitwiseor_241 (
        .y(_T_442),
        .a(_T_441),
        .b(_T_411)
    );
    wire csrValid;
    BITWISEOR #(.width(1)) bitwiseor_242 (
        .y(csrValid),
        .a(_T_442),
        .b(_T_415)
    );
    wire [1:0] _T_443;
    BITS #(.width(12), .high(11), .low(10)) bits_243 (
        .y(_T_443),
        .in(csr_addr)
    );
    wire [1:0] _T_444;
    BITWISENOT #(.width(2)) bitwisenot_244 (
        .y(_T_444),
        .in(_T_443)
    );
    wire _T_446;
    wire [1:0] _WTEMP_29;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_245 (
        .y(_WTEMP_29),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(2)) u_eq_246 (
        .y(_T_446),
        .a(_T_444),
        .b(_WTEMP_29)
    );
    wire _T_447;
    EQ_UNSIGNED #(.width(12)) u_eq_247 (
        .y(_T_447),
        .a(csr_addr),
        .b(12'h301)
    );
    wire _T_448;
    BITWISEOR #(.width(1)) bitwiseor_248 (
        .y(_T_448),
        .a(_T_446),
        .b(_T_447)
    );
    wire _T_449;
    EQ_UNSIGNED #(.width(12)) u_eq_249 (
        .y(_T_449),
        .a(csr_addr),
        .b(12'h302)
    );
    wire csrRO;
    BITWISEOR #(.width(1)) bitwiseor_250 (
        .y(csrRO),
        .a(_T_448),
        .b(_T_449)
    );
    wire _T_450;
    EQ_UNSIGNED #(.width(3)) u_eq_251 (
        .y(_T_450),
        .a(io_cmd),
        .b(3'h1)
    );
    wire _T_451;
    BITS #(.width(3), .high(1), .low(1)) bits_252 (
        .y(_T_451),
        .in(io_cmd)
    );
    wire _T_453;
    wire [4:0] _WTEMP_30;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_253 (
        .y(_WTEMP_30),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(5)) u_neq_254 (
        .y(_T_453),
        .a(rs1_addr),
        .b(_WTEMP_30)
    );
    wire _T_454;
    BITWISEAND #(.width(1)) bitwiseand_255 (
        .y(_T_454),
        .a(_T_451),
        .b(_T_453)
    );
    wire wen;
    BITWISEOR #(.width(1)) bitwiseor_256 (
        .y(wen),
        .a(_T_450),
        .b(_T_454)
    );
    wire [31:0] _T_456;
    BITWISEOR #(.width(32)) bitwiseor_257 (
        .y(_T_456),
        .a(io_out),
        .b(io_in)
    );
    wire [31:0] _T_457;
    BITWISENOT #(.width(32)) bitwisenot_258 (
        .y(_T_457),
        .in(io_in)
    );
    wire [31:0] _T_458;
    BITWISEAND #(.width(32)) bitwiseand_259 (
        .y(_T_458),
        .a(io_out),
        .b(_T_457)
    );
    wire _T_459;
    EQ_UNSIGNED #(.width(3)) u_eq_260 (
        .y(_T_459),
        .a(3'h3),
        .b(io_cmd)
    );
    wire [31:0] _T_460;
    wire [31:0] _WTEMP_31;
    PAD_UNSIGNED #(.width(1), .n(32)) u_pad_261 (
        .y(_WTEMP_31),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(32)) u_mux_262 (
        .y(_T_460),
        .sel(_T_459),
        .a(_T_458),
        .b(_WTEMP_31)
    );
    wire _T_461;
    EQ_UNSIGNED #(.width(3)) u_eq_263 (
        .y(_T_461),
        .a(3'h2),
        .b(io_cmd)
    );
    wire [31:0] _T_462;
    MUX_UNSIGNED #(.width(32)) u_mux_264 (
        .y(_T_462),
        .sel(_T_461),
        .a(_T_456),
        .b(_T_460)
    );
    wire _T_463;
    EQ_UNSIGNED #(.width(3)) u_eq_265 (
        .y(_T_463),
        .a(3'h1),
        .b(io_cmd)
    );
    wire [31:0] wdata;
    MUX_UNSIGNED #(.width(32)) u_mux_266 (
        .y(wdata),
        .sel(_T_463),
        .a(io_in),
        .b(_T_462)
    );
    wire _T_464;
    BITS #(.width(32), .high(1), .low(1)) bits_267 (
        .y(_T_464),
        .in(io_addr)
    );
    wire iaddrInvalid;
    BITWISEAND #(.width(1)) bitwiseand_268 (
        .y(iaddrInvalid),
        .a(io_pc_check),
        .b(_T_464)
    );
    wire [1:0] _T_519;
    BITS #(.width(32), .high(1), .low(0)) bits_269 (
        .y(_T_519),
        .in(io_addr)
    );
    wire _T_521;
    wire [1:0] _WTEMP_32;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_270 (
        .y(_WTEMP_32),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(2)) u_neq_271 (
        .y(_T_521),
        .a(_T_519),
        .b(_WTEMP_32)
    );
    wire _T_522;
    BITS #(.width(32), .high(0), .low(0)) bits_272 (
        .y(_T_522),
        .in(io_addr)
    );
    wire _T_523;
    BITS #(.width(32), .high(0), .low(0)) bits_273 (
        .y(_T_523),
        .in(io_addr)
    );
    wire _T_524;
    EQ_UNSIGNED #(.width(3)) u_eq_274 (
        .y(_T_524),
        .a(3'h4),
        .b(io_ld_type)
    );
    wire _T_525;
    MUX_UNSIGNED #(.width(1)) u_mux_275 (
        .y(_T_525),
        .sel(_T_524),
        .a(_T_523),
        .b(1'h0)
    );
    wire _T_526;
    EQ_UNSIGNED #(.width(3)) u_eq_276 (
        .y(_T_526),
        .a(3'h2),
        .b(io_ld_type)
    );
    wire _T_527;
    MUX_UNSIGNED #(.width(1)) u_mux_277 (
        .y(_T_527),
        .sel(_T_526),
        .a(_T_522),
        .b(_T_525)
    );
    wire _T_528;
    EQ_UNSIGNED #(.width(3)) u_eq_278 (
        .y(_T_528),
        .a(3'h1),
        .b(io_ld_type)
    );
    wire laddrInvalid;
    MUX_UNSIGNED #(.width(1)) u_mux_279 (
        .y(laddrInvalid),
        .sel(_T_528),
        .a(_T_521),
        .b(_T_527)
    );
    wire [1:0] _T_530;
    BITS #(.width(32), .high(1), .low(0)) bits_280 (
        .y(_T_530),
        .in(io_addr)
    );
    wire _T_532;
    wire [1:0] _WTEMP_33;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_281 (
        .y(_WTEMP_33),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(2)) u_neq_282 (
        .y(_T_532),
        .a(_T_530),
        .b(_WTEMP_33)
    );
    wire _T_533;
    BITS #(.width(32), .high(0), .low(0)) bits_283 (
        .y(_T_533),
        .in(io_addr)
    );
    wire _T_534;
    EQ_UNSIGNED #(.width(2)) u_eq_284 (
        .y(_T_534),
        .a(2'h2),
        .b(io_st_type)
    );
    wire _T_535;
    MUX_UNSIGNED #(.width(1)) u_mux_285 (
        .y(_T_535),
        .sel(_T_534),
        .a(_T_533),
        .b(1'h0)
    );
    wire _T_536;
    EQ_UNSIGNED #(.width(2)) u_eq_286 (
        .y(_T_536),
        .a(2'h1),
        .b(io_st_type)
    );
    wire saddrInvalid;
    MUX_UNSIGNED #(.width(1)) u_mux_287 (
        .y(saddrInvalid),
        .sel(_T_536),
        .a(_T_532),
        .b(_T_535)
    );
    wire _T_537;
    BITWISEOR #(.width(1)) bitwiseor_288 (
        .y(_T_537),
        .a(io_illegal),
        .b(iaddrInvalid)
    );
    wire _T_538;
    BITWISEOR #(.width(1)) bitwiseor_289 (
        .y(_T_538),
        .a(_T_537),
        .b(laddrInvalid)
    );
    wire _T_539;
    BITWISEOR #(.width(1)) bitwiseor_290 (
        .y(_T_539),
        .a(_T_538),
        .b(saddrInvalid)
    );
    wire [1:0] _T_540;
    BITS #(.width(3), .high(1), .low(0)) bits_291 (
        .y(_T_540),
        .in(io_cmd)
    );
    wire _T_542;
    wire [1:0] _WTEMP_34;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_292 (
        .y(_WTEMP_34),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(2)) u_neq_293 (
        .y(_T_542),
        .a(_T_540),
        .b(_WTEMP_34)
    );
    wire _T_544;
    EQ_UNSIGNED #(.width(1)) u_eq_294 (
        .y(_T_544),
        .a(csrValid),
        .b(1'h0)
    );
    wire _T_546;
    EQ_UNSIGNED #(.width(1)) u_eq_295 (
        .y(_T_546),
        .a(privValid),
        .b(1'h0)
    );
    wire _T_547;
    BITWISEOR #(.width(1)) bitwiseor_296 (
        .y(_T_547),
        .a(_T_544),
        .b(_T_546)
    );
    wire _T_548;
    BITWISEAND #(.width(1)) bitwiseand_297 (
        .y(_T_548),
        .a(_T_542),
        .b(_T_547)
    );
    wire _T_549;
    BITWISEOR #(.width(1)) bitwiseor_298 (
        .y(_T_549),
        .a(_T_539),
        .b(_T_548)
    );
    wire _T_550;
    BITWISEAND #(.width(1)) bitwiseand_299 (
        .y(_T_550),
        .a(wen),
        .b(csrRO)
    );
    wire _T_551;
    BITWISEOR #(.width(1)) bitwiseor_300 (
        .y(_T_551),
        .a(_T_549),
        .b(_T_550)
    );
    wire _T_553;
    EQ_UNSIGNED #(.width(1)) u_eq_301 (
        .y(_T_553),
        .a(privValid),
        .b(1'h0)
    );
    wire _T_554;
    BITWISEAND #(.width(1)) bitwiseand_302 (
        .y(_T_554),
        .a(privInst),
        .b(_T_553)
    );
    wire _T_555;
    BITWISEOR #(.width(1)) bitwiseor_303 (
        .y(_T_555),
        .a(_T_551),
        .b(_T_554)
    );
    wire _T_556;
    BITWISEOR #(.width(1)) bitwiseor_304 (
        .y(_T_556),
        .a(_T_555),
        .b(isEcall)
    );
    wire _T_557;
    BITWISEOR #(.width(1)) bitwiseor_305 (
        .y(_T_557),
        .a(_T_556),
        .b(isEbreak)
    );
    wire [7:0] _T_558;
    SHL_UNSIGNED #(.width(2), .n(6)) u_shl_306 (
        .y(_T_558),
        .in(_PRV__q)
    );
    wire [32:0] _T_559;
    wire [31:0] _WTEMP_35;
    PAD_UNSIGNED #(.width(8), .n(32)) u_pad_307 (
        .y(_WTEMP_35),
        .in(_T_558)
    );
    ADD_UNSIGNED #(.width(32)) u_add_308 (
        .y(_T_559),
        .a(32'h100),
        .b(_WTEMP_35)
    );
    wire [31:0] _T_560;
    TAIL #(.width(33), .n(1)) tail_309 (
        .y(_T_560),
        .in(_T_559)
    );
    wire [32:0] _T_562;
    wire [31:0] _WTEMP_36;
    PAD_UNSIGNED #(.width(1), .n(32)) u_pad_310 (
        .y(_WTEMP_36),
        .in(1'h1)
    );
    ADD_UNSIGNED #(.width(32)) u_add_311 (
        .y(_T_562),
        .a(_time___q),
        .b(_WTEMP_36)
    );
    wire [31:0] _T_563;
    TAIL #(.width(33), .n(1)) tail_312 (
        .y(_T_563),
        .in(_T_562)
    );
    wire [31:0] _T_564;
    BITWISENOT #(.width(32)) bitwisenot_313 (
        .y(_T_564),
        .in(_time___q)
    );
    wire _T_566;
    wire [31:0] _WTEMP_37;
    PAD_UNSIGNED #(.width(1), .n(32)) u_pad_314 (
        .y(_WTEMP_37),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(32)) u_eq_315 (
        .y(_T_566),
        .a(_T_564),
        .b(_WTEMP_37)
    );
    wire [32:0] _T_568;
    wire [31:0] _WTEMP_38;
    PAD_UNSIGNED #(.width(1), .n(32)) u_pad_316 (
        .y(_WTEMP_38),
        .in(1'h1)
    );
    ADD_UNSIGNED #(.width(32)) u_add_317 (
        .y(_T_568),
        .a(_timeh__q),
        .b(_WTEMP_38)
    );
    wire [31:0] _T_569;
    TAIL #(.width(33), .n(1)) tail_318 (
        .y(_T_569),
        .in(_T_568)
    );
    wire [31:0] _GEN_1;
    MUX_UNSIGNED #(.width(32)) u_mux_319 (
        .y(_GEN_1),
        .sel(_T_566),
        .a(_T_569),
        .b(_timeh__q)
    );
    wire [32:0] _T_571;
    wire [31:0] _WTEMP_39;
    PAD_UNSIGNED #(.width(1), .n(32)) u_pad_320 (
        .y(_WTEMP_39),
        .in(1'h1)
    );
    ADD_UNSIGNED #(.width(32)) u_add_321 (
        .y(_T_571),
        .a(_cycle__q),
        .b(_WTEMP_39)
    );
    wire [31:0] _T_572;
    TAIL #(.width(33), .n(1)) tail_322 (
        .y(_T_572),
        .in(_T_571)
    );
    wire [31:0] _T_573;
    BITWISENOT #(.width(32)) bitwisenot_323 (
        .y(_T_573),
        .in(_cycle__q)
    );
    wire _T_575;
    wire [31:0] _WTEMP_40;
    PAD_UNSIGNED #(.width(1), .n(32)) u_pad_324 (
        .y(_WTEMP_40),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(32)) u_eq_325 (
        .y(_T_575),
        .a(_T_573),
        .b(_WTEMP_40)
    );
    wire [32:0] _T_577;
    wire [31:0] _WTEMP_41;
    PAD_UNSIGNED #(.width(1), .n(32)) u_pad_326 (
        .y(_WTEMP_41),
        .in(1'h1)
    );
    ADD_UNSIGNED #(.width(32)) u_add_327 (
        .y(_T_577),
        .a(_cycleh__q),
        .b(_WTEMP_41)
    );
    wire [31:0] _T_578;
    TAIL #(.width(33), .n(1)) tail_328 (
        .y(_T_578),
        .in(_T_577)
    );
    wire [31:0] _GEN_2;
    MUX_UNSIGNED #(.width(32)) u_mux_329 (
        .y(_GEN_2),
        .sel(_T_575),
        .a(_T_578),
        .b(_cycleh__q)
    );
    wire _T_580;
    NEQ_UNSIGNED #(.width(32)) u_neq_330 (
        .y(_T_580),
        .a(io_inst),
        .b(32'h13)
    );
    wire _T_582;
    EQ_UNSIGNED #(.width(1)) u_eq_331 (
        .y(_T_582),
        .a(io_expt),
        .b(1'h0)
    );
    wire _T_583;
    BITWISEOR #(.width(1)) bitwiseor_332 (
        .y(_T_583),
        .a(_T_582),
        .b(isEcall)
    );
    wire _T_584;
    BITWISEOR #(.width(1)) bitwiseor_333 (
        .y(_T_584),
        .a(_T_583),
        .b(isEbreak)
    );
    wire _T_585;
    BITWISEAND #(.width(1)) bitwiseand_334 (
        .y(_T_585),
        .a(_T_580),
        .b(_T_584)
    );
    wire _T_587;
    EQ_UNSIGNED #(.width(1)) u_eq_335 (
        .y(_T_587),
        .a(io_stall),
        .b(1'h0)
    );
    wire isInstRet;
    BITWISEAND #(.width(1)) bitwiseand_336 (
        .y(isInstRet),
        .a(_T_585),
        .b(_T_587)
    );
    wire [32:0] _T_589;
    wire [31:0] _WTEMP_42;
    PAD_UNSIGNED #(.width(1), .n(32)) u_pad_337 (
        .y(_WTEMP_42),
        .in(1'h1)
    );
    ADD_UNSIGNED #(.width(32)) u_add_338 (
        .y(_T_589),
        .a(_instret__q),
        .b(_WTEMP_42)
    );
    wire [31:0] _T_590;
    TAIL #(.width(33), .n(1)) tail_339 (
        .y(_T_590),
        .in(_T_589)
    );
    wire [31:0] _GEN_3;
    MUX_UNSIGNED #(.width(32)) u_mux_340 (
        .y(_GEN_3),
        .sel(isInstRet),
        .a(_T_590),
        .b(_instret__q)
    );
    wire [31:0] _T_591;
    BITWISENOT #(.width(32)) bitwisenot_341 (
        .y(_T_591),
        .in(_instret__q)
    );
    wire _T_593;
    wire [31:0] _WTEMP_43;
    PAD_UNSIGNED #(.width(1), .n(32)) u_pad_342 (
        .y(_WTEMP_43),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(32)) u_eq_343 (
        .y(_T_593),
        .a(_T_591),
        .b(_WTEMP_43)
    );
    wire _T_594;
    BITWISEAND #(.width(1)) bitwiseand_344 (
        .y(_T_594),
        .a(isInstRet),
        .b(_T_593)
    );
    wire [32:0] _T_596;
    wire [31:0] _WTEMP_44;
    PAD_UNSIGNED #(.width(1), .n(32)) u_pad_345 (
        .y(_WTEMP_44),
        .in(1'h1)
    );
    ADD_UNSIGNED #(.width(32)) u_add_346 (
        .y(_T_596),
        .a(_instreth__q),
        .b(_WTEMP_44)
    );
    wire [31:0] _T_597;
    TAIL #(.width(33), .n(1)) tail_347 (
        .y(_T_597),
        .in(_T_596)
    );
    wire [31:0] _GEN_4;
    MUX_UNSIGNED #(.width(32)) u_mux_348 (
        .y(_GEN_4),
        .sel(_T_594),
        .a(_T_597),
        .b(_instreth__q)
    );
    wire _T_599;
    EQ_UNSIGNED #(.width(1)) u_eq_349 (
        .y(_T_599),
        .a(io_stall),
        .b(1'h0)
    );
    wire [29:0] _T_600;
    SHR_UNSIGNED #(.width(32), .n(2)) u_shr_350 (
        .y(_T_600),
        .in(io_pc)
    );
    wire [31:0] _T_601;
    SHL_UNSIGNED #(.width(30), .n(2)) u_shl_351 (
        .y(_T_601),
        .in(_T_600)
    );
    wire [4:0] _T_608;
    wire [3:0] _WTEMP_45;
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_352 (
        .y(_WTEMP_45),
        .in(_PRV__q)
    );
    ADD_UNSIGNED #(.width(4)) u_add_353 (
        .y(_T_608),
        .a(4'h8),
        .b(_WTEMP_45)
    );
    wire [3:0] _T_609;
    TAIL #(.width(5), .n(1)) tail_354 (
        .y(_T_609),
        .in(_T_608)
    );
    wire [1:0] _T_610;
    MUX_UNSIGNED #(.width(2)) u_mux_355 (
        .y(_T_610),
        .sel(isEbreak),
        .a(2'h3),
        .b(2'h2)
    );
    wire [3:0] _T_611;
    wire [3:0] _WTEMP_46;
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_356 (
        .y(_WTEMP_46),
        .in(_T_610)
    );
    MUX_UNSIGNED #(.width(4)) u_mux_357 (
        .y(_T_611),
        .sel(isEcall),
        .a(_T_609),
        .b(_WTEMP_46)
    );
    wire [3:0] _T_612;
    wire [3:0] _WTEMP_47;
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_358 (
        .y(_WTEMP_47),
        .in(3'h6)
    );
    MUX_UNSIGNED #(.width(4)) u_mux_359 (
        .y(_T_612),
        .sel(saddrInvalid),
        .a(_WTEMP_47),
        .b(_T_611)
    );
    wire [3:0] _T_613;
    wire [3:0] _WTEMP_48;
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_360 (
        .y(_WTEMP_48),
        .in(3'h4)
    );
    MUX_UNSIGNED #(.width(4)) u_mux_361 (
        .y(_T_613),
        .sel(laddrInvalid),
        .a(_WTEMP_48),
        .b(_T_612)
    );
    wire [3:0] _T_614;
    wire [3:0] _WTEMP_49;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_362 (
        .y(_WTEMP_49),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(4)) u_mux_363 (
        .y(_T_614),
        .sel(iaddrInvalid),
        .a(_WTEMP_49),
        .b(_T_613)
    );
    wire _T_616;
    BITWISEOR #(.width(1)) bitwiseor_364 (
        .y(_T_616),
        .a(iaddrInvalid),
        .b(laddrInvalid)
    );
    wire _T_617;
    BITWISEOR #(.width(1)) bitwiseor_365 (
        .y(_T_617),
        .a(_T_616),
        .b(saddrInvalid)
    );
    wire [31:0] _GEN_5;
    MUX_UNSIGNED #(.width(32)) u_mux_366 (
        .y(_GEN_5),
        .sel(_T_617),
        .a(io_addr),
        .b(_mbadaddr__q)
    );
    wire [31:0] _GEN_6;
    MUX_UNSIGNED #(.width(32)) u_mux_367 (
        .y(_GEN_6),
        .sel(io_expt),
        .a(_T_601),
        .b(_mepc__q)
    );
    wire [31:0] _GEN_7;
    wire [31:0] _WTEMP_50;
    PAD_UNSIGNED #(.width(4), .n(32)) u_pad_368 (
        .y(_WTEMP_50),
        .in(_T_614)
    );
    MUX_UNSIGNED #(.width(32)) u_mux_369 (
        .y(_GEN_7),
        .sel(io_expt),
        .a(_WTEMP_50),
        .b(_mcause__q)
    );
    wire [1:0] _GEN_8;
    MUX_UNSIGNED #(.width(2)) u_mux_370 (
        .y(_GEN_8),
        .sel(io_expt),
        .a(2'h3),
        .b(_PRV__q)
    );
    wire _GEN_9;
    MUX_UNSIGNED #(.width(1)) u_mux_371 (
        .y(_GEN_9),
        .sel(io_expt),
        .a(1'h0),
        .b(_IE__q)
    );
    wire [1:0] _GEN_10;
    MUX_UNSIGNED #(.width(2)) u_mux_372 (
        .y(_GEN_10),
        .sel(io_expt),
        .a(_PRV__q),
        .b(_PRV1__q)
    );
    wire _GEN_11;
    MUX_UNSIGNED #(.width(1)) u_mux_373 (
        .y(_GEN_11),
        .sel(io_expt),
        .a(_IE__q),
        .b(_IE1__q)
    );
    wire [31:0] _GEN_12;
    MUX_UNSIGNED #(.width(32)) u_mux_374 (
        .y(_GEN_12),
        .sel(io_expt),
        .a(_GEN_5),
        .b(_mbadaddr__q)
    );
    wire _T_619;
    EQ_UNSIGNED #(.width(1)) u_eq_375 (
        .y(_T_619),
        .a(io_expt),
        .b(1'h0)
    );
    wire _T_620;
    BITWISEAND #(.width(1)) bitwiseand_376 (
        .y(_T_620),
        .a(_T_619),
        .b(isEret)
    );
    wire [1:0] _GEN_13;
    MUX_UNSIGNED #(.width(2)) u_mux_377 (
        .y(_GEN_13),
        .sel(_T_620),
        .a(_PRV1__q),
        .b(_GEN_8)
    );
    wire _GEN_14;
    MUX_UNSIGNED #(.width(1)) u_mux_378 (
        .y(_GEN_14),
        .sel(_T_620),
        .a(_IE1__q),
        .b(_GEN_9)
    );
    wire [1:0] _GEN_15;
    MUX_UNSIGNED #(.width(2)) u_mux_379 (
        .y(_GEN_15),
        .sel(_T_620),
        .a(2'h0),
        .b(_GEN_10)
    );
    wire _GEN_16;
    MUX_UNSIGNED #(.width(1)) u_mux_380 (
        .y(_GEN_16),
        .sel(_T_620),
        .a(1'h1),
        .b(_GEN_11)
    );
    wire _T_623;
    EQ_UNSIGNED #(.width(1)) u_eq_381 (
        .y(_T_623),
        .a(io_expt),
        .b(1'h0)
    );
    wire _T_625;
    EQ_UNSIGNED #(.width(1)) u_eq_382 (
        .y(_T_625),
        .a(isEret),
        .b(1'h0)
    );
    wire _T_626;
    BITWISEAND #(.width(1)) bitwiseand_383 (
        .y(_T_626),
        .a(_T_623),
        .b(_T_625)
    );
    wire _T_627;
    BITWISEAND #(.width(1)) bitwiseand_384 (
        .y(_T_627),
        .a(_T_626),
        .b(wen)
    );
    wire _T_628;
    EQ_UNSIGNED #(.width(12)) u_eq_385 (
        .y(_T_628),
        .a(csr_addr),
        .b(12'h300)
    );
    wire [1:0] _T_629;
    BITS #(.width(32), .high(5), .low(4)) bits_386 (
        .y(_T_629),
        .in(wdata)
    );
    wire _T_630;
    BITS #(.width(32), .high(3), .low(3)) bits_387 (
        .y(_T_630),
        .in(wdata)
    );
    wire [1:0] _T_631;
    BITS #(.width(32), .high(2), .low(1)) bits_388 (
        .y(_T_631),
        .in(wdata)
    );
    wire _T_632;
    BITS #(.width(32), .high(0), .low(0)) bits_389 (
        .y(_T_632),
        .in(wdata)
    );
    wire [1:0] _GEN_17;
    MUX_UNSIGNED #(.width(2)) u_mux_390 (
        .y(_GEN_17),
        .sel(_T_628),
        .a(_T_629),
        .b(_GEN_15)
    );
    wire _GEN_18;
    MUX_UNSIGNED #(.width(1)) u_mux_391 (
        .y(_GEN_18),
        .sel(_T_628),
        .a(_T_630),
        .b(_GEN_16)
    );
    wire [1:0] _GEN_19;
    MUX_UNSIGNED #(.width(2)) u_mux_392 (
        .y(_GEN_19),
        .sel(_T_628),
        .a(_T_631),
        .b(_GEN_13)
    );
    wire _GEN_20;
    MUX_UNSIGNED #(.width(1)) u_mux_393 (
        .y(_GEN_20),
        .sel(_T_628),
        .a(_T_632),
        .b(_GEN_14)
    );
    wire _T_633;
    EQ_UNSIGNED #(.width(12)) u_eq_394 (
        .y(_T_633),
        .a(csr_addr),
        .b(12'h344)
    );
    wire _T_635;
    EQ_UNSIGNED #(.width(1)) u_eq_395 (
        .y(_T_635),
        .a(_T_628),
        .b(1'h0)
    );
    wire _T_636;
    BITWISEAND #(.width(1)) bitwiseand_396 (
        .y(_T_636),
        .a(_T_635),
        .b(_T_633)
    );
    wire _T_637;
    BITS #(.width(32), .high(7), .low(7)) bits_397 (
        .y(_T_637),
        .in(wdata)
    );
    wire _T_638;
    BITS #(.width(32), .high(3), .low(3)) bits_398 (
        .y(_T_638),
        .in(wdata)
    );
    wire _GEN_21;
    MUX_UNSIGNED #(.width(1)) u_mux_399 (
        .y(_GEN_21),
        .sel(_T_636),
        .a(_T_637),
        .b(_MTIP__q)
    );
    wire _GEN_22;
    MUX_UNSIGNED #(.width(1)) u_mux_400 (
        .y(_GEN_22),
        .sel(_T_636),
        .a(_T_638),
        .b(_MSIP__q)
    );
    wire _T_639;
    EQ_UNSIGNED #(.width(12)) u_eq_401 (
        .y(_T_639),
        .a(csr_addr),
        .b(12'h304)
    );
    wire _T_641;
    EQ_UNSIGNED #(.width(1)) u_eq_402 (
        .y(_T_641),
        .a(_T_628),
        .b(1'h0)
    );
    wire _T_643;
    EQ_UNSIGNED #(.width(1)) u_eq_403 (
        .y(_T_643),
        .a(_T_633),
        .b(1'h0)
    );
    wire _T_644;
    BITWISEAND #(.width(1)) bitwiseand_404 (
        .y(_T_644),
        .a(_T_641),
        .b(_T_643)
    );
    wire _T_645;
    BITWISEAND #(.width(1)) bitwiseand_405 (
        .y(_T_645),
        .a(_T_644),
        .b(_T_639)
    );
    wire _T_646;
    BITS #(.width(32), .high(7), .low(7)) bits_406 (
        .y(_T_646),
        .in(wdata)
    );
    wire _T_647;
    BITS #(.width(32), .high(3), .low(3)) bits_407 (
        .y(_T_647),
        .in(wdata)
    );
    wire _GEN_23;
    MUX_UNSIGNED #(.width(1)) u_mux_408 (
        .y(_GEN_23),
        .sel(_T_645),
        .a(_T_646),
        .b(_MTIE__q)
    );
    wire _GEN_24;
    MUX_UNSIGNED #(.width(1)) u_mux_409 (
        .y(_GEN_24),
        .sel(_T_645),
        .a(_T_647),
        .b(_MSIE__q)
    );
    wire _T_648;
    EQ_UNSIGNED #(.width(12)) u_eq_410 (
        .y(_T_648),
        .a(csr_addr),
        .b(12'h701)
    );
    wire _T_650;
    EQ_UNSIGNED #(.width(1)) u_eq_411 (
        .y(_T_650),
        .a(_T_628),
        .b(1'h0)
    );
    wire _T_652;
    EQ_UNSIGNED #(.width(1)) u_eq_412 (
        .y(_T_652),
        .a(_T_633),
        .b(1'h0)
    );
    wire _T_653;
    BITWISEAND #(.width(1)) bitwiseand_413 (
        .y(_T_653),
        .a(_T_650),
        .b(_T_652)
    );
    wire _T_655;
    EQ_UNSIGNED #(.width(1)) u_eq_414 (
        .y(_T_655),
        .a(_T_639),
        .b(1'h0)
    );
    wire _T_656;
    BITWISEAND #(.width(1)) bitwiseand_415 (
        .y(_T_656),
        .a(_T_653),
        .b(_T_655)
    );
    wire _T_657;
    BITWISEAND #(.width(1)) bitwiseand_416 (
        .y(_T_657),
        .a(_T_656),
        .b(_T_648)
    );
    wire [31:0] _GEN_25;
    MUX_UNSIGNED #(.width(32)) u_mux_417 (
        .y(_GEN_25),
        .sel(_T_657),
        .a(wdata),
        .b(_T_563)
    );
    wire _T_658;
    EQ_UNSIGNED #(.width(12)) u_eq_418 (
        .y(_T_658),
        .a(csr_addr),
        .b(12'h741)
    );
    wire _T_660;
    EQ_UNSIGNED #(.width(1)) u_eq_419 (
        .y(_T_660),
        .a(_T_628),
        .b(1'h0)
    );
    wire _T_662;
    EQ_UNSIGNED #(.width(1)) u_eq_420 (
        .y(_T_662),
        .a(_T_633),
        .b(1'h0)
    );
    wire _T_663;
    BITWISEAND #(.width(1)) bitwiseand_421 (
        .y(_T_663),
        .a(_T_660),
        .b(_T_662)
    );
    wire _T_665;
    EQ_UNSIGNED #(.width(1)) u_eq_422 (
        .y(_T_665),
        .a(_T_639),
        .b(1'h0)
    );
    wire _T_666;
    BITWISEAND #(.width(1)) bitwiseand_423 (
        .y(_T_666),
        .a(_T_663),
        .b(_T_665)
    );
    wire _T_668;
    EQ_UNSIGNED #(.width(1)) u_eq_424 (
        .y(_T_668),
        .a(_T_648),
        .b(1'h0)
    );
    wire _T_669;
    BITWISEAND #(.width(1)) bitwiseand_425 (
        .y(_T_669),
        .a(_T_666),
        .b(_T_668)
    );
    wire _T_670;
    BITWISEAND #(.width(1)) bitwiseand_426 (
        .y(_T_670),
        .a(_T_669),
        .b(_T_658)
    );
    wire [31:0] _GEN_26;
    MUX_UNSIGNED #(.width(32)) u_mux_427 (
        .y(_GEN_26),
        .sel(_T_670),
        .a(wdata),
        .b(_GEN_1)
    );
    wire _T_671;
    EQ_UNSIGNED #(.width(12)) u_eq_428 (
        .y(_T_671),
        .a(csr_addr),
        .b(12'h321)
    );
    wire _T_673;
    EQ_UNSIGNED #(.width(1)) u_eq_429 (
        .y(_T_673),
        .a(_T_628),
        .b(1'h0)
    );
    wire _T_675;
    EQ_UNSIGNED #(.width(1)) u_eq_430 (
        .y(_T_675),
        .a(_T_633),
        .b(1'h0)
    );
    wire _T_676;
    BITWISEAND #(.width(1)) bitwiseand_431 (
        .y(_T_676),
        .a(_T_673),
        .b(_T_675)
    );
    wire _T_678;
    EQ_UNSIGNED #(.width(1)) u_eq_432 (
        .y(_T_678),
        .a(_T_639),
        .b(1'h0)
    );
    wire _T_679;
    BITWISEAND #(.width(1)) bitwiseand_433 (
        .y(_T_679),
        .a(_T_676),
        .b(_T_678)
    );
    wire _T_681;
    EQ_UNSIGNED #(.width(1)) u_eq_434 (
        .y(_T_681),
        .a(_T_648),
        .b(1'h0)
    );
    wire _T_682;
    BITWISEAND #(.width(1)) bitwiseand_435 (
        .y(_T_682),
        .a(_T_679),
        .b(_T_681)
    );
    wire _T_684;
    EQ_UNSIGNED #(.width(1)) u_eq_436 (
        .y(_T_684),
        .a(_T_658),
        .b(1'h0)
    );
    wire _T_685;
    BITWISEAND #(.width(1)) bitwiseand_437 (
        .y(_T_685),
        .a(_T_682),
        .b(_T_684)
    );
    wire _T_686;
    BITWISEAND #(.width(1)) bitwiseand_438 (
        .y(_T_686),
        .a(_T_685),
        .b(_T_671)
    );
    wire [31:0] _GEN_27;
    MUX_UNSIGNED #(.width(32)) u_mux_439 (
        .y(_GEN_27),
        .sel(_T_686),
        .a(wdata),
        .b(_mtimecmp__q)
    );
    wire _T_687;
    EQ_UNSIGNED #(.width(12)) u_eq_440 (
        .y(_T_687),
        .a(csr_addr),
        .b(12'h340)
    );
    wire _T_689;
    EQ_UNSIGNED #(.width(1)) u_eq_441 (
        .y(_T_689),
        .a(_T_628),
        .b(1'h0)
    );
    wire _T_691;
    EQ_UNSIGNED #(.width(1)) u_eq_442 (
        .y(_T_691),
        .a(_T_633),
        .b(1'h0)
    );
    wire _T_692;
    BITWISEAND #(.width(1)) bitwiseand_443 (
        .y(_T_692),
        .a(_T_689),
        .b(_T_691)
    );
    wire _T_694;
    EQ_UNSIGNED #(.width(1)) u_eq_444 (
        .y(_T_694),
        .a(_T_639),
        .b(1'h0)
    );
    wire _T_695;
    BITWISEAND #(.width(1)) bitwiseand_445 (
        .y(_T_695),
        .a(_T_692),
        .b(_T_694)
    );
    wire _T_697;
    EQ_UNSIGNED #(.width(1)) u_eq_446 (
        .y(_T_697),
        .a(_T_648),
        .b(1'h0)
    );
    wire _T_698;
    BITWISEAND #(.width(1)) bitwiseand_447 (
        .y(_T_698),
        .a(_T_695),
        .b(_T_697)
    );
    wire _T_700;
    EQ_UNSIGNED #(.width(1)) u_eq_448 (
        .y(_T_700),
        .a(_T_658),
        .b(1'h0)
    );
    wire _T_701;
    BITWISEAND #(.width(1)) bitwiseand_449 (
        .y(_T_701),
        .a(_T_698),
        .b(_T_700)
    );
    wire _T_703;
    EQ_UNSIGNED #(.width(1)) u_eq_450 (
        .y(_T_703),
        .a(_T_671),
        .b(1'h0)
    );
    wire _T_704;
    BITWISEAND #(.width(1)) bitwiseand_451 (
        .y(_T_704),
        .a(_T_701),
        .b(_T_703)
    );
    wire _T_705;
    BITWISEAND #(.width(1)) bitwiseand_452 (
        .y(_T_705),
        .a(_T_704),
        .b(_T_687)
    );
    wire [31:0] _GEN_28;
    MUX_UNSIGNED #(.width(32)) u_mux_453 (
        .y(_GEN_28),
        .sel(_T_705),
        .a(wdata),
        .b(_mscratch__q)
    );
    wire _T_706;
    EQ_UNSIGNED #(.width(12)) u_eq_454 (
        .y(_T_706),
        .a(csr_addr),
        .b(12'h341)
    );
    wire _T_708;
    EQ_UNSIGNED #(.width(1)) u_eq_455 (
        .y(_T_708),
        .a(_T_628),
        .b(1'h0)
    );
    wire _T_710;
    EQ_UNSIGNED #(.width(1)) u_eq_456 (
        .y(_T_710),
        .a(_T_633),
        .b(1'h0)
    );
    wire _T_711;
    BITWISEAND #(.width(1)) bitwiseand_457 (
        .y(_T_711),
        .a(_T_708),
        .b(_T_710)
    );
    wire _T_713;
    EQ_UNSIGNED #(.width(1)) u_eq_458 (
        .y(_T_713),
        .a(_T_639),
        .b(1'h0)
    );
    wire _T_714;
    BITWISEAND #(.width(1)) bitwiseand_459 (
        .y(_T_714),
        .a(_T_711),
        .b(_T_713)
    );
    wire _T_716;
    EQ_UNSIGNED #(.width(1)) u_eq_460 (
        .y(_T_716),
        .a(_T_648),
        .b(1'h0)
    );
    wire _T_717;
    BITWISEAND #(.width(1)) bitwiseand_461 (
        .y(_T_717),
        .a(_T_714),
        .b(_T_716)
    );
    wire _T_719;
    EQ_UNSIGNED #(.width(1)) u_eq_462 (
        .y(_T_719),
        .a(_T_658),
        .b(1'h0)
    );
    wire _T_720;
    BITWISEAND #(.width(1)) bitwiseand_463 (
        .y(_T_720),
        .a(_T_717),
        .b(_T_719)
    );
    wire _T_722;
    EQ_UNSIGNED #(.width(1)) u_eq_464 (
        .y(_T_722),
        .a(_T_671),
        .b(1'h0)
    );
    wire _T_723;
    BITWISEAND #(.width(1)) bitwiseand_465 (
        .y(_T_723),
        .a(_T_720),
        .b(_T_722)
    );
    wire _T_725;
    EQ_UNSIGNED #(.width(1)) u_eq_466 (
        .y(_T_725),
        .a(_T_687),
        .b(1'h0)
    );
    wire _T_726;
    BITWISEAND #(.width(1)) bitwiseand_467 (
        .y(_T_726),
        .a(_T_723),
        .b(_T_725)
    );
    wire _T_727;
    BITWISEAND #(.width(1)) bitwiseand_468 (
        .y(_T_727),
        .a(_T_726),
        .b(_T_706)
    );
    wire [31:0] _T_729;
    DSHR_UNSIGNED #(.width_in(32), .width_n(2)) u_dshr_469 (
        .y(_T_729),
        .in(wdata),
        .n(2'h2)
    );
    wire [34:0] _T_731;
    DSHL_UNSIGNED #(.width_in(32), .width_n(2)) u_dshl_470 (
        .y(_T_731),
        .in(_T_729),
        .n(2'h2)
    );
    wire [34:0] _GEN_29;
    wire [34:0] _WTEMP_51;
    PAD_UNSIGNED #(.width(32), .n(35)) u_pad_471 (
        .y(_WTEMP_51),
        .in(_GEN_6)
    );
    MUX_UNSIGNED #(.width(35)) u_mux_472 (
        .y(_GEN_29),
        .sel(_T_727),
        .a(_T_731),
        .b(_WTEMP_51)
    );
    wire _T_732;
    EQ_UNSIGNED #(.width(12)) u_eq_473 (
        .y(_T_732),
        .a(csr_addr),
        .b(12'h342)
    );
    wire _T_734;
    EQ_UNSIGNED #(.width(1)) u_eq_474 (
        .y(_T_734),
        .a(_T_628),
        .b(1'h0)
    );
    wire _T_736;
    EQ_UNSIGNED #(.width(1)) u_eq_475 (
        .y(_T_736),
        .a(_T_633),
        .b(1'h0)
    );
    wire _T_737;
    BITWISEAND #(.width(1)) bitwiseand_476 (
        .y(_T_737),
        .a(_T_734),
        .b(_T_736)
    );
    wire _T_739;
    EQ_UNSIGNED #(.width(1)) u_eq_477 (
        .y(_T_739),
        .a(_T_639),
        .b(1'h0)
    );
    wire _T_740;
    BITWISEAND #(.width(1)) bitwiseand_478 (
        .y(_T_740),
        .a(_T_737),
        .b(_T_739)
    );
    wire _T_742;
    EQ_UNSIGNED #(.width(1)) u_eq_479 (
        .y(_T_742),
        .a(_T_648),
        .b(1'h0)
    );
    wire _T_743;
    BITWISEAND #(.width(1)) bitwiseand_480 (
        .y(_T_743),
        .a(_T_740),
        .b(_T_742)
    );
    wire _T_745;
    EQ_UNSIGNED #(.width(1)) u_eq_481 (
        .y(_T_745),
        .a(_T_658),
        .b(1'h0)
    );
    wire _T_746;
    BITWISEAND #(.width(1)) bitwiseand_482 (
        .y(_T_746),
        .a(_T_743),
        .b(_T_745)
    );
    wire _T_748;
    EQ_UNSIGNED #(.width(1)) u_eq_483 (
        .y(_T_748),
        .a(_T_671),
        .b(1'h0)
    );
    wire _T_749;
    BITWISEAND #(.width(1)) bitwiseand_484 (
        .y(_T_749),
        .a(_T_746),
        .b(_T_748)
    );
    wire _T_751;
    EQ_UNSIGNED #(.width(1)) u_eq_485 (
        .y(_T_751),
        .a(_T_687),
        .b(1'h0)
    );
    wire _T_752;
    BITWISEAND #(.width(1)) bitwiseand_486 (
        .y(_T_752),
        .a(_T_749),
        .b(_T_751)
    );
    wire _T_754;
    EQ_UNSIGNED #(.width(1)) u_eq_487 (
        .y(_T_754),
        .a(_T_706),
        .b(1'h0)
    );
    wire _T_755;
    BITWISEAND #(.width(1)) bitwiseand_488 (
        .y(_T_755),
        .a(_T_752),
        .b(_T_754)
    );
    wire _T_756;
    BITWISEAND #(.width(1)) bitwiseand_489 (
        .y(_T_756),
        .a(_T_755),
        .b(_T_732)
    );
    wire [31:0] _T_758;
    BITWISEAND #(.width(32)) bitwiseand_490 (
        .y(_T_758),
        .a(wdata),
        .b(32'h8000000F)
    );
    wire [31:0] _GEN_30;
    MUX_UNSIGNED #(.width(32)) u_mux_491 (
        .y(_GEN_30),
        .sel(_T_756),
        .a(_T_758),
        .b(_GEN_7)
    );
    wire _T_759;
    EQ_UNSIGNED #(.width(12)) u_eq_492 (
        .y(_T_759),
        .a(csr_addr),
        .b(12'h343)
    );
    wire _T_761;
    EQ_UNSIGNED #(.width(1)) u_eq_493 (
        .y(_T_761),
        .a(_T_628),
        .b(1'h0)
    );
    wire _T_763;
    EQ_UNSIGNED #(.width(1)) u_eq_494 (
        .y(_T_763),
        .a(_T_633),
        .b(1'h0)
    );
    wire _T_764;
    BITWISEAND #(.width(1)) bitwiseand_495 (
        .y(_T_764),
        .a(_T_761),
        .b(_T_763)
    );
    wire _T_766;
    EQ_UNSIGNED #(.width(1)) u_eq_496 (
        .y(_T_766),
        .a(_T_639),
        .b(1'h0)
    );
    wire _T_767;
    BITWISEAND #(.width(1)) bitwiseand_497 (
        .y(_T_767),
        .a(_T_764),
        .b(_T_766)
    );
    wire _T_769;
    EQ_UNSIGNED #(.width(1)) u_eq_498 (
        .y(_T_769),
        .a(_T_648),
        .b(1'h0)
    );
    wire _T_770;
    BITWISEAND #(.width(1)) bitwiseand_499 (
        .y(_T_770),
        .a(_T_767),
        .b(_T_769)
    );
    wire _T_772;
    EQ_UNSIGNED #(.width(1)) u_eq_500 (
        .y(_T_772),
        .a(_T_658),
        .b(1'h0)
    );
    wire _T_773;
    BITWISEAND #(.width(1)) bitwiseand_501 (
        .y(_T_773),
        .a(_T_770),
        .b(_T_772)
    );
    wire _T_775;
    EQ_UNSIGNED #(.width(1)) u_eq_502 (
        .y(_T_775),
        .a(_T_671),
        .b(1'h0)
    );
    wire _T_776;
    BITWISEAND #(.width(1)) bitwiseand_503 (
        .y(_T_776),
        .a(_T_773),
        .b(_T_775)
    );
    wire _T_778;
    EQ_UNSIGNED #(.width(1)) u_eq_504 (
        .y(_T_778),
        .a(_T_687),
        .b(1'h0)
    );
    wire _T_779;
    BITWISEAND #(.width(1)) bitwiseand_505 (
        .y(_T_779),
        .a(_T_776),
        .b(_T_778)
    );
    wire _T_781;
    EQ_UNSIGNED #(.width(1)) u_eq_506 (
        .y(_T_781),
        .a(_T_706),
        .b(1'h0)
    );
    wire _T_782;
    BITWISEAND #(.width(1)) bitwiseand_507 (
        .y(_T_782),
        .a(_T_779),
        .b(_T_781)
    );
    wire _T_784;
    EQ_UNSIGNED #(.width(1)) u_eq_508 (
        .y(_T_784),
        .a(_T_732),
        .b(1'h0)
    );
    wire _T_785;
    BITWISEAND #(.width(1)) bitwiseand_509 (
        .y(_T_785),
        .a(_T_782),
        .b(_T_784)
    );
    wire _T_786;
    BITWISEAND #(.width(1)) bitwiseand_510 (
        .y(_T_786),
        .a(_T_785),
        .b(_T_759)
    );
    wire [31:0] _GEN_31;
    MUX_UNSIGNED #(.width(32)) u_mux_511 (
        .y(_GEN_31),
        .sel(_T_786),
        .a(wdata),
        .b(_GEN_12)
    );
    wire _T_787;
    EQ_UNSIGNED #(.width(12)) u_eq_512 (
        .y(_T_787),
        .a(csr_addr),
        .b(12'h780)
    );
    wire _T_789;
    EQ_UNSIGNED #(.width(1)) u_eq_513 (
        .y(_T_789),
        .a(_T_628),
        .b(1'h0)
    );
    wire _T_791;
    EQ_UNSIGNED #(.width(1)) u_eq_514 (
        .y(_T_791),
        .a(_T_633),
        .b(1'h0)
    );
    wire _T_792;
    BITWISEAND #(.width(1)) bitwiseand_515 (
        .y(_T_792),
        .a(_T_789),
        .b(_T_791)
    );
    wire _T_794;
    EQ_UNSIGNED #(.width(1)) u_eq_516 (
        .y(_T_794),
        .a(_T_639),
        .b(1'h0)
    );
    wire _T_795;
    BITWISEAND #(.width(1)) bitwiseand_517 (
        .y(_T_795),
        .a(_T_792),
        .b(_T_794)
    );
    wire _T_797;
    EQ_UNSIGNED #(.width(1)) u_eq_518 (
        .y(_T_797),
        .a(_T_648),
        .b(1'h0)
    );
    wire _T_798;
    BITWISEAND #(.width(1)) bitwiseand_519 (
        .y(_T_798),
        .a(_T_795),
        .b(_T_797)
    );
    wire _T_800;
    EQ_UNSIGNED #(.width(1)) u_eq_520 (
        .y(_T_800),
        .a(_T_658),
        .b(1'h0)
    );
    wire _T_801;
    BITWISEAND #(.width(1)) bitwiseand_521 (
        .y(_T_801),
        .a(_T_798),
        .b(_T_800)
    );
    wire _T_803;
    EQ_UNSIGNED #(.width(1)) u_eq_522 (
        .y(_T_803),
        .a(_T_671),
        .b(1'h0)
    );
    wire _T_804;
    BITWISEAND #(.width(1)) bitwiseand_523 (
        .y(_T_804),
        .a(_T_801),
        .b(_T_803)
    );
    wire _T_806;
    EQ_UNSIGNED #(.width(1)) u_eq_524 (
        .y(_T_806),
        .a(_T_687),
        .b(1'h0)
    );
    wire _T_807;
    BITWISEAND #(.width(1)) bitwiseand_525 (
        .y(_T_807),
        .a(_T_804),
        .b(_T_806)
    );
    wire _T_809;
    EQ_UNSIGNED #(.width(1)) u_eq_526 (
        .y(_T_809),
        .a(_T_706),
        .b(1'h0)
    );
    wire _T_810;
    BITWISEAND #(.width(1)) bitwiseand_527 (
        .y(_T_810),
        .a(_T_807),
        .b(_T_809)
    );
    wire _T_812;
    EQ_UNSIGNED #(.width(1)) u_eq_528 (
        .y(_T_812),
        .a(_T_732),
        .b(1'h0)
    );
    wire _T_813;
    BITWISEAND #(.width(1)) bitwiseand_529 (
        .y(_T_813),
        .a(_T_810),
        .b(_T_812)
    );
    wire _T_815;
    EQ_UNSIGNED #(.width(1)) u_eq_530 (
        .y(_T_815),
        .a(_T_759),
        .b(1'h0)
    );
    wire _T_816;
    BITWISEAND #(.width(1)) bitwiseand_531 (
        .y(_T_816),
        .a(_T_813),
        .b(_T_815)
    );
    wire _T_817;
    BITWISEAND #(.width(1)) bitwiseand_532 (
        .y(_T_817),
        .a(_T_816),
        .b(_T_787)
    );
    wire [31:0] _GEN_32;
    MUX_UNSIGNED #(.width(32)) u_mux_533 (
        .y(_GEN_32),
        .sel(_T_817),
        .a(wdata),
        .b(_mtohost__q)
    );
    wire _T_818;
    EQ_UNSIGNED #(.width(12)) u_eq_534 (
        .y(_T_818),
        .a(csr_addr),
        .b(12'h781)
    );
    wire _T_820;
    EQ_UNSIGNED #(.width(1)) u_eq_535 (
        .y(_T_820),
        .a(_T_628),
        .b(1'h0)
    );
    wire _T_822;
    EQ_UNSIGNED #(.width(1)) u_eq_536 (
        .y(_T_822),
        .a(_T_633),
        .b(1'h0)
    );
    wire _T_823;
    BITWISEAND #(.width(1)) bitwiseand_537 (
        .y(_T_823),
        .a(_T_820),
        .b(_T_822)
    );
    wire _T_825;
    EQ_UNSIGNED #(.width(1)) u_eq_538 (
        .y(_T_825),
        .a(_T_639),
        .b(1'h0)
    );
    wire _T_826;
    BITWISEAND #(.width(1)) bitwiseand_539 (
        .y(_T_826),
        .a(_T_823),
        .b(_T_825)
    );
    wire _T_828;
    EQ_UNSIGNED #(.width(1)) u_eq_540 (
        .y(_T_828),
        .a(_T_648),
        .b(1'h0)
    );
    wire _T_829;
    BITWISEAND #(.width(1)) bitwiseand_541 (
        .y(_T_829),
        .a(_T_826),
        .b(_T_828)
    );
    wire _T_831;
    EQ_UNSIGNED #(.width(1)) u_eq_542 (
        .y(_T_831),
        .a(_T_658),
        .b(1'h0)
    );
    wire _T_832;
    BITWISEAND #(.width(1)) bitwiseand_543 (
        .y(_T_832),
        .a(_T_829),
        .b(_T_831)
    );
    wire _T_834;
    EQ_UNSIGNED #(.width(1)) u_eq_544 (
        .y(_T_834),
        .a(_T_671),
        .b(1'h0)
    );
    wire _T_835;
    BITWISEAND #(.width(1)) bitwiseand_545 (
        .y(_T_835),
        .a(_T_832),
        .b(_T_834)
    );
    wire _T_837;
    EQ_UNSIGNED #(.width(1)) u_eq_546 (
        .y(_T_837),
        .a(_T_687),
        .b(1'h0)
    );
    wire _T_838;
    BITWISEAND #(.width(1)) bitwiseand_547 (
        .y(_T_838),
        .a(_T_835),
        .b(_T_837)
    );
    wire _T_840;
    EQ_UNSIGNED #(.width(1)) u_eq_548 (
        .y(_T_840),
        .a(_T_706),
        .b(1'h0)
    );
    wire _T_841;
    BITWISEAND #(.width(1)) bitwiseand_549 (
        .y(_T_841),
        .a(_T_838),
        .b(_T_840)
    );
    wire _T_843;
    EQ_UNSIGNED #(.width(1)) u_eq_550 (
        .y(_T_843),
        .a(_T_732),
        .b(1'h0)
    );
    wire _T_844;
    BITWISEAND #(.width(1)) bitwiseand_551 (
        .y(_T_844),
        .a(_T_841),
        .b(_T_843)
    );
    wire _T_846;
    EQ_UNSIGNED #(.width(1)) u_eq_552 (
        .y(_T_846),
        .a(_T_759),
        .b(1'h0)
    );
    wire _T_847;
    BITWISEAND #(.width(1)) bitwiseand_553 (
        .y(_T_847),
        .a(_T_844),
        .b(_T_846)
    );
    wire _T_849;
    EQ_UNSIGNED #(.width(1)) u_eq_554 (
        .y(_T_849),
        .a(_T_787),
        .b(1'h0)
    );
    wire _T_850;
    BITWISEAND #(.width(1)) bitwiseand_555 (
        .y(_T_850),
        .a(_T_847),
        .b(_T_849)
    );
    wire _T_851;
    BITWISEAND #(.width(1)) bitwiseand_556 (
        .y(_T_851),
        .a(_T_850),
        .b(_T_818)
    );
    wire [31:0] _GEN_33;
    MUX_UNSIGNED #(.width(32)) u_mux_557 (
        .y(_GEN_33),
        .sel(_T_851),
        .a(wdata),
        .b(_GEN_0)
    );
    wire _T_852;
    EQ_UNSIGNED #(.width(12)) u_eq_558 (
        .y(_T_852),
        .a(csr_addr),
        .b(12'h900)
    );
    wire _T_854;
    EQ_UNSIGNED #(.width(1)) u_eq_559 (
        .y(_T_854),
        .a(_T_628),
        .b(1'h0)
    );
    wire _T_856;
    EQ_UNSIGNED #(.width(1)) u_eq_560 (
        .y(_T_856),
        .a(_T_633),
        .b(1'h0)
    );
    wire _T_857;
    BITWISEAND #(.width(1)) bitwiseand_561 (
        .y(_T_857),
        .a(_T_854),
        .b(_T_856)
    );
    wire _T_859;
    EQ_UNSIGNED #(.width(1)) u_eq_562 (
        .y(_T_859),
        .a(_T_639),
        .b(1'h0)
    );
    wire _T_860;
    BITWISEAND #(.width(1)) bitwiseand_563 (
        .y(_T_860),
        .a(_T_857),
        .b(_T_859)
    );
    wire _T_862;
    EQ_UNSIGNED #(.width(1)) u_eq_564 (
        .y(_T_862),
        .a(_T_648),
        .b(1'h0)
    );
    wire _T_863;
    BITWISEAND #(.width(1)) bitwiseand_565 (
        .y(_T_863),
        .a(_T_860),
        .b(_T_862)
    );
    wire _T_865;
    EQ_UNSIGNED #(.width(1)) u_eq_566 (
        .y(_T_865),
        .a(_T_658),
        .b(1'h0)
    );
    wire _T_866;
    BITWISEAND #(.width(1)) bitwiseand_567 (
        .y(_T_866),
        .a(_T_863),
        .b(_T_865)
    );
    wire _T_868;
    EQ_UNSIGNED #(.width(1)) u_eq_568 (
        .y(_T_868),
        .a(_T_671),
        .b(1'h0)
    );
    wire _T_869;
    BITWISEAND #(.width(1)) bitwiseand_569 (
        .y(_T_869),
        .a(_T_866),
        .b(_T_868)
    );
    wire _T_871;
    EQ_UNSIGNED #(.width(1)) u_eq_570 (
        .y(_T_871),
        .a(_T_687),
        .b(1'h0)
    );
    wire _T_872;
    BITWISEAND #(.width(1)) bitwiseand_571 (
        .y(_T_872),
        .a(_T_869),
        .b(_T_871)
    );
    wire _T_874;
    EQ_UNSIGNED #(.width(1)) u_eq_572 (
        .y(_T_874),
        .a(_T_706),
        .b(1'h0)
    );
    wire _T_875;
    BITWISEAND #(.width(1)) bitwiseand_573 (
        .y(_T_875),
        .a(_T_872),
        .b(_T_874)
    );
    wire _T_877;
    EQ_UNSIGNED #(.width(1)) u_eq_574 (
        .y(_T_877),
        .a(_T_732),
        .b(1'h0)
    );
    wire _T_878;
    BITWISEAND #(.width(1)) bitwiseand_575 (
        .y(_T_878),
        .a(_T_875),
        .b(_T_877)
    );
    wire _T_880;
    EQ_UNSIGNED #(.width(1)) u_eq_576 (
        .y(_T_880),
        .a(_T_759),
        .b(1'h0)
    );
    wire _T_881;
    BITWISEAND #(.width(1)) bitwiseand_577 (
        .y(_T_881),
        .a(_T_878),
        .b(_T_880)
    );
    wire _T_883;
    EQ_UNSIGNED #(.width(1)) u_eq_578 (
        .y(_T_883),
        .a(_T_787),
        .b(1'h0)
    );
    wire _T_884;
    BITWISEAND #(.width(1)) bitwiseand_579 (
        .y(_T_884),
        .a(_T_881),
        .b(_T_883)
    );
    wire _T_886;
    EQ_UNSIGNED #(.width(1)) u_eq_580 (
        .y(_T_886),
        .a(_T_818),
        .b(1'h0)
    );
    wire _T_887;
    BITWISEAND #(.width(1)) bitwiseand_581 (
        .y(_T_887),
        .a(_T_884),
        .b(_T_886)
    );
    wire _T_888;
    BITWISEAND #(.width(1)) bitwiseand_582 (
        .y(_T_888),
        .a(_T_887),
        .b(_T_852)
    );
    wire [31:0] _GEN_34;
    MUX_UNSIGNED #(.width(32)) u_mux_583 (
        .y(_GEN_34),
        .sel(_T_888),
        .a(wdata),
        .b(_T_572)
    );
    wire _T_889;
    EQ_UNSIGNED #(.width(12)) u_eq_584 (
        .y(_T_889),
        .a(csr_addr),
        .b(12'h901)
    );
    wire _T_891;
    EQ_UNSIGNED #(.width(1)) u_eq_585 (
        .y(_T_891),
        .a(_T_628),
        .b(1'h0)
    );
    wire _T_893;
    EQ_UNSIGNED #(.width(1)) u_eq_586 (
        .y(_T_893),
        .a(_T_633),
        .b(1'h0)
    );
    wire _T_894;
    BITWISEAND #(.width(1)) bitwiseand_587 (
        .y(_T_894),
        .a(_T_891),
        .b(_T_893)
    );
    wire _T_896;
    EQ_UNSIGNED #(.width(1)) u_eq_588 (
        .y(_T_896),
        .a(_T_639),
        .b(1'h0)
    );
    wire _T_897;
    BITWISEAND #(.width(1)) bitwiseand_589 (
        .y(_T_897),
        .a(_T_894),
        .b(_T_896)
    );
    wire _T_899;
    EQ_UNSIGNED #(.width(1)) u_eq_590 (
        .y(_T_899),
        .a(_T_648),
        .b(1'h0)
    );
    wire _T_900;
    BITWISEAND #(.width(1)) bitwiseand_591 (
        .y(_T_900),
        .a(_T_897),
        .b(_T_899)
    );
    wire _T_902;
    EQ_UNSIGNED #(.width(1)) u_eq_592 (
        .y(_T_902),
        .a(_T_658),
        .b(1'h0)
    );
    wire _T_903;
    BITWISEAND #(.width(1)) bitwiseand_593 (
        .y(_T_903),
        .a(_T_900),
        .b(_T_902)
    );
    wire _T_905;
    EQ_UNSIGNED #(.width(1)) u_eq_594 (
        .y(_T_905),
        .a(_T_671),
        .b(1'h0)
    );
    wire _T_906;
    BITWISEAND #(.width(1)) bitwiseand_595 (
        .y(_T_906),
        .a(_T_903),
        .b(_T_905)
    );
    wire _T_908;
    EQ_UNSIGNED #(.width(1)) u_eq_596 (
        .y(_T_908),
        .a(_T_687),
        .b(1'h0)
    );
    wire _T_909;
    BITWISEAND #(.width(1)) bitwiseand_597 (
        .y(_T_909),
        .a(_T_906),
        .b(_T_908)
    );
    wire _T_911;
    EQ_UNSIGNED #(.width(1)) u_eq_598 (
        .y(_T_911),
        .a(_T_706),
        .b(1'h0)
    );
    wire _T_912;
    BITWISEAND #(.width(1)) bitwiseand_599 (
        .y(_T_912),
        .a(_T_909),
        .b(_T_911)
    );
    wire _T_914;
    EQ_UNSIGNED #(.width(1)) u_eq_600 (
        .y(_T_914),
        .a(_T_732),
        .b(1'h0)
    );
    wire _T_915;
    BITWISEAND #(.width(1)) bitwiseand_601 (
        .y(_T_915),
        .a(_T_912),
        .b(_T_914)
    );
    wire _T_917;
    EQ_UNSIGNED #(.width(1)) u_eq_602 (
        .y(_T_917),
        .a(_T_759),
        .b(1'h0)
    );
    wire _T_918;
    BITWISEAND #(.width(1)) bitwiseand_603 (
        .y(_T_918),
        .a(_T_915),
        .b(_T_917)
    );
    wire _T_920;
    EQ_UNSIGNED #(.width(1)) u_eq_604 (
        .y(_T_920),
        .a(_T_787),
        .b(1'h0)
    );
    wire _T_921;
    BITWISEAND #(.width(1)) bitwiseand_605 (
        .y(_T_921),
        .a(_T_918),
        .b(_T_920)
    );
    wire _T_923;
    EQ_UNSIGNED #(.width(1)) u_eq_606 (
        .y(_T_923),
        .a(_T_818),
        .b(1'h0)
    );
    wire _T_924;
    BITWISEAND #(.width(1)) bitwiseand_607 (
        .y(_T_924),
        .a(_T_921),
        .b(_T_923)
    );
    wire _T_926;
    EQ_UNSIGNED #(.width(1)) u_eq_608 (
        .y(_T_926),
        .a(_T_852),
        .b(1'h0)
    );
    wire _T_927;
    BITWISEAND #(.width(1)) bitwiseand_609 (
        .y(_T_927),
        .a(_T_924),
        .b(_T_926)
    );
    wire _T_928;
    BITWISEAND #(.width(1)) bitwiseand_610 (
        .y(_T_928),
        .a(_T_927),
        .b(_T_889)
    );
    wire [31:0] _GEN_35;
    MUX_UNSIGNED #(.width(32)) u_mux_611 (
        .y(_GEN_35),
        .sel(_T_928),
        .a(wdata),
        .b(_GEN_25)
    );
    wire _T_929;
    EQ_UNSIGNED #(.width(12)) u_eq_612 (
        .y(_T_929),
        .a(csr_addr),
        .b(12'h902)
    );
    wire _T_931;
    EQ_UNSIGNED #(.width(1)) u_eq_613 (
        .y(_T_931),
        .a(_T_628),
        .b(1'h0)
    );
    wire _T_933;
    EQ_UNSIGNED #(.width(1)) u_eq_614 (
        .y(_T_933),
        .a(_T_633),
        .b(1'h0)
    );
    wire _T_934;
    BITWISEAND #(.width(1)) bitwiseand_615 (
        .y(_T_934),
        .a(_T_931),
        .b(_T_933)
    );
    wire _T_936;
    EQ_UNSIGNED #(.width(1)) u_eq_616 (
        .y(_T_936),
        .a(_T_639),
        .b(1'h0)
    );
    wire _T_937;
    BITWISEAND #(.width(1)) bitwiseand_617 (
        .y(_T_937),
        .a(_T_934),
        .b(_T_936)
    );
    wire _T_939;
    EQ_UNSIGNED #(.width(1)) u_eq_618 (
        .y(_T_939),
        .a(_T_648),
        .b(1'h0)
    );
    wire _T_940;
    BITWISEAND #(.width(1)) bitwiseand_619 (
        .y(_T_940),
        .a(_T_937),
        .b(_T_939)
    );
    wire _T_942;
    EQ_UNSIGNED #(.width(1)) u_eq_620 (
        .y(_T_942),
        .a(_T_658),
        .b(1'h0)
    );
    wire _T_943;
    BITWISEAND #(.width(1)) bitwiseand_621 (
        .y(_T_943),
        .a(_T_940),
        .b(_T_942)
    );
    wire _T_945;
    EQ_UNSIGNED #(.width(1)) u_eq_622 (
        .y(_T_945),
        .a(_T_671),
        .b(1'h0)
    );
    wire _T_946;
    BITWISEAND #(.width(1)) bitwiseand_623 (
        .y(_T_946),
        .a(_T_943),
        .b(_T_945)
    );
    wire _T_948;
    EQ_UNSIGNED #(.width(1)) u_eq_624 (
        .y(_T_948),
        .a(_T_687),
        .b(1'h0)
    );
    wire _T_949;
    BITWISEAND #(.width(1)) bitwiseand_625 (
        .y(_T_949),
        .a(_T_946),
        .b(_T_948)
    );
    wire _T_951;
    EQ_UNSIGNED #(.width(1)) u_eq_626 (
        .y(_T_951),
        .a(_T_706),
        .b(1'h0)
    );
    wire _T_952;
    BITWISEAND #(.width(1)) bitwiseand_627 (
        .y(_T_952),
        .a(_T_949),
        .b(_T_951)
    );
    wire _T_954;
    EQ_UNSIGNED #(.width(1)) u_eq_628 (
        .y(_T_954),
        .a(_T_732),
        .b(1'h0)
    );
    wire _T_955;
    BITWISEAND #(.width(1)) bitwiseand_629 (
        .y(_T_955),
        .a(_T_952),
        .b(_T_954)
    );
    wire _T_957;
    EQ_UNSIGNED #(.width(1)) u_eq_630 (
        .y(_T_957),
        .a(_T_759),
        .b(1'h0)
    );
    wire _T_958;
    BITWISEAND #(.width(1)) bitwiseand_631 (
        .y(_T_958),
        .a(_T_955),
        .b(_T_957)
    );
    wire _T_960;
    EQ_UNSIGNED #(.width(1)) u_eq_632 (
        .y(_T_960),
        .a(_T_787),
        .b(1'h0)
    );
    wire _T_961;
    BITWISEAND #(.width(1)) bitwiseand_633 (
        .y(_T_961),
        .a(_T_958),
        .b(_T_960)
    );
    wire _T_963;
    EQ_UNSIGNED #(.width(1)) u_eq_634 (
        .y(_T_963),
        .a(_T_818),
        .b(1'h0)
    );
    wire _T_964;
    BITWISEAND #(.width(1)) bitwiseand_635 (
        .y(_T_964),
        .a(_T_961),
        .b(_T_963)
    );
    wire _T_966;
    EQ_UNSIGNED #(.width(1)) u_eq_636 (
        .y(_T_966),
        .a(_T_852),
        .b(1'h0)
    );
    wire _T_967;
    BITWISEAND #(.width(1)) bitwiseand_637 (
        .y(_T_967),
        .a(_T_964),
        .b(_T_966)
    );
    wire _T_969;
    EQ_UNSIGNED #(.width(1)) u_eq_638 (
        .y(_T_969),
        .a(_T_889),
        .b(1'h0)
    );
    wire _T_970;
    BITWISEAND #(.width(1)) bitwiseand_639 (
        .y(_T_970),
        .a(_T_967),
        .b(_T_969)
    );
    wire _T_971;
    BITWISEAND #(.width(1)) bitwiseand_640 (
        .y(_T_971),
        .a(_T_970),
        .b(_T_929)
    );
    wire [31:0] _GEN_36;
    MUX_UNSIGNED #(.width(32)) u_mux_641 (
        .y(_GEN_36),
        .sel(_T_971),
        .a(wdata),
        .b(_GEN_3)
    );
    wire _T_972;
    EQ_UNSIGNED #(.width(12)) u_eq_642 (
        .y(_T_972),
        .a(csr_addr),
        .b(12'h980)
    );
    wire _T_974;
    EQ_UNSIGNED #(.width(1)) u_eq_643 (
        .y(_T_974),
        .a(_T_628),
        .b(1'h0)
    );
    wire _T_976;
    EQ_UNSIGNED #(.width(1)) u_eq_644 (
        .y(_T_976),
        .a(_T_633),
        .b(1'h0)
    );
    wire _T_977;
    BITWISEAND #(.width(1)) bitwiseand_645 (
        .y(_T_977),
        .a(_T_974),
        .b(_T_976)
    );
    wire _T_979;
    EQ_UNSIGNED #(.width(1)) u_eq_646 (
        .y(_T_979),
        .a(_T_639),
        .b(1'h0)
    );
    wire _T_980;
    BITWISEAND #(.width(1)) bitwiseand_647 (
        .y(_T_980),
        .a(_T_977),
        .b(_T_979)
    );
    wire _T_982;
    EQ_UNSIGNED #(.width(1)) u_eq_648 (
        .y(_T_982),
        .a(_T_648),
        .b(1'h0)
    );
    wire _T_983;
    BITWISEAND #(.width(1)) bitwiseand_649 (
        .y(_T_983),
        .a(_T_980),
        .b(_T_982)
    );
    wire _T_985;
    EQ_UNSIGNED #(.width(1)) u_eq_650 (
        .y(_T_985),
        .a(_T_658),
        .b(1'h0)
    );
    wire _T_986;
    BITWISEAND #(.width(1)) bitwiseand_651 (
        .y(_T_986),
        .a(_T_983),
        .b(_T_985)
    );
    wire _T_988;
    EQ_UNSIGNED #(.width(1)) u_eq_652 (
        .y(_T_988),
        .a(_T_671),
        .b(1'h0)
    );
    wire _T_989;
    BITWISEAND #(.width(1)) bitwiseand_653 (
        .y(_T_989),
        .a(_T_986),
        .b(_T_988)
    );
    wire _T_991;
    EQ_UNSIGNED #(.width(1)) u_eq_654 (
        .y(_T_991),
        .a(_T_687),
        .b(1'h0)
    );
    wire _T_992;
    BITWISEAND #(.width(1)) bitwiseand_655 (
        .y(_T_992),
        .a(_T_989),
        .b(_T_991)
    );
    wire _T_994;
    EQ_UNSIGNED #(.width(1)) u_eq_656 (
        .y(_T_994),
        .a(_T_706),
        .b(1'h0)
    );
    wire _T_995;
    BITWISEAND #(.width(1)) bitwiseand_657 (
        .y(_T_995),
        .a(_T_992),
        .b(_T_994)
    );
    wire _T_997;
    EQ_UNSIGNED #(.width(1)) u_eq_658 (
        .y(_T_997),
        .a(_T_732),
        .b(1'h0)
    );
    wire _T_998;
    BITWISEAND #(.width(1)) bitwiseand_659 (
        .y(_T_998),
        .a(_T_995),
        .b(_T_997)
    );
    wire _T_1000;
    EQ_UNSIGNED #(.width(1)) u_eq_660 (
        .y(_T_1000),
        .a(_T_759),
        .b(1'h0)
    );
    wire _T_1001;
    BITWISEAND #(.width(1)) bitwiseand_661 (
        .y(_T_1001),
        .a(_T_998),
        .b(_T_1000)
    );
    wire _T_1003;
    EQ_UNSIGNED #(.width(1)) u_eq_662 (
        .y(_T_1003),
        .a(_T_787),
        .b(1'h0)
    );
    wire _T_1004;
    BITWISEAND #(.width(1)) bitwiseand_663 (
        .y(_T_1004),
        .a(_T_1001),
        .b(_T_1003)
    );
    wire _T_1006;
    EQ_UNSIGNED #(.width(1)) u_eq_664 (
        .y(_T_1006),
        .a(_T_818),
        .b(1'h0)
    );
    wire _T_1007;
    BITWISEAND #(.width(1)) bitwiseand_665 (
        .y(_T_1007),
        .a(_T_1004),
        .b(_T_1006)
    );
    wire _T_1009;
    EQ_UNSIGNED #(.width(1)) u_eq_666 (
        .y(_T_1009),
        .a(_T_852),
        .b(1'h0)
    );
    wire _T_1010;
    BITWISEAND #(.width(1)) bitwiseand_667 (
        .y(_T_1010),
        .a(_T_1007),
        .b(_T_1009)
    );
    wire _T_1012;
    EQ_UNSIGNED #(.width(1)) u_eq_668 (
        .y(_T_1012),
        .a(_T_889),
        .b(1'h0)
    );
    wire _T_1013;
    BITWISEAND #(.width(1)) bitwiseand_669 (
        .y(_T_1013),
        .a(_T_1010),
        .b(_T_1012)
    );
    wire _T_1015;
    EQ_UNSIGNED #(.width(1)) u_eq_670 (
        .y(_T_1015),
        .a(_T_929),
        .b(1'h0)
    );
    wire _T_1016;
    BITWISEAND #(.width(1)) bitwiseand_671 (
        .y(_T_1016),
        .a(_T_1013),
        .b(_T_1015)
    );
    wire _T_1017;
    BITWISEAND #(.width(1)) bitwiseand_672 (
        .y(_T_1017),
        .a(_T_1016),
        .b(_T_972)
    );
    wire [31:0] _GEN_37;
    MUX_UNSIGNED #(.width(32)) u_mux_673 (
        .y(_GEN_37),
        .sel(_T_1017),
        .a(wdata),
        .b(_GEN_2)
    );
    wire _T_1018;
    EQ_UNSIGNED #(.width(12)) u_eq_674 (
        .y(_T_1018),
        .a(csr_addr),
        .b(12'h981)
    );
    wire _T_1020;
    EQ_UNSIGNED #(.width(1)) u_eq_675 (
        .y(_T_1020),
        .a(_T_628),
        .b(1'h0)
    );
    wire _T_1022;
    EQ_UNSIGNED #(.width(1)) u_eq_676 (
        .y(_T_1022),
        .a(_T_633),
        .b(1'h0)
    );
    wire _T_1023;
    BITWISEAND #(.width(1)) bitwiseand_677 (
        .y(_T_1023),
        .a(_T_1020),
        .b(_T_1022)
    );
    wire _T_1025;
    EQ_UNSIGNED #(.width(1)) u_eq_678 (
        .y(_T_1025),
        .a(_T_639),
        .b(1'h0)
    );
    wire _T_1026;
    BITWISEAND #(.width(1)) bitwiseand_679 (
        .y(_T_1026),
        .a(_T_1023),
        .b(_T_1025)
    );
    wire _T_1028;
    EQ_UNSIGNED #(.width(1)) u_eq_680 (
        .y(_T_1028),
        .a(_T_648),
        .b(1'h0)
    );
    wire _T_1029;
    BITWISEAND #(.width(1)) bitwiseand_681 (
        .y(_T_1029),
        .a(_T_1026),
        .b(_T_1028)
    );
    wire _T_1031;
    EQ_UNSIGNED #(.width(1)) u_eq_682 (
        .y(_T_1031),
        .a(_T_658),
        .b(1'h0)
    );
    wire _T_1032;
    BITWISEAND #(.width(1)) bitwiseand_683 (
        .y(_T_1032),
        .a(_T_1029),
        .b(_T_1031)
    );
    wire _T_1034;
    EQ_UNSIGNED #(.width(1)) u_eq_684 (
        .y(_T_1034),
        .a(_T_671),
        .b(1'h0)
    );
    wire _T_1035;
    BITWISEAND #(.width(1)) bitwiseand_685 (
        .y(_T_1035),
        .a(_T_1032),
        .b(_T_1034)
    );
    wire _T_1037;
    EQ_UNSIGNED #(.width(1)) u_eq_686 (
        .y(_T_1037),
        .a(_T_687),
        .b(1'h0)
    );
    wire _T_1038;
    BITWISEAND #(.width(1)) bitwiseand_687 (
        .y(_T_1038),
        .a(_T_1035),
        .b(_T_1037)
    );
    wire _T_1040;
    EQ_UNSIGNED #(.width(1)) u_eq_688 (
        .y(_T_1040),
        .a(_T_706),
        .b(1'h0)
    );
    wire _T_1041;
    BITWISEAND #(.width(1)) bitwiseand_689 (
        .y(_T_1041),
        .a(_T_1038),
        .b(_T_1040)
    );
    wire _T_1043;
    EQ_UNSIGNED #(.width(1)) u_eq_690 (
        .y(_T_1043),
        .a(_T_732),
        .b(1'h0)
    );
    wire _T_1044;
    BITWISEAND #(.width(1)) bitwiseand_691 (
        .y(_T_1044),
        .a(_T_1041),
        .b(_T_1043)
    );
    wire _T_1046;
    EQ_UNSIGNED #(.width(1)) u_eq_692 (
        .y(_T_1046),
        .a(_T_759),
        .b(1'h0)
    );
    wire _T_1047;
    BITWISEAND #(.width(1)) bitwiseand_693 (
        .y(_T_1047),
        .a(_T_1044),
        .b(_T_1046)
    );
    wire _T_1049;
    EQ_UNSIGNED #(.width(1)) u_eq_694 (
        .y(_T_1049),
        .a(_T_787),
        .b(1'h0)
    );
    wire _T_1050;
    BITWISEAND #(.width(1)) bitwiseand_695 (
        .y(_T_1050),
        .a(_T_1047),
        .b(_T_1049)
    );
    wire _T_1052;
    EQ_UNSIGNED #(.width(1)) u_eq_696 (
        .y(_T_1052),
        .a(_T_818),
        .b(1'h0)
    );
    wire _T_1053;
    BITWISEAND #(.width(1)) bitwiseand_697 (
        .y(_T_1053),
        .a(_T_1050),
        .b(_T_1052)
    );
    wire _T_1055;
    EQ_UNSIGNED #(.width(1)) u_eq_698 (
        .y(_T_1055),
        .a(_T_852),
        .b(1'h0)
    );
    wire _T_1056;
    BITWISEAND #(.width(1)) bitwiseand_699 (
        .y(_T_1056),
        .a(_T_1053),
        .b(_T_1055)
    );
    wire _T_1058;
    EQ_UNSIGNED #(.width(1)) u_eq_700 (
        .y(_T_1058),
        .a(_T_889),
        .b(1'h0)
    );
    wire _T_1059;
    BITWISEAND #(.width(1)) bitwiseand_701 (
        .y(_T_1059),
        .a(_T_1056),
        .b(_T_1058)
    );
    wire _T_1061;
    EQ_UNSIGNED #(.width(1)) u_eq_702 (
        .y(_T_1061),
        .a(_T_929),
        .b(1'h0)
    );
    wire _T_1062;
    BITWISEAND #(.width(1)) bitwiseand_703 (
        .y(_T_1062),
        .a(_T_1059),
        .b(_T_1061)
    );
    wire _T_1064;
    EQ_UNSIGNED #(.width(1)) u_eq_704 (
        .y(_T_1064),
        .a(_T_972),
        .b(1'h0)
    );
    wire _T_1065;
    BITWISEAND #(.width(1)) bitwiseand_705 (
        .y(_T_1065),
        .a(_T_1062),
        .b(_T_1064)
    );
    wire _T_1066;
    BITWISEAND #(.width(1)) bitwiseand_706 (
        .y(_T_1066),
        .a(_T_1065),
        .b(_T_1018)
    );
    wire [31:0] _GEN_38;
    MUX_UNSIGNED #(.width(32)) u_mux_707 (
        .y(_GEN_38),
        .sel(_T_1066),
        .a(wdata),
        .b(_GEN_26)
    );
    wire _T_1067;
    EQ_UNSIGNED #(.width(12)) u_eq_708 (
        .y(_T_1067),
        .a(csr_addr),
        .b(12'h982)
    );
    wire _T_1069;
    EQ_UNSIGNED #(.width(1)) u_eq_709 (
        .y(_T_1069),
        .a(_T_628),
        .b(1'h0)
    );
    wire _T_1071;
    EQ_UNSIGNED #(.width(1)) u_eq_710 (
        .y(_T_1071),
        .a(_T_633),
        .b(1'h0)
    );
    wire _T_1072;
    BITWISEAND #(.width(1)) bitwiseand_711 (
        .y(_T_1072),
        .a(_T_1069),
        .b(_T_1071)
    );
    wire _T_1074;
    EQ_UNSIGNED #(.width(1)) u_eq_712 (
        .y(_T_1074),
        .a(_T_639),
        .b(1'h0)
    );
    wire _T_1075;
    BITWISEAND #(.width(1)) bitwiseand_713 (
        .y(_T_1075),
        .a(_T_1072),
        .b(_T_1074)
    );
    wire _T_1077;
    EQ_UNSIGNED #(.width(1)) u_eq_714 (
        .y(_T_1077),
        .a(_T_648),
        .b(1'h0)
    );
    wire _T_1078;
    BITWISEAND #(.width(1)) bitwiseand_715 (
        .y(_T_1078),
        .a(_T_1075),
        .b(_T_1077)
    );
    wire _T_1080;
    EQ_UNSIGNED #(.width(1)) u_eq_716 (
        .y(_T_1080),
        .a(_T_658),
        .b(1'h0)
    );
    wire _T_1081;
    BITWISEAND #(.width(1)) bitwiseand_717 (
        .y(_T_1081),
        .a(_T_1078),
        .b(_T_1080)
    );
    wire _T_1083;
    EQ_UNSIGNED #(.width(1)) u_eq_718 (
        .y(_T_1083),
        .a(_T_671),
        .b(1'h0)
    );
    wire _T_1084;
    BITWISEAND #(.width(1)) bitwiseand_719 (
        .y(_T_1084),
        .a(_T_1081),
        .b(_T_1083)
    );
    wire _T_1086;
    EQ_UNSIGNED #(.width(1)) u_eq_720 (
        .y(_T_1086),
        .a(_T_687),
        .b(1'h0)
    );
    wire _T_1087;
    BITWISEAND #(.width(1)) bitwiseand_721 (
        .y(_T_1087),
        .a(_T_1084),
        .b(_T_1086)
    );
    wire _T_1089;
    EQ_UNSIGNED #(.width(1)) u_eq_722 (
        .y(_T_1089),
        .a(_T_706),
        .b(1'h0)
    );
    wire _T_1090;
    BITWISEAND #(.width(1)) bitwiseand_723 (
        .y(_T_1090),
        .a(_T_1087),
        .b(_T_1089)
    );
    wire _T_1092;
    EQ_UNSIGNED #(.width(1)) u_eq_724 (
        .y(_T_1092),
        .a(_T_732),
        .b(1'h0)
    );
    wire _T_1093;
    BITWISEAND #(.width(1)) bitwiseand_725 (
        .y(_T_1093),
        .a(_T_1090),
        .b(_T_1092)
    );
    wire _T_1095;
    EQ_UNSIGNED #(.width(1)) u_eq_726 (
        .y(_T_1095),
        .a(_T_759),
        .b(1'h0)
    );
    wire _T_1096;
    BITWISEAND #(.width(1)) bitwiseand_727 (
        .y(_T_1096),
        .a(_T_1093),
        .b(_T_1095)
    );
    wire _T_1098;
    EQ_UNSIGNED #(.width(1)) u_eq_728 (
        .y(_T_1098),
        .a(_T_787),
        .b(1'h0)
    );
    wire _T_1099;
    BITWISEAND #(.width(1)) bitwiseand_729 (
        .y(_T_1099),
        .a(_T_1096),
        .b(_T_1098)
    );
    wire _T_1101;
    EQ_UNSIGNED #(.width(1)) u_eq_730 (
        .y(_T_1101),
        .a(_T_818),
        .b(1'h0)
    );
    wire _T_1102;
    BITWISEAND #(.width(1)) bitwiseand_731 (
        .y(_T_1102),
        .a(_T_1099),
        .b(_T_1101)
    );
    wire _T_1104;
    EQ_UNSIGNED #(.width(1)) u_eq_732 (
        .y(_T_1104),
        .a(_T_852),
        .b(1'h0)
    );
    wire _T_1105;
    BITWISEAND #(.width(1)) bitwiseand_733 (
        .y(_T_1105),
        .a(_T_1102),
        .b(_T_1104)
    );
    wire _T_1107;
    EQ_UNSIGNED #(.width(1)) u_eq_734 (
        .y(_T_1107),
        .a(_T_889),
        .b(1'h0)
    );
    wire _T_1108;
    BITWISEAND #(.width(1)) bitwiseand_735 (
        .y(_T_1108),
        .a(_T_1105),
        .b(_T_1107)
    );
    wire _T_1110;
    EQ_UNSIGNED #(.width(1)) u_eq_736 (
        .y(_T_1110),
        .a(_T_929),
        .b(1'h0)
    );
    wire _T_1111;
    BITWISEAND #(.width(1)) bitwiseand_737 (
        .y(_T_1111),
        .a(_T_1108),
        .b(_T_1110)
    );
    wire _T_1113;
    EQ_UNSIGNED #(.width(1)) u_eq_738 (
        .y(_T_1113),
        .a(_T_972),
        .b(1'h0)
    );
    wire _T_1114;
    BITWISEAND #(.width(1)) bitwiseand_739 (
        .y(_T_1114),
        .a(_T_1111),
        .b(_T_1113)
    );
    wire _T_1116;
    EQ_UNSIGNED #(.width(1)) u_eq_740 (
        .y(_T_1116),
        .a(_T_1018),
        .b(1'h0)
    );
    wire _T_1117;
    BITWISEAND #(.width(1)) bitwiseand_741 (
        .y(_T_1117),
        .a(_T_1114),
        .b(_T_1116)
    );
    wire _T_1118;
    BITWISEAND #(.width(1)) bitwiseand_742 (
        .y(_T_1118),
        .a(_T_1117),
        .b(_T_1067)
    );
    wire [31:0] _GEN_39;
    MUX_UNSIGNED #(.width(32)) u_mux_743 (
        .y(_GEN_39),
        .sel(_T_1118),
        .a(wdata),
        .b(_GEN_4)
    );
    wire [1:0] _GEN_40;
    MUX_UNSIGNED #(.width(2)) u_mux_744 (
        .y(_GEN_40),
        .sel(_T_627),
        .a(_GEN_17),
        .b(_GEN_15)
    );
    wire _GEN_41;
    MUX_UNSIGNED #(.width(1)) u_mux_745 (
        .y(_GEN_41),
        .sel(_T_627),
        .a(_GEN_18),
        .b(_GEN_16)
    );
    wire [1:0] _GEN_42;
    MUX_UNSIGNED #(.width(2)) u_mux_746 (
        .y(_GEN_42),
        .sel(_T_627),
        .a(_GEN_19),
        .b(_GEN_13)
    );
    wire _GEN_43;
    MUX_UNSIGNED #(.width(1)) u_mux_747 (
        .y(_GEN_43),
        .sel(_T_627),
        .a(_GEN_20),
        .b(_GEN_14)
    );
    wire _GEN_44;
    MUX_UNSIGNED #(.width(1)) u_mux_748 (
        .y(_GEN_44),
        .sel(_T_627),
        .a(_GEN_21),
        .b(_MTIP__q)
    );
    wire _GEN_45;
    MUX_UNSIGNED #(.width(1)) u_mux_749 (
        .y(_GEN_45),
        .sel(_T_627),
        .a(_GEN_22),
        .b(_MSIP__q)
    );
    wire _GEN_46;
    MUX_UNSIGNED #(.width(1)) u_mux_750 (
        .y(_GEN_46),
        .sel(_T_627),
        .a(_GEN_23),
        .b(_MTIE__q)
    );
    wire _GEN_47;
    MUX_UNSIGNED #(.width(1)) u_mux_751 (
        .y(_GEN_47),
        .sel(_T_627),
        .a(_GEN_24),
        .b(_MSIE__q)
    );
    wire [31:0] _GEN_48;
    MUX_UNSIGNED #(.width(32)) u_mux_752 (
        .y(_GEN_48),
        .sel(_T_627),
        .a(_GEN_35),
        .b(_T_563)
    );
    wire [31:0] _GEN_49;
    MUX_UNSIGNED #(.width(32)) u_mux_753 (
        .y(_GEN_49),
        .sel(_T_627),
        .a(_GEN_38),
        .b(_GEN_1)
    );
    wire [31:0] _GEN_50;
    MUX_UNSIGNED #(.width(32)) u_mux_754 (
        .y(_GEN_50),
        .sel(_T_627),
        .a(_GEN_27),
        .b(_mtimecmp__q)
    );
    wire [31:0] _GEN_51;
    MUX_UNSIGNED #(.width(32)) u_mux_755 (
        .y(_GEN_51),
        .sel(_T_627),
        .a(_GEN_28),
        .b(_mscratch__q)
    );
    wire [34:0] _GEN_52;
    wire [34:0] _WTEMP_52;
    PAD_UNSIGNED #(.width(32), .n(35)) u_pad_756 (
        .y(_WTEMP_52),
        .in(_GEN_6)
    );
    MUX_UNSIGNED #(.width(35)) u_mux_757 (
        .y(_GEN_52),
        .sel(_T_627),
        .a(_GEN_29),
        .b(_WTEMP_52)
    );
    wire [31:0] _GEN_53;
    MUX_UNSIGNED #(.width(32)) u_mux_758 (
        .y(_GEN_53),
        .sel(_T_627),
        .a(_GEN_30),
        .b(_GEN_7)
    );
    wire [31:0] _GEN_54;
    MUX_UNSIGNED #(.width(32)) u_mux_759 (
        .y(_GEN_54),
        .sel(_T_627),
        .a(_GEN_31),
        .b(_GEN_12)
    );
    wire [31:0] _GEN_55;
    MUX_UNSIGNED #(.width(32)) u_mux_760 (
        .y(_GEN_55),
        .sel(_T_627),
        .a(_GEN_32),
        .b(_mtohost__q)
    );
    wire [31:0] _GEN_56;
    MUX_UNSIGNED #(.width(32)) u_mux_761 (
        .y(_GEN_56),
        .sel(_T_627),
        .a(_GEN_33),
        .b(_GEN_0)
    );
    wire [31:0] _GEN_57;
    MUX_UNSIGNED #(.width(32)) u_mux_762 (
        .y(_GEN_57),
        .sel(_T_627),
        .a(_GEN_34),
        .b(_T_572)
    );
    wire [31:0] _GEN_58;
    MUX_UNSIGNED #(.width(32)) u_mux_763 (
        .y(_GEN_58),
        .sel(_T_627),
        .a(_GEN_36),
        .b(_GEN_3)
    );
    wire [31:0] _GEN_59;
    MUX_UNSIGNED #(.width(32)) u_mux_764 (
        .y(_GEN_59),
        .sel(_T_627),
        .a(_GEN_37),
        .b(_GEN_2)
    );
    wire [31:0] _GEN_60;
    MUX_UNSIGNED #(.width(32)) u_mux_765 (
        .y(_GEN_60),
        .sel(_T_627),
        .a(_GEN_39),
        .b(_GEN_4)
    );
    wire [34:0] _GEN_61;
    wire [34:0] _WTEMP_53;
    PAD_UNSIGNED #(.width(32), .n(35)) u_pad_766 (
        .y(_WTEMP_53),
        .in(_mepc__q)
    );
    MUX_UNSIGNED #(.width(35)) u_mux_767 (
        .y(_GEN_61),
        .sel(_T_599),
        .a(_GEN_52),
        .b(_WTEMP_53)
    );
    wire [31:0] _GEN_62;
    MUX_UNSIGNED #(.width(32)) u_mux_768 (
        .y(_GEN_62),
        .sel(_T_599),
        .a(_GEN_53),
        .b(_mcause__q)
    );
    wire [1:0] _GEN_63;
    MUX_UNSIGNED #(.width(2)) u_mux_769 (
        .y(_GEN_63),
        .sel(_T_599),
        .a(_GEN_42),
        .b(_PRV__q)
    );
    wire _GEN_64;
    MUX_UNSIGNED #(.width(1)) u_mux_770 (
        .y(_GEN_64),
        .sel(_T_599),
        .a(_GEN_43),
        .b(_IE__q)
    );
    wire [1:0] _GEN_65;
    MUX_UNSIGNED #(.width(2)) u_mux_771 (
        .y(_GEN_65),
        .sel(_T_599),
        .a(_GEN_40),
        .b(_PRV1__q)
    );
    wire _GEN_66;
    MUX_UNSIGNED #(.width(1)) u_mux_772 (
        .y(_GEN_66),
        .sel(_T_599),
        .a(_GEN_41),
        .b(_IE1__q)
    );
    wire [31:0] _GEN_67;
    MUX_UNSIGNED #(.width(32)) u_mux_773 (
        .y(_GEN_67),
        .sel(_T_599),
        .a(_GEN_54),
        .b(_mbadaddr__q)
    );
    wire _GEN_68;
    MUX_UNSIGNED #(.width(1)) u_mux_774 (
        .y(_GEN_68),
        .sel(_T_599),
        .a(_GEN_44),
        .b(_MTIP__q)
    );
    wire _GEN_69;
    MUX_UNSIGNED #(.width(1)) u_mux_775 (
        .y(_GEN_69),
        .sel(_T_599),
        .a(_GEN_45),
        .b(_MSIP__q)
    );
    wire _GEN_70;
    MUX_UNSIGNED #(.width(1)) u_mux_776 (
        .y(_GEN_70),
        .sel(_T_599),
        .a(_GEN_46),
        .b(_MTIE__q)
    );
    wire _GEN_71;
    MUX_UNSIGNED #(.width(1)) u_mux_777 (
        .y(_GEN_71),
        .sel(_T_599),
        .a(_GEN_47),
        .b(_MSIE__q)
    );
    wire [31:0] _GEN_72;
    MUX_UNSIGNED #(.width(32)) u_mux_778 (
        .y(_GEN_72),
        .sel(_T_599),
        .a(_GEN_48),
        .b(_T_563)
    );
    wire [31:0] _GEN_73;
    MUX_UNSIGNED #(.width(32)) u_mux_779 (
        .y(_GEN_73),
        .sel(_T_599),
        .a(_GEN_49),
        .b(_GEN_1)
    );
    wire [31:0] _GEN_74;
    MUX_UNSIGNED #(.width(32)) u_mux_780 (
        .y(_GEN_74),
        .sel(_T_599),
        .a(_GEN_50),
        .b(_mtimecmp__q)
    );
    wire [31:0] _GEN_75;
    MUX_UNSIGNED #(.width(32)) u_mux_781 (
        .y(_GEN_75),
        .sel(_T_599),
        .a(_GEN_51),
        .b(_mscratch__q)
    );
    wire [31:0] _GEN_76;
    MUX_UNSIGNED #(.width(32)) u_mux_782 (
        .y(_GEN_76),
        .sel(_T_599),
        .a(_GEN_55),
        .b(_mtohost__q)
    );
    wire [31:0] _GEN_77;
    MUX_UNSIGNED #(.width(32)) u_mux_783 (
        .y(_GEN_77),
        .sel(_T_599),
        .a(_GEN_56),
        .b(_GEN_0)
    );
    wire [31:0] _GEN_78;
    MUX_UNSIGNED #(.width(32)) u_mux_784 (
        .y(_GEN_78),
        .sel(_T_599),
        .a(_GEN_57),
        .b(_T_572)
    );
    wire [31:0] _GEN_79;
    MUX_UNSIGNED #(.width(32)) u_mux_785 (
        .y(_GEN_79),
        .sel(_T_599),
        .a(_GEN_58),
        .b(_GEN_3)
    );
    wire [31:0] _GEN_80;
    MUX_UNSIGNED #(.width(32)) u_mux_786 (
        .y(_GEN_80),
        .sel(_T_599),
        .a(_GEN_59),
        .b(_GEN_2)
    );
    wire [31:0] _GEN_81;
    MUX_UNSIGNED #(.width(32)) u_mux_787 (
        .y(_GEN_81),
        .sel(_T_599),
        .a(_GEN_60),
        .b(_GEN_4)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_788 (
        .y(_IE__d),
        .sel(reset),
        .a(1'h0),
        .b(_GEN_64)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_789 (
        .y(_IE1__d),
        .sel(reset),
        .a(1'h0),
        .b(_GEN_66)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_790 (
        .y(_MSIE__d),
        .sel(reset),
        .a(1'h0),
        .b(_GEN_71)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_791 (
        .y(_MSIP__d),
        .sel(reset),
        .a(1'h0),
        .b(_GEN_69)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_792 (
        .y(_MTIE__d),
        .sel(reset),
        .a(1'h0),
        .b(_GEN_70)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_793 (
        .y(_MTIP__d),
        .sel(reset),
        .a(1'h0),
        .b(_GEN_68)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_794 (
        .y(_PRV__d),
        .sel(reset),
        .a(2'h3),
        .b(_GEN_63)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_795 (
        .y(_PRV1__d),
        .sel(reset),
        .a(2'h3),
        .b(_GEN_65)
    );
    MUX_UNSIGNED #(.width(32)) u_mux_796 (
        .y(_cycle__d),
        .sel(reset),
        .a(32'h0),
        .b(_GEN_78)
    );
    MUX_UNSIGNED #(.width(32)) u_mux_797 (
        .y(_cycleh__d),
        .sel(reset),
        .a(32'h0),
        .b(_GEN_80)
    );
    MUX_UNSIGNED #(.width(32)) u_mux_798 (
        .y(_instret__d),
        .sel(reset),
        .a(32'h0),
        .b(_GEN_79)
    );
    MUX_UNSIGNED #(.width(32)) u_mux_799 (
        .y(_instreth__d),
        .sel(reset),
        .a(32'h0),
        .b(_GEN_81)
    );
    assign io_epc = _mepc__q;
    assign io_evec = _T_560;
    assign io_expt = _T_557;
    assign io_host_tohost = _mtohost__q;
    assign io_out = _T_281;
    assign _mbadaddr__d = _GEN_67;
    assign _mcause__d = _GEN_62;
    BITS #(.width(35), .high(31), .low(0)) bits_800 (
        .y(_mepc__d),
        .in(_GEN_61)
    );
    assign _mfromhost__d = _GEN_77;
    assign _mscratch__d = _GEN_75;
    assign _mtimecmp__d = _GEN_74;
    MUX_UNSIGNED #(.width(32)) u_mux_801 (
        .y(_mtohost__d),
        .sel(reset),
        .a(32'h0),
        .b(_GEN_76)
    );
    MUX_UNSIGNED #(.width(32)) u_mux_802 (
        .y(_time___d),
        .sel(reset),
        .a(32'h0),
        .b(_GEN_72)
    );
    MUX_UNSIGNED #(.width(32)) u_mux_803 (
        .y(_timeh__d),
        .sel(reset),
        .a(32'h0),
        .b(_GEN_73)
    );
endmodule //CSR
module DFF_POSCLK(q, d, clk);
    parameter width = 4;
    output reg [width-1:0] q;
    input [width-1:0] d;
    input clk;
    always @(posedge clk) begin
        q <= d;
    end
endmodule // DFF_POSCLK
module BITS(y, in);
    parameter width = 4;
    parameter high = 2;
    parameter low = 0;
    output [high-low:0] y;
    input [width-1:0] in;
    assign y = in[high:low];
endmodule // BITS
module CAT(y, a, b);
    parameter width_a = 4;
    parameter width_b = 4;
    output [width_a+width_b-1:0] y;
    input [width_a-1:0] a;
    input [width_b-1:0] b;
    assign y = {a, b};
endmodule // CAT
module MUX_UNSIGNED(y, sel, a, b);
    parameter width = 4;
    output [width-1:0] y;
    input sel;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = sel ? a : b;
endmodule // MUX_UNSIGNED
module BITWISEAND(y, a, b);
    parameter width = 4;
    output [width-1:0] y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a & b;
endmodule // BITWISEAND
module EQ_UNSIGNED(y, a, b);
    parameter width = 4;
    output y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a == b;
endmodule // EQ_UNSIGNED
module PAD_UNSIGNED(y, in);
    parameter width = 4;
    parameter n = 4;
    output [(n > width ? n : width)-1:0] y;
    input [width-1:0] in;
    assign y = (n > width) ? {{(n - width){1'b0}}, in} : in;
endmodule // PAD_UNSIGNED
module LEQ_UNSIGNED(y, a, b);
    parameter width = 4;
    output y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a <= b;
endmodule // LEQ_UNSIGNED
module BITWISEOR(y, a, b);
    parameter width = 4;
    output [width-1:0] y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a | b;
endmodule // BITWISEOR
module BITWISENOT(y, in);
    parameter width = 4;
    output [width-1:0] y;
    input [width-1:0] in;
    assign y = ~in;
endmodule // BITWISENOT
module NEQ_UNSIGNED(y, a, b);
    parameter width = 4;
    output y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a != b;
endmodule // NEQ_UNSIGNED
module SHL_UNSIGNED(y, in);
    parameter width = 4;
    parameter n = 4;
    output [width+n-1:0] y;
    input [width-1:0] in;
    wire [width+n-1:0] temp;
    assign temp = {{n{1'b0}}, in};
    assign y = temp << n;
endmodule // SHL_UNSIGNED
module ADD_UNSIGNED(y, a, b);
    parameter width = 4;
    output [width:0] y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a + b;
endmodule // ADD_UNSIGNED
module TAIL(y, in);
    parameter width = 4;
    parameter n = 2;
    output [width-n-1:0] y;
    input [width-1:0] in;
    assign y = in[width-n-1:0];
endmodule // TAIL
module SHR_UNSIGNED(y, in);
    parameter width = 4;
    parameter n = 2;
    output [(n < width ? (width-n-1) : 0):0] y;
    input [width-1:0] in;
    assign y = n < width ? in[width-1:n] : 1'b0;
endmodule // SHR_UNSIGNED
module DSHR_UNSIGNED(y, in, n);
    parameter width_in = 4;
    parameter width_n = 2;
    output [width_in-1:0] y;
    input [width_in-1:0] in;
    input [width_n-1:0] n;
    assign y = in >> n;
endmodule // DSHR_UNSIGNED
module DSHL_UNSIGNED(y, in, n);
    parameter width_in = 4;
    parameter width_n = 2;
    output [(width_in+2**width_n-1)-1:0] y;
    input [width_in-1:0] in;
    input [width_n-1:0] n;
    wire [(width_in+2**width_n-1)-1:0] temp;
    assign temp = {{(2**width_n-1){1'b0}}, in};
    assign y = temp << n;
endmodule // DSHL_UNSIGNED
module RegFile(
    input clock,
    input reset,
    input [4:0] io_raddr1,
    input [4:0] io_raddr2,
    output [31:0] io_rdata1,
    output [31:0] io_rdata2,
    input io_wen,
    input [4:0] io_waddr,
    input [31:0] io_wdata
);
    wire [31:0] regs__T_20_data;
    wire regs__T_20_clk;
    wire regs__T_20_en;
    wire [4:0] regs__T_20_addr;
    wire [31:0] regs__T_25_data;
    wire regs__T_25_clk;
    wire regs__T_25_en;
    wire [4:0] regs__T_25_addr;
    wire regs__T_31_clk;
    wire regs__T_31_en;
    wire regs__T_31_mask;
    wire [4:0] regs__T_31_addr;
    wire [31:0] regs__T_31_data;
    wire [63:0] regs_read_datas;
    wire [1:0] regs_read_clks;
    wire [1:0] regs_read_ens;
    wire [9:0] regs_read_addrs;
    wire regs_write_clks;
    wire regs_write_ens;
    wire regs_write_masks;
    wire [4:0] regs_write_addrs;
    wire [31:0] regs_write_datas;
    BITS #(.width(64), .high(31), .low(0)) bits_804 (
        .y(regs__T_20_data),
        .in(regs_read_datas)
    );
    BITS #(.width(64), .high(63), .low(32)) bits_805 (
        .y(regs__T_25_data),
        .in(regs_read_datas)
    );
    CAT #(.width_a(1), .width_b(1)) cat_806 (
        .y(regs_read_clks),
        .a(regs__T_25_clk),
        .b(regs__T_20_clk)
    );
    CAT #(.width_a(1), .width_b(1)) cat_807 (
        .y(regs_read_ens),
        .a(regs__T_25_en),
        .b(regs__T_20_en)
    );
    CAT #(.width_a(5), .width_b(5)) cat_808 (
        .y(regs_read_addrs),
        .a(regs__T_25_addr),
        .b(regs__T_20_addr)
    );
    assign regs_write_datas = regs__T_31_data;
    assign regs_write_clks = regs__T_31_clk;
    assign regs_write_ens = regs__T_31_en;
    assign regs_write_addrs = regs__T_31_addr;
    assign regs_write_masks = regs__T_31_mask;
    MRMWMEM #(.depth(32), .addrbits(5), .width(32), .readernum(2), .writernum(1), .isSyncRead(0)) regs (
        .read_datas(regs_read_datas),
        .read_clks(regs_read_clks),
        .read_ens(regs_read_ens),
        .read_addrs(regs_read_addrs),
        .write_clks(regs_write_clks),
        .write_ens(regs_write_ens),
        .write_masks(regs_write_masks),
        .write_addrs(regs_write_addrs),
        .write_datas(regs_write_datas)
    );
    wire _T_19;
    wire [4:0] _WTEMP_54;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_809 (
        .y(_WTEMP_54),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(5)) u_neq_810 (
        .y(_T_19),
        .a(io_raddr1),
        .b(_WTEMP_54)
    );
    wire [31:0] _T_22;
    wire [31:0] _WTEMP_55;
    PAD_UNSIGNED #(.width(1), .n(32)) u_pad_811 (
        .y(_WTEMP_55),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(32)) u_mux_812 (
        .y(_T_22),
        .sel(_T_19),
        .a(regs__T_20_data),
        .b(_WTEMP_55)
    );
    wire _T_24;
    wire [4:0] _WTEMP_56;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_813 (
        .y(_WTEMP_56),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(5)) u_neq_814 (
        .y(_T_24),
        .a(io_raddr2),
        .b(_WTEMP_56)
    );
    wire [31:0] _T_27;
    wire [31:0] _WTEMP_57;
    PAD_UNSIGNED #(.width(1), .n(32)) u_pad_815 (
        .y(_WTEMP_57),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(32)) u_mux_816 (
        .y(_T_27),
        .sel(_T_24),
        .a(regs__T_25_data),
        .b(_WTEMP_57)
    );
    wire _T_29;
    wire [4:0] _WTEMP_58;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_817 (
        .y(_WTEMP_58),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(5)) u_neq_818 (
        .y(_T_29),
        .a(io_waddr),
        .b(_WTEMP_58)
    );
    wire _T_30;
    BITWISEAND #(.width(1)) bitwiseand_819 (
        .y(_T_30),
        .a(io_wen),
        .b(_T_29)
    );
    wire [4:0] _GEN_0;
    assign _GEN_0 = io_waddr;
    wire _GEN_1;
    assign _GEN_1 = clock;
    wire _GEN_2;
    MUX_UNSIGNED #(.width(1)) u_mux_820 (
        .y(_GEN_2),
        .sel(_T_30),
        .a(1'h1),
        .b(1'h0)
    );
    wire [31:0] _GEN_3;
    assign _GEN_3 = io_wdata;
    assign io_rdata1 = _T_22;
    assign io_rdata2 = _T_27;
    assign regs__T_20_addr = io_raddr1;
    assign regs__T_20_clk = clock;
    assign regs__T_20_en = 1'h1;
    assign regs__T_25_addr = io_raddr2;
    assign regs__T_25_clk = clock;
    assign regs__T_25_en = 1'h1;
    assign regs__T_31_addr = _GEN_0;
    assign regs__T_31_clk = _GEN_1;
    assign regs__T_31_data = _GEN_3;
    assign regs__T_31_en = _GEN_2;
    assign regs__T_31_mask = _GEN_2;
endmodule //RegFile
module MRMWMEM(read_datas, read_clks, read_ens, read_addrs, write_clks, write_ens, write_masks, write_addrs, write_datas);
    parameter depth = 16;
    parameter addrbits = 4;
    parameter width = 32;
    parameter readernum = 2;
    parameter writernum = 2;
    parameter isSyncRead = 0;
    output [(width*readernum-1):0] read_datas;
    input [(1*readernum-1):0] read_clks;
    input [(1*readernum-1):0] read_ens;
    input [(addrbits*readernum-1):0] read_addrs;
    input [1*writernum-1:0] write_clks;
    input [1*writernum-1:0] write_ens;
    input [1*writernum-1:0] write_masks;
    input [(addrbits*writernum-1):0] write_addrs;
    input [(width*writernum-1):0] write_datas;
    reg [width-1:0] memcore [0:depth-1];
    wire [(addrbits*readernum-1):0] final_read_addrs;
    genvar gv_n;
    generate
        for (gv_n = 0; gv_n < readernum; gv_n = gv_n + 1) begin: get_final_raddrs
            if (isSyncRead) begin: raddr_processor
                reg [addrbits-1:0] read_addr_pipe_0;
                always @(posedge read_clks[gv_n]) begin
                    if (read_ens[gv_n]) begin
                        read_addr_pipe_0 <= read_addrs[gv_n*addrbits +: addrbits];
                    end
                end
                assign final_read_addrs[gv_n*addrbits +: addrbits] = read_addr_pipe_0;
            end else begin: raddr_processor
                assign final_read_addrs[gv_n*addrbits +: addrbits] = read_addrs[gv_n*addrbits +: addrbits];
            end
        end
    endgenerate
    genvar gv_k;
    generate
        for (gv_k = 0; gv_k < readernum; gv_k = gv_k + 1) begin: form_read_datas
            assign read_datas[gv_k*width +: width] = memcore[final_read_addrs[gv_k*addrbits +: addrbits]];
        end
    endgenerate
    integer i;
    always @(posedge write_clks[0]) begin
        for (i = 0; i < writernum; i = i + 1) begin
            if (write_ens[i] & write_masks[i]) begin
                memcore[write_addrs[i*addrbits +: addrbits]] <= write_datas[i*width +: width];
            end
        end
    end
endmodule // MRMWMEM
module ALUArea(
    input clock,
    input reset,
    input [31:0] io_A,
    input [31:0] io_B,
    input [3:0] io_alu_op,
    output [31:0] io_out,
    output [31:0] io_sum
);
    wire _T_12;
    BITS #(.width(4), .high(0), .low(0)) bits_821 (
        .y(_T_12),
        .in(io_alu_op)
    );
    wire [32:0] _T_14;
    wire [31:0] _WTEMP_59;
    PAD_UNSIGNED #(.width(1), .n(32)) u_pad_822 (
        .y(_WTEMP_59),
        .in(1'h0)
    );
    SUB_UNSIGNED #(.width(32)) u_sub_823 (
        .y(_T_14),
        .a(_WTEMP_59),
        .b(io_B)
    );
    wire [31:0] _T_15;
    TAIL #(.width(33), .n(1)) tail_824 (
        .y(_T_15),
        .in(_T_14)
    );
    wire [31:0] _T_16;
    MUX_UNSIGNED #(.width(32)) u_mux_825 (
        .y(_T_16),
        .sel(_T_12),
        .a(_T_15),
        .b(io_B)
    );
    wire [32:0] _T_17;
    ADD_UNSIGNED #(.width(32)) u_add_826 (
        .y(_T_17),
        .a(io_A),
        .b(_T_16)
    );
    wire [31:0] sum;
    TAIL #(.width(33), .n(1)) tail_827 (
        .y(sum),
        .in(_T_17)
    );
    wire _T_18;
    BITS #(.width(32), .high(31), .low(31)) bits_828 (
        .y(_T_18),
        .in(io_A)
    );
    wire _T_19;
    BITS #(.width(32), .high(31), .low(31)) bits_829 (
        .y(_T_19),
        .in(io_B)
    );
    wire _T_20;
    EQ_UNSIGNED #(.width(1)) u_eq_830 (
        .y(_T_20),
        .a(_T_18),
        .b(_T_19)
    );
    wire _T_21;
    BITS #(.width(32), .high(31), .low(31)) bits_831 (
        .y(_T_21),
        .in(sum)
    );
    wire _T_22;
    BITS #(.width(4), .high(1), .low(1)) bits_832 (
        .y(_T_22),
        .in(io_alu_op)
    );
    wire _T_23;
    BITS #(.width(32), .high(31), .low(31)) bits_833 (
        .y(_T_23),
        .in(io_B)
    );
    wire _T_24;
    BITS #(.width(32), .high(31), .low(31)) bits_834 (
        .y(_T_24),
        .in(io_A)
    );
    wire _T_25;
    MUX_UNSIGNED #(.width(1)) u_mux_835 (
        .y(_T_25),
        .sel(_T_22),
        .a(_T_23),
        .b(_T_24)
    );
    wire cmp;
    MUX_UNSIGNED #(.width(1)) u_mux_836 (
        .y(cmp),
        .sel(_T_20),
        .a(_T_21),
        .b(_T_25)
    );
    wire [4:0] shamt;
    BITS #(.width(32), .high(4), .low(0)) bits_837 (
        .y(shamt),
        .in(io_B)
    );
    wire _T_26;
    BITS #(.width(4), .high(3), .low(3)) bits_838 (
        .y(_T_26),
        .in(io_alu_op)
    );
    wire [31:0] _T_29;
    assign _T_29 = 32'hFFFF0000;
    wire [31:0] _T_30;
    assign _T_30 = 32'hFFFF;
    wire [15:0] _T_31;
    SHR_UNSIGNED #(.width(32), .n(16)) u_shr_839 (
        .y(_T_31),
        .in(io_A)
    );
    wire [31:0] _T_32;
    wire [31:0] _WTEMP_60;
    PAD_UNSIGNED #(.width(16), .n(32)) u_pad_840 (
        .y(_WTEMP_60),
        .in(_T_31)
    );
    BITWISEAND #(.width(32)) bitwiseand_841 (
        .y(_T_32),
        .a(_WTEMP_60),
        .b(_T_30)
    );
    wire [15:0] _T_33;
    BITS #(.width(32), .high(15), .low(0)) bits_842 (
        .y(_T_33),
        .in(io_A)
    );
    wire [31:0] _T_34;
    SHL_UNSIGNED #(.width(16), .n(16)) u_shl_843 (
        .y(_T_34),
        .in(_T_33)
    );
    wire [31:0] _T_35;
    assign _T_35 = 32'hFFFF0000;
    wire [31:0] _T_36;
    BITWISEAND #(.width(32)) bitwiseand_844 (
        .y(_T_36),
        .a(_T_34),
        .b(_T_35)
    );
    wire [31:0] _T_37;
    BITWISEOR #(.width(32)) bitwiseor_845 (
        .y(_T_37),
        .a(_T_32),
        .b(_T_36)
    );
    wire [23:0] _T_38;
    assign _T_38 = 24'hFFFF;
    wire [31:0] _T_39;
    assign _T_39 = 32'hFFFF00;
    wire [31:0] _T_40;
    assign _T_40 = 32'hFF00FF;
    wire [23:0] _T_41;
    SHR_UNSIGNED #(.width(32), .n(8)) u_shr_846 (
        .y(_T_41),
        .in(_T_37)
    );
    wire [31:0] _T_42;
    wire [31:0] _WTEMP_61;
    PAD_UNSIGNED #(.width(24), .n(32)) u_pad_847 (
        .y(_WTEMP_61),
        .in(_T_41)
    );
    BITWISEAND #(.width(32)) bitwiseand_848 (
        .y(_T_42),
        .a(_WTEMP_61),
        .b(_T_40)
    );
    wire [23:0] _T_43;
    BITS #(.width(32), .high(23), .low(0)) bits_849 (
        .y(_T_43),
        .in(_T_37)
    );
    wire [31:0] _T_44;
    SHL_UNSIGNED #(.width(24), .n(8)) u_shl_850 (
        .y(_T_44),
        .in(_T_43)
    );
    wire [31:0] _T_45;
    assign _T_45 = 32'hFF00FF00;
    wire [31:0] _T_46;
    BITWISEAND #(.width(32)) bitwiseand_851 (
        .y(_T_46),
        .a(_T_44),
        .b(_T_45)
    );
    wire [31:0] _T_47;
    BITWISEOR #(.width(32)) bitwiseor_852 (
        .y(_T_47),
        .a(_T_42),
        .b(_T_46)
    );
    wire [27:0] _T_48;
    assign _T_48 = 28'hFF00FF;
    wire [31:0] _T_49;
    assign _T_49 = 32'hFF00FF0;
    wire [31:0] _T_50;
    assign _T_50 = 32'hF0F0F0F;
    wire [27:0] _T_51;
    SHR_UNSIGNED #(.width(32), .n(4)) u_shr_853 (
        .y(_T_51),
        .in(_T_47)
    );
    wire [31:0] _T_52;
    wire [31:0] _WTEMP_62;
    PAD_UNSIGNED #(.width(28), .n(32)) u_pad_854 (
        .y(_WTEMP_62),
        .in(_T_51)
    );
    BITWISEAND #(.width(32)) bitwiseand_855 (
        .y(_T_52),
        .a(_WTEMP_62),
        .b(_T_50)
    );
    wire [27:0] _T_53;
    BITS #(.width(32), .high(27), .low(0)) bits_856 (
        .y(_T_53),
        .in(_T_47)
    );
    wire [31:0] _T_54;
    SHL_UNSIGNED #(.width(28), .n(4)) u_shl_857 (
        .y(_T_54),
        .in(_T_53)
    );
    wire [31:0] _T_55;
    assign _T_55 = 32'hF0F0F0F0;
    wire [31:0] _T_56;
    BITWISEAND #(.width(32)) bitwiseand_858 (
        .y(_T_56),
        .a(_T_54),
        .b(_T_55)
    );
    wire [31:0] _T_57;
    BITWISEOR #(.width(32)) bitwiseor_859 (
        .y(_T_57),
        .a(_T_52),
        .b(_T_56)
    );
    wire [29:0] _T_58;
    assign _T_58 = 30'hF0F0F0F;
    wire [31:0] _T_59;
    assign _T_59 = 32'h3C3C3C3C;
    wire [31:0] _T_60;
    assign _T_60 = 32'h33333333;
    wire [29:0] _T_61;
    SHR_UNSIGNED #(.width(32), .n(2)) u_shr_860 (
        .y(_T_61),
        .in(_T_57)
    );
    wire [31:0] _T_62;
    wire [31:0] _WTEMP_63;
    PAD_UNSIGNED #(.width(30), .n(32)) u_pad_861 (
        .y(_WTEMP_63),
        .in(_T_61)
    );
    BITWISEAND #(.width(32)) bitwiseand_862 (
        .y(_T_62),
        .a(_WTEMP_63),
        .b(_T_60)
    );
    wire [29:0] _T_63;
    BITS #(.width(32), .high(29), .low(0)) bits_863 (
        .y(_T_63),
        .in(_T_57)
    );
    wire [31:0] _T_64;
    SHL_UNSIGNED #(.width(30), .n(2)) u_shl_864 (
        .y(_T_64),
        .in(_T_63)
    );
    wire [31:0] _T_65;
    assign _T_65 = 32'hCCCCCCCC;
    wire [31:0] _T_66;
    BITWISEAND #(.width(32)) bitwiseand_865 (
        .y(_T_66),
        .a(_T_64),
        .b(_T_65)
    );
    wire [31:0] _T_67;
    BITWISEOR #(.width(32)) bitwiseor_866 (
        .y(_T_67),
        .a(_T_62),
        .b(_T_66)
    );
    wire [30:0] _T_68;
    assign _T_68 = 31'h33333333;
    wire [31:0] _T_69;
    assign _T_69 = 32'h66666666;
    wire [31:0] _T_70;
    assign _T_70 = 32'h55555555;
    wire [30:0] _T_71;
    SHR_UNSIGNED #(.width(32), .n(1)) u_shr_867 (
        .y(_T_71),
        .in(_T_67)
    );
    wire [31:0] _T_72;
    wire [31:0] _WTEMP_64;
    PAD_UNSIGNED #(.width(31), .n(32)) u_pad_868 (
        .y(_WTEMP_64),
        .in(_T_71)
    );
    BITWISEAND #(.width(32)) bitwiseand_869 (
        .y(_T_72),
        .a(_WTEMP_64),
        .b(_T_70)
    );
    wire [30:0] _T_73;
    BITS #(.width(32), .high(30), .low(0)) bits_870 (
        .y(_T_73),
        .in(_T_67)
    );
    wire [31:0] _T_74;
    SHL_UNSIGNED #(.width(31), .n(1)) u_shl_871 (
        .y(_T_74),
        .in(_T_73)
    );
    wire [31:0] _T_75;
    assign _T_75 = 32'hAAAAAAAA;
    wire [31:0] _T_76;
    BITWISEAND #(.width(32)) bitwiseand_872 (
        .y(_T_76),
        .a(_T_74),
        .b(_T_75)
    );
    wire [31:0] _T_77;
    BITWISEOR #(.width(32)) bitwiseor_873 (
        .y(_T_77),
        .a(_T_72),
        .b(_T_76)
    );
    wire [31:0] shin;
    MUX_UNSIGNED #(.width(32)) u_mux_874 (
        .y(shin),
        .sel(_T_26),
        .a(io_A),
        .b(_T_77)
    );
    wire _T_78;
    BITS #(.width(4), .high(0), .low(0)) bits_875 (
        .y(_T_78),
        .in(io_alu_op)
    );
    wire _T_79;
    BITS #(.width(32), .high(31), .low(31)) bits_876 (
        .y(_T_79),
        .in(shin)
    );
    wire _T_80;
    BITWISEAND #(.width(1)) bitwiseand_877 (
        .y(_T_80),
        .a(_T_78),
        .b(_T_79)
    );
    wire [32:0] _T_81;
    CAT #(.width_a(1), .width_b(32)) cat_878 (
        .y(_T_81),
        .a(_T_80),
        .b(shin)
    );
    wire [32:0] _T_82;
    ASSINT #(.width(33)) assint_879 (
        .y(_T_82),
        .in(_T_81)
    );
    wire [32:0] _T_83;
    DSHR_SIGNED #(.width_in(33), .width_n(5)) s_dshr_880 (
        .y(_T_83),
        .in(_T_82),
        .n(shamt)
    );
    wire [31:0] shiftr;
    BITS #(.width(33), .high(31), .low(0)) bits_881 (
        .y(shiftr),
        .in(_T_83)
    );
    wire [31:0] _T_86;
    assign _T_86 = 32'hFFFF0000;
    wire [31:0] _T_87;
    assign _T_87 = 32'hFFFF;
    wire [15:0] _T_88;
    SHR_UNSIGNED #(.width(32), .n(16)) u_shr_882 (
        .y(_T_88),
        .in(shiftr)
    );
    wire [31:0] _T_89;
    wire [31:0] _WTEMP_65;
    PAD_UNSIGNED #(.width(16), .n(32)) u_pad_883 (
        .y(_WTEMP_65),
        .in(_T_88)
    );
    BITWISEAND #(.width(32)) bitwiseand_884 (
        .y(_T_89),
        .a(_WTEMP_65),
        .b(_T_87)
    );
    wire [15:0] _T_90;
    BITS #(.width(32), .high(15), .low(0)) bits_885 (
        .y(_T_90),
        .in(shiftr)
    );
    wire [31:0] _T_91;
    SHL_UNSIGNED #(.width(16), .n(16)) u_shl_886 (
        .y(_T_91),
        .in(_T_90)
    );
    wire [31:0] _T_92;
    assign _T_92 = 32'hFFFF0000;
    wire [31:0] _T_93;
    BITWISEAND #(.width(32)) bitwiseand_887 (
        .y(_T_93),
        .a(_T_91),
        .b(_T_92)
    );
    wire [31:0] _T_94;
    BITWISEOR #(.width(32)) bitwiseor_888 (
        .y(_T_94),
        .a(_T_89),
        .b(_T_93)
    );
    wire [23:0] _T_95;
    assign _T_95 = 24'hFFFF;
    wire [31:0] _T_96;
    assign _T_96 = 32'hFFFF00;
    wire [31:0] _T_97;
    assign _T_97 = 32'hFF00FF;
    wire [23:0] _T_98;
    SHR_UNSIGNED #(.width(32), .n(8)) u_shr_889 (
        .y(_T_98),
        .in(_T_94)
    );
    wire [31:0] _T_99;
    wire [31:0] _WTEMP_66;
    PAD_UNSIGNED #(.width(24), .n(32)) u_pad_890 (
        .y(_WTEMP_66),
        .in(_T_98)
    );
    BITWISEAND #(.width(32)) bitwiseand_891 (
        .y(_T_99),
        .a(_WTEMP_66),
        .b(_T_97)
    );
    wire [23:0] _T_100;
    BITS #(.width(32), .high(23), .low(0)) bits_892 (
        .y(_T_100),
        .in(_T_94)
    );
    wire [31:0] _T_101;
    SHL_UNSIGNED #(.width(24), .n(8)) u_shl_893 (
        .y(_T_101),
        .in(_T_100)
    );
    wire [31:0] _T_102;
    assign _T_102 = 32'hFF00FF00;
    wire [31:0] _T_103;
    BITWISEAND #(.width(32)) bitwiseand_894 (
        .y(_T_103),
        .a(_T_101),
        .b(_T_102)
    );
    wire [31:0] _T_104;
    BITWISEOR #(.width(32)) bitwiseor_895 (
        .y(_T_104),
        .a(_T_99),
        .b(_T_103)
    );
    wire [27:0] _T_105;
    assign _T_105 = 28'hFF00FF;
    wire [31:0] _T_106;
    assign _T_106 = 32'hFF00FF0;
    wire [31:0] _T_107;
    assign _T_107 = 32'hF0F0F0F;
    wire [27:0] _T_108;
    SHR_UNSIGNED #(.width(32), .n(4)) u_shr_896 (
        .y(_T_108),
        .in(_T_104)
    );
    wire [31:0] _T_109;
    wire [31:0] _WTEMP_67;
    PAD_UNSIGNED #(.width(28), .n(32)) u_pad_897 (
        .y(_WTEMP_67),
        .in(_T_108)
    );
    BITWISEAND #(.width(32)) bitwiseand_898 (
        .y(_T_109),
        .a(_WTEMP_67),
        .b(_T_107)
    );
    wire [27:0] _T_110;
    BITS #(.width(32), .high(27), .low(0)) bits_899 (
        .y(_T_110),
        .in(_T_104)
    );
    wire [31:0] _T_111;
    SHL_UNSIGNED #(.width(28), .n(4)) u_shl_900 (
        .y(_T_111),
        .in(_T_110)
    );
    wire [31:0] _T_112;
    assign _T_112 = 32'hF0F0F0F0;
    wire [31:0] _T_113;
    BITWISEAND #(.width(32)) bitwiseand_901 (
        .y(_T_113),
        .a(_T_111),
        .b(_T_112)
    );
    wire [31:0] _T_114;
    BITWISEOR #(.width(32)) bitwiseor_902 (
        .y(_T_114),
        .a(_T_109),
        .b(_T_113)
    );
    wire [29:0] _T_115;
    assign _T_115 = 30'hF0F0F0F;
    wire [31:0] _T_116;
    assign _T_116 = 32'h3C3C3C3C;
    wire [31:0] _T_117;
    assign _T_117 = 32'h33333333;
    wire [29:0] _T_118;
    SHR_UNSIGNED #(.width(32), .n(2)) u_shr_903 (
        .y(_T_118),
        .in(_T_114)
    );
    wire [31:0] _T_119;
    wire [31:0] _WTEMP_68;
    PAD_UNSIGNED #(.width(30), .n(32)) u_pad_904 (
        .y(_WTEMP_68),
        .in(_T_118)
    );
    BITWISEAND #(.width(32)) bitwiseand_905 (
        .y(_T_119),
        .a(_WTEMP_68),
        .b(_T_117)
    );
    wire [29:0] _T_120;
    BITS #(.width(32), .high(29), .low(0)) bits_906 (
        .y(_T_120),
        .in(_T_114)
    );
    wire [31:0] _T_121;
    SHL_UNSIGNED #(.width(30), .n(2)) u_shl_907 (
        .y(_T_121),
        .in(_T_120)
    );
    wire [31:0] _T_122;
    assign _T_122 = 32'hCCCCCCCC;
    wire [31:0] _T_123;
    BITWISEAND #(.width(32)) bitwiseand_908 (
        .y(_T_123),
        .a(_T_121),
        .b(_T_122)
    );
    wire [31:0] _T_124;
    BITWISEOR #(.width(32)) bitwiseor_909 (
        .y(_T_124),
        .a(_T_119),
        .b(_T_123)
    );
    wire [30:0] _T_125;
    assign _T_125 = 31'h33333333;
    wire [31:0] _T_126;
    assign _T_126 = 32'h66666666;
    wire [31:0] _T_127;
    assign _T_127 = 32'h55555555;
    wire [30:0] _T_128;
    SHR_UNSIGNED #(.width(32), .n(1)) u_shr_910 (
        .y(_T_128),
        .in(_T_124)
    );
    wire [31:0] _T_129;
    wire [31:0] _WTEMP_69;
    PAD_UNSIGNED #(.width(31), .n(32)) u_pad_911 (
        .y(_WTEMP_69),
        .in(_T_128)
    );
    BITWISEAND #(.width(32)) bitwiseand_912 (
        .y(_T_129),
        .a(_WTEMP_69),
        .b(_T_127)
    );
    wire [30:0] _T_130;
    BITS #(.width(32), .high(30), .low(0)) bits_913 (
        .y(_T_130),
        .in(_T_124)
    );
    wire [31:0] _T_131;
    SHL_UNSIGNED #(.width(31), .n(1)) u_shl_914 (
        .y(_T_131),
        .in(_T_130)
    );
    wire [31:0] _T_132;
    assign _T_132 = 32'hAAAAAAAA;
    wire [31:0] _T_133;
    BITWISEAND #(.width(32)) bitwiseand_915 (
        .y(_T_133),
        .a(_T_131),
        .b(_T_132)
    );
    wire [31:0] shiftl;
    BITWISEOR #(.width(32)) bitwiseor_916 (
        .y(shiftl),
        .a(_T_129),
        .b(_T_133)
    );
    wire _T_134;
    EQ_UNSIGNED #(.width(4)) u_eq_917 (
        .y(_T_134),
        .a(io_alu_op),
        .b(4'h0)
    );
    wire _T_135;
    EQ_UNSIGNED #(.width(4)) u_eq_918 (
        .y(_T_135),
        .a(io_alu_op),
        .b(4'h1)
    );
    wire _T_136;
    BITWISEOR #(.width(1)) bitwiseor_919 (
        .y(_T_136),
        .a(_T_134),
        .b(_T_135)
    );
    wire _T_137;
    EQ_UNSIGNED #(.width(4)) u_eq_920 (
        .y(_T_137),
        .a(io_alu_op),
        .b(4'h5)
    );
    wire _T_138;
    EQ_UNSIGNED #(.width(4)) u_eq_921 (
        .y(_T_138),
        .a(io_alu_op),
        .b(4'h7)
    );
    wire _T_139;
    BITWISEOR #(.width(1)) bitwiseor_922 (
        .y(_T_139),
        .a(_T_137),
        .b(_T_138)
    );
    wire _T_140;
    EQ_UNSIGNED #(.width(4)) u_eq_923 (
        .y(_T_140),
        .a(io_alu_op),
        .b(4'h9)
    );
    wire _T_141;
    EQ_UNSIGNED #(.width(4)) u_eq_924 (
        .y(_T_141),
        .a(io_alu_op),
        .b(4'h8)
    );
    wire _T_142;
    BITWISEOR #(.width(1)) bitwiseor_925 (
        .y(_T_142),
        .a(_T_140),
        .b(_T_141)
    );
    wire _T_143;
    EQ_UNSIGNED #(.width(4)) u_eq_926 (
        .y(_T_143),
        .a(io_alu_op),
        .b(4'h6)
    );
    wire _T_144;
    EQ_UNSIGNED #(.width(4)) u_eq_927 (
        .y(_T_144),
        .a(io_alu_op),
        .b(4'h2)
    );
    wire [31:0] _T_145;
    BITWISEAND #(.width(32)) bitwiseand_928 (
        .y(_T_145),
        .a(io_A),
        .b(io_B)
    );
    wire _T_146;
    EQ_UNSIGNED #(.width(4)) u_eq_929 (
        .y(_T_146),
        .a(io_alu_op),
        .b(4'h3)
    );
    wire [31:0] _T_147;
    BITWISEOR #(.width(32)) bitwiseor_930 (
        .y(_T_147),
        .a(io_A),
        .b(io_B)
    );
    wire _T_148;
    EQ_UNSIGNED #(.width(4)) u_eq_931 (
        .y(_T_148),
        .a(io_alu_op),
        .b(4'h4)
    );
    wire [31:0] _T_149;
    BITWISEXOR #(.width(32)) bitwisexor_932 (
        .y(_T_149),
        .a(io_A),
        .b(io_B)
    );
    wire _T_150;
    EQ_UNSIGNED #(.width(4)) u_eq_933 (
        .y(_T_150),
        .a(io_alu_op),
        .b(4'hA)
    );
    wire [31:0] _T_151;
    MUX_UNSIGNED #(.width(32)) u_mux_934 (
        .y(_T_151),
        .sel(_T_150),
        .a(io_A),
        .b(io_B)
    );
    wire [31:0] _T_152;
    MUX_UNSIGNED #(.width(32)) u_mux_935 (
        .y(_T_152),
        .sel(_T_148),
        .a(_T_149),
        .b(_T_151)
    );
    wire [31:0] _T_153;
    MUX_UNSIGNED #(.width(32)) u_mux_936 (
        .y(_T_153),
        .sel(_T_146),
        .a(_T_147),
        .b(_T_152)
    );
    wire [31:0] _T_154;
    MUX_UNSIGNED #(.width(32)) u_mux_937 (
        .y(_T_154),
        .sel(_T_144),
        .a(_T_145),
        .b(_T_153)
    );
    wire [31:0] _T_155;
    MUX_UNSIGNED #(.width(32)) u_mux_938 (
        .y(_T_155),
        .sel(_T_143),
        .a(shiftl),
        .b(_T_154)
    );
    wire [31:0] _T_156;
    MUX_UNSIGNED #(.width(32)) u_mux_939 (
        .y(_T_156),
        .sel(_T_142),
        .a(shiftr),
        .b(_T_155)
    );
    wire _T_157;
    SHL_UNSIGNED #(.width(1), .n(0)) u_shl_940 (
        .y(_T_157),
        .in(cmp)
    );
    wire [31:0] _T_158;
    wire [31:0] _WTEMP_70;
    PAD_UNSIGNED #(.width(1), .n(32)) u_pad_941 (
        .y(_WTEMP_70),
        .in(_T_157)
    );
    MUX_UNSIGNED #(.width(32)) u_mux_942 (
        .y(_T_158),
        .sel(_T_139),
        .a(_WTEMP_70),
        .b(_T_156)
    );
    wire [31:0] out;
    MUX_UNSIGNED #(.width(32)) u_mux_943 (
        .y(out),
        .sel(_T_136),
        .a(sum),
        .b(_T_158)
    );
    assign io_out = out;
    assign io_sum = sum;
endmodule //ALUArea
module SUB_UNSIGNED(y, a, b);
    parameter width = 4;
    output [width:0] y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a - b;
endmodule // SUB_UNSIGNED
module ASSINT(y, in);
    parameter width = 4;
    output [width-1:0] y;
    input [width-1:0] in;
    assign y = $signed(in);
endmodule // ASSINT
module DSHR_SIGNED(y, in, n);
    parameter width_in = 4;
    parameter width_n = 2;
    output [width_in-1:0] y;
    input [width_in-1:0] in;
    input [width_n-1:0] n;
    assign y = $signed(in) >>> n;
endmodule // DSHR_SIGNED
module BITWISEXOR(y, a, b);
    parameter width = 4;
    output [width-1:0] y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a ^ b;
endmodule // BITWISEXOR
module ImmGenWire(
    input clock,
    input reset,
    input [31:0] io_inst,
    input [2:0] io_sel,
    output [31:0] io_out
);
    wire [11:0] _T_8;
    BITS #(.width(32), .high(31), .low(20)) bits_944 (
        .y(_T_8),
        .in(io_inst)
    );
    wire [11:0] Iimm;
    ASSINT #(.width(12)) assint_945 (
        .y(Iimm),
        .in(_T_8)
    );
    wire [6:0] _T_9;
    BITS #(.width(32), .high(31), .low(25)) bits_946 (
        .y(_T_9),
        .in(io_inst)
    );
    wire [4:0] _T_10;
    BITS #(.width(32), .high(11), .low(7)) bits_947 (
        .y(_T_10),
        .in(io_inst)
    );
    wire [11:0] _T_11;
    CAT #(.width_a(7), .width_b(5)) cat_948 (
        .y(_T_11),
        .a(_T_9),
        .b(_T_10)
    );
    wire [11:0] Simm;
    ASSINT #(.width(12)) assint_949 (
        .y(Simm),
        .in(_T_11)
    );
    wire _T_12;
    BITS #(.width(32), .high(31), .low(31)) bits_950 (
        .y(_T_12),
        .in(io_inst)
    );
    wire _T_13;
    BITS #(.width(32), .high(7), .low(7)) bits_951 (
        .y(_T_13),
        .in(io_inst)
    );
    wire [5:0] _T_14;
    BITS #(.width(32), .high(30), .low(25)) bits_952 (
        .y(_T_14),
        .in(io_inst)
    );
    wire [3:0] _T_15;
    BITS #(.width(32), .high(11), .low(8)) bits_953 (
        .y(_T_15),
        .in(io_inst)
    );
    wire [4:0] _T_17;
    CAT #(.width_a(4), .width_b(1)) cat_954 (
        .y(_T_17),
        .a(_T_15),
        .b(1'h0)
    );
    wire [1:0] _T_18;
    CAT #(.width_a(1), .width_b(1)) cat_955 (
        .y(_T_18),
        .a(_T_12),
        .b(_T_13)
    );
    wire [7:0] _T_19;
    CAT #(.width_a(2), .width_b(6)) cat_956 (
        .y(_T_19),
        .a(_T_18),
        .b(_T_14)
    );
    wire [12:0] _T_20;
    CAT #(.width_a(8), .width_b(5)) cat_957 (
        .y(_T_20),
        .a(_T_19),
        .b(_T_17)
    );
    wire [12:0] Bimm;
    ASSINT #(.width(13)) assint_958 (
        .y(Bimm),
        .in(_T_20)
    );
    wire [19:0] _T_21;
    BITS #(.width(32), .high(31), .low(12)) bits_959 (
        .y(_T_21),
        .in(io_inst)
    );
    wire [31:0] _T_23;
    CAT #(.width_a(20), .width_b(12)) cat_960 (
        .y(_T_23),
        .a(_T_21),
        .b(12'h0)
    );
    wire [31:0] Uimm;
    ASSINT #(.width(32)) assint_961 (
        .y(Uimm),
        .in(_T_23)
    );
    wire _T_24;
    BITS #(.width(32), .high(31), .low(31)) bits_962 (
        .y(_T_24),
        .in(io_inst)
    );
    wire [7:0] _T_25;
    BITS #(.width(32), .high(19), .low(12)) bits_963 (
        .y(_T_25),
        .in(io_inst)
    );
    wire _T_26;
    BITS #(.width(32), .high(20), .low(20)) bits_964 (
        .y(_T_26),
        .in(io_inst)
    );
    wire [5:0] _T_27;
    BITS #(.width(32), .high(30), .low(25)) bits_965 (
        .y(_T_27),
        .in(io_inst)
    );
    wire [3:0] _T_28;
    BITS #(.width(32), .high(24), .low(21)) bits_966 (
        .y(_T_28),
        .in(io_inst)
    );
    wire [9:0] _T_30;
    CAT #(.width_a(6), .width_b(4)) cat_967 (
        .y(_T_30),
        .a(_T_27),
        .b(_T_28)
    );
    wire [10:0] _T_31;
    CAT #(.width_a(10), .width_b(1)) cat_968 (
        .y(_T_31),
        .a(_T_30),
        .b(1'h0)
    );
    wire [8:0] _T_32;
    CAT #(.width_a(1), .width_b(8)) cat_969 (
        .y(_T_32),
        .a(_T_24),
        .b(_T_25)
    );
    wire [9:0] _T_33;
    CAT #(.width_a(9), .width_b(1)) cat_970 (
        .y(_T_33),
        .a(_T_32),
        .b(_T_26)
    );
    wire [20:0] _T_34;
    CAT #(.width_a(10), .width_b(11)) cat_971 (
        .y(_T_34),
        .a(_T_33),
        .b(_T_31)
    );
    wire [20:0] Jimm;
    ASSINT #(.width(21)) assint_972 (
        .y(Jimm),
        .in(_T_34)
    );
    wire [4:0] _T_35;
    BITS #(.width(32), .high(19), .low(15)) bits_973 (
        .y(_T_35),
        .in(io_inst)
    );
    wire [5:0] Zimm;
    CVT_UNSIGNED #(.width(5)) u_cvt_974 (
        .y(Zimm),
        .in(_T_35)
    );
    wire [11:0] _T_37;
    wire [11:0] _WTEMP_71;
    PAD_SIGNED #(.width(2), .n(12)) s_pad_975 (
        .y(_WTEMP_71),
        .in(-2'sh2)
    );
    BITWISEAND #(.width(12)) bitwiseand_976 (
        .y(_T_37),
        .a(Iimm),
        .b(_WTEMP_71)
    );
    wire [11:0] _T_38;
    ASSINT #(.width(12)) assint_977 (
        .y(_T_38),
        .in(_T_37)
    );
    wire _T_39;
    EQ_UNSIGNED #(.width(3)) u_eq_978 (
        .y(_T_39),
        .a(3'h6),
        .b(io_sel)
    );
    wire [11:0] _T_40;
    wire [11:0] _WTEMP_72;
    PAD_SIGNED #(.width(6), .n(12)) s_pad_979 (
        .y(_WTEMP_72),
        .in(Zimm)
    );
    MUX_SIGNED #(.width(12)) s_mux_980 (
        .y(_T_40),
        .sel(_T_39),
        .a(_WTEMP_72),
        .b(_T_38)
    );
    wire _T_41;
    EQ_UNSIGNED #(.width(3)) u_eq_981 (
        .y(_T_41),
        .a(3'h4),
        .b(io_sel)
    );
    wire [20:0] _T_42;
    wire [20:0] _WTEMP_73;
    PAD_SIGNED #(.width(12), .n(21)) s_pad_982 (
        .y(_WTEMP_73),
        .in(_T_40)
    );
    MUX_SIGNED #(.width(21)) s_mux_983 (
        .y(_T_42),
        .sel(_T_41),
        .a(Jimm),
        .b(_WTEMP_73)
    );
    wire _T_43;
    EQ_UNSIGNED #(.width(3)) u_eq_984 (
        .y(_T_43),
        .a(3'h3),
        .b(io_sel)
    );
    wire [31:0] _T_44;
    wire [31:0] _WTEMP_74;
    PAD_SIGNED #(.width(21), .n(32)) s_pad_985 (
        .y(_WTEMP_74),
        .in(_T_42)
    );
    MUX_SIGNED #(.width(32)) s_mux_986 (
        .y(_T_44),
        .sel(_T_43),
        .a(Uimm),
        .b(_WTEMP_74)
    );
    wire _T_45;
    EQ_UNSIGNED #(.width(3)) u_eq_987 (
        .y(_T_45),
        .a(3'h5),
        .b(io_sel)
    );
    wire [31:0] _T_46;
    wire [31:0] _WTEMP_75;
    PAD_SIGNED #(.width(13), .n(32)) s_pad_988 (
        .y(_WTEMP_75),
        .in(Bimm)
    );
    MUX_SIGNED #(.width(32)) s_mux_989 (
        .y(_T_46),
        .sel(_T_45),
        .a(_WTEMP_75),
        .b(_T_44)
    );
    wire _T_47;
    EQ_UNSIGNED #(.width(3)) u_eq_990 (
        .y(_T_47),
        .a(3'h2),
        .b(io_sel)
    );
    wire [31:0] _T_48;
    wire [31:0] _WTEMP_76;
    PAD_SIGNED #(.width(12), .n(32)) s_pad_991 (
        .y(_WTEMP_76),
        .in(Simm)
    );
    MUX_SIGNED #(.width(32)) s_mux_992 (
        .y(_T_48),
        .sel(_T_47),
        .a(_WTEMP_76),
        .b(_T_46)
    );
    wire _T_49;
    EQ_UNSIGNED #(.width(3)) u_eq_993 (
        .y(_T_49),
        .a(3'h1),
        .b(io_sel)
    );
    wire [31:0] _T_50;
    wire [31:0] _WTEMP_77;
    PAD_SIGNED #(.width(12), .n(32)) s_pad_994 (
        .y(_WTEMP_77),
        .in(Iimm)
    );
    MUX_SIGNED #(.width(32)) s_mux_995 (
        .y(_T_50),
        .sel(_T_49),
        .a(_WTEMP_77),
        .b(_T_48)
    );
    wire [31:0] _T_51;
    ASUINT #(.width(32)) asuint_996 (
        .y(_T_51),
        .in(_T_50)
    );
    assign io_out = _T_51;
endmodule //ImmGenWire
module CVT_UNSIGNED(y, in);
    parameter width = 4;
    output [width:0] y;
    input [width-1:0] in;
    assign y = $signed({1'b0, in});
endmodule // CVT_UNSIGNED
module PAD_SIGNED(y, in);
    parameter width = 4;
    parameter n = 4;
    output [(n > width ? n : width)-1:0] y;
    input [width-1:0] in;
    assign y = n > width ? {{(n - width){in[width-1]}}, in} : in;
endmodule // PAD_SIGNED
module MUX_SIGNED(y, sel, a, b);
    parameter width = 4;
    output [width-1:0] y;
    input sel;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = sel ? $signed(a) : $signed(b);
endmodule // MUX_SIGNED
module ASUINT(y, in);
    parameter width = 4;
    output [width-1:0] y;
    input [width-1:0] in;
    assign y = $unsigned(in);
endmodule // ASUINT
module BrCondArea(
    input clock,
    input reset,
    input [31:0] io_rs1,
    input [31:0] io_rs2,
    input [2:0] io_br_type,
    output io_taken
);
    wire [32:0] _T_10;
    SUB_UNSIGNED #(.width(32)) u_sub_997 (
        .y(_T_10),
        .a(io_rs1),
        .b(io_rs2)
    );
    wire [31:0] diff;
    TAIL #(.width(33), .n(1)) tail_998 (
        .y(diff),
        .in(_T_10)
    );
    wire neq;
    wire [31:0] _WTEMP_78;
    PAD_UNSIGNED #(.width(1), .n(32)) u_pad_999 (
        .y(_WTEMP_78),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(32)) u_neq_1000 (
        .y(neq),
        .a(diff),
        .b(_WTEMP_78)
    );
    wire eq;
    EQ_UNSIGNED #(.width(1)) u_eq_1001 (
        .y(eq),
        .a(neq),
        .b(1'h0)
    );
    wire _T_13;
    BITS #(.width(32), .high(31), .low(31)) bits_1002 (
        .y(_T_13),
        .in(io_rs1)
    );
    wire _T_14;
    BITS #(.width(32), .high(31), .low(31)) bits_1003 (
        .y(_T_14),
        .in(io_rs2)
    );
    wire isSameSign;
    EQ_UNSIGNED #(.width(1)) u_eq_1004 (
        .y(isSameSign),
        .a(_T_13),
        .b(_T_14)
    );
    wire _T_15;
    BITS #(.width(32), .high(31), .low(31)) bits_1005 (
        .y(_T_15),
        .in(diff)
    );
    wire _T_16;
    BITS #(.width(32), .high(31), .low(31)) bits_1006 (
        .y(_T_16),
        .in(io_rs1)
    );
    wire lt;
    MUX_UNSIGNED #(.width(1)) u_mux_1007 (
        .y(lt),
        .sel(isSameSign),
        .a(_T_15),
        .b(_T_16)
    );
    wire _T_17;
    BITS #(.width(32), .high(31), .low(31)) bits_1008 (
        .y(_T_17),
        .in(diff)
    );
    wire _T_18;
    BITS #(.width(32), .high(31), .low(31)) bits_1009 (
        .y(_T_18),
        .in(io_rs2)
    );
    wire ltu;
    MUX_UNSIGNED #(.width(1)) u_mux_1010 (
        .y(ltu),
        .sel(isSameSign),
        .a(_T_17),
        .b(_T_18)
    );
    wire ge;
    EQ_UNSIGNED #(.width(1)) u_eq_1011 (
        .y(ge),
        .a(lt),
        .b(1'h0)
    );
    wire geu;
    EQ_UNSIGNED #(.width(1)) u_eq_1012 (
        .y(geu),
        .a(ltu),
        .b(1'h0)
    );
    wire _T_21;
    EQ_UNSIGNED #(.width(3)) u_eq_1013 (
        .y(_T_21),
        .a(io_br_type),
        .b(3'h3)
    );
    wire _T_22;
    BITWISEAND #(.width(1)) bitwiseand_1014 (
        .y(_T_22),
        .a(_T_21),
        .b(eq)
    );
    wire _T_23;
    EQ_UNSIGNED #(.width(3)) u_eq_1015 (
        .y(_T_23),
        .a(io_br_type),
        .b(3'h6)
    );
    wire _T_24;
    BITWISEAND #(.width(1)) bitwiseand_1016 (
        .y(_T_24),
        .a(_T_23),
        .b(neq)
    );
    wire _T_25;
    BITWISEOR #(.width(1)) bitwiseor_1017 (
        .y(_T_25),
        .a(_T_22),
        .b(_T_24)
    );
    wire _T_26;
    EQ_UNSIGNED #(.width(3)) u_eq_1018 (
        .y(_T_26),
        .a(io_br_type),
        .b(3'h2)
    );
    wire _T_27;
    BITWISEAND #(.width(1)) bitwiseand_1019 (
        .y(_T_27),
        .a(_T_26),
        .b(lt)
    );
    wire _T_28;
    BITWISEOR #(.width(1)) bitwiseor_1020 (
        .y(_T_28),
        .a(_T_25),
        .b(_T_27)
    );
    wire _T_29;
    EQ_UNSIGNED #(.width(3)) u_eq_1021 (
        .y(_T_29),
        .a(io_br_type),
        .b(3'h5)
    );
    wire _T_30;
    BITWISEAND #(.width(1)) bitwiseand_1022 (
        .y(_T_30),
        .a(_T_29),
        .b(ge)
    );
    wire _T_31;
    BITWISEOR #(.width(1)) bitwiseor_1023 (
        .y(_T_31),
        .a(_T_28),
        .b(_T_30)
    );
    wire _T_32;
    EQ_UNSIGNED #(.width(3)) u_eq_1024 (
        .y(_T_32),
        .a(io_br_type),
        .b(3'h1)
    );
    wire _T_33;
    BITWISEAND #(.width(1)) bitwiseand_1025 (
        .y(_T_33),
        .a(_T_32),
        .b(ltu)
    );
    wire _T_34;
    BITWISEOR #(.width(1)) bitwiseor_1026 (
        .y(_T_34),
        .a(_T_31),
        .b(_T_33)
    );
    wire _T_35;
    EQ_UNSIGNED #(.width(3)) u_eq_1027 (
        .y(_T_35),
        .a(io_br_type),
        .b(3'h4)
    );
    wire _T_36;
    BITWISEAND #(.width(1)) bitwiseand_1028 (
        .y(_T_36),
        .a(_T_35),
        .b(geu)
    );
    wire _T_37;
    BITWISEOR #(.width(1)) bitwiseor_1029 (
        .y(_T_37),
        .a(_T_34),
        .b(_T_36)
    );
    assign io_taken = _T_37;
endmodule //BrCondArea
module Control(
    input clock,
    input reset,
    input [31:0] io_inst,
    output [1:0] io_pc_sel,
    output io_inst_kill,
    output io_A_sel,
    output io_B_sel,
    output [2:0] io_imm_sel,
    output [3:0] io_alu_op,
    output [2:0] io_br_type,
    output [1:0] io_st_type,
    output [2:0] io_ld_type,
    output [1:0] io_wb_sel,
    output io_wb_en,
    output [2:0] io_csr_cmd,
    output io_illegal
);
    wire [31:0] _T_32;
    wire [31:0] _WTEMP_103;
    PAD_UNSIGNED #(.width(7), .n(32)) u_pad_1204 (
        .y(_WTEMP_103),
        .in(7'h7F)
    );
    BITWISEAND #(.width(32)) bitwiseand_1205 (
        .y(_T_32),
        .a(io_inst),
        .b(_WTEMP_103)
    );
    wire _T_33;
    wire [31:0] _WTEMP_104;
    PAD_UNSIGNED #(.width(6), .n(32)) u_pad_1206 (
        .y(_WTEMP_104),
        .in(6'h37)
    );
    EQ_UNSIGNED #(.width(32)) u_eq_1207 (
        .y(_T_33),
        .a(_WTEMP_104),
        .b(_T_32)
    );
    wire [31:0] _T_36;
    wire [31:0] _WTEMP_105;
    PAD_UNSIGNED #(.width(7), .n(32)) u_pad_1208 (
        .y(_WTEMP_105),
        .in(7'h7F)
    );
    BITWISEAND #(.width(32)) bitwiseand_1209 (
        .y(_T_36),
        .a(io_inst),
        .b(_WTEMP_105)
    );
    wire _T_37;
    wire [31:0] _WTEMP_106;
    PAD_UNSIGNED #(.width(5), .n(32)) u_pad_1210 (
        .y(_WTEMP_106),
        .in(5'h17)
    );
    EQ_UNSIGNED #(.width(32)) u_eq_1211 (
        .y(_T_37),
        .a(_WTEMP_106),
        .b(_T_36)
    );
    wire [31:0] _T_40;
    wire [31:0] _WTEMP_107;
    PAD_UNSIGNED #(.width(7), .n(32)) u_pad_1212 (
        .y(_WTEMP_107),
        .in(7'h7F)
    );
    BITWISEAND #(.width(32)) bitwiseand_1213 (
        .y(_T_40),
        .a(io_inst),
        .b(_WTEMP_107)
    );
    wire _T_41;
    wire [31:0] _WTEMP_108;
    PAD_UNSIGNED #(.width(7), .n(32)) u_pad_1214 (
        .y(_WTEMP_108),
        .in(7'h6F)
    );
    EQ_UNSIGNED #(.width(32)) u_eq_1215 (
        .y(_T_41),
        .a(_WTEMP_108),
        .b(_T_40)
    );
    wire [31:0] _T_44;
    wire [31:0] _WTEMP_109;
    PAD_UNSIGNED #(.width(15), .n(32)) u_pad_1216 (
        .y(_WTEMP_109),
        .in(15'h707F)
    );
    BITWISEAND #(.width(32)) bitwiseand_1217 (
        .y(_T_44),
        .a(io_inst),
        .b(_WTEMP_109)
    );
    wire _T_45;
    wire [31:0] _WTEMP_110;
    PAD_UNSIGNED #(.width(7), .n(32)) u_pad_1218 (
        .y(_WTEMP_110),
        .in(7'h67)
    );
    EQ_UNSIGNED #(.width(32)) u_eq_1219 (
        .y(_T_45),
        .a(_WTEMP_110),
        .b(_T_44)
    );
    wire [31:0] _T_48;
    wire [31:0] _WTEMP_111;
    PAD_UNSIGNED #(.width(15), .n(32)) u_pad_1220 (
        .y(_WTEMP_111),
        .in(15'h707F)
    );
    BITWISEAND #(.width(32)) bitwiseand_1221 (
        .y(_T_48),
        .a(io_inst),
        .b(_WTEMP_111)
    );
    wire _T_49;
    wire [31:0] _WTEMP_112;
    PAD_UNSIGNED #(.width(7), .n(32)) u_pad_1222 (
        .y(_WTEMP_112),
        .in(7'h63)
    );
    EQ_UNSIGNED #(.width(32)) u_eq_1223 (
        .y(_T_49),
        .a(_WTEMP_112),
        .b(_T_48)
    );
    wire [31:0] _T_52;
    wire [31:0] _WTEMP_113;
    PAD_UNSIGNED #(.width(15), .n(32)) u_pad_1224 (
        .y(_WTEMP_113),
        .in(15'h707F)
    );
    BITWISEAND #(.width(32)) bitwiseand_1225 (
        .y(_T_52),
        .a(io_inst),
        .b(_WTEMP_113)
    );
    wire _T_53;
    wire [31:0] _WTEMP_114;
    PAD_UNSIGNED #(.width(13), .n(32)) u_pad_1226 (
        .y(_WTEMP_114),
        .in(13'h1063)
    );
    EQ_UNSIGNED #(.width(32)) u_eq_1227 (
        .y(_T_53),
        .a(_WTEMP_114),
        .b(_T_52)
    );
    wire [31:0] _T_56;
    wire [31:0] _WTEMP_115;
    PAD_UNSIGNED #(.width(15), .n(32)) u_pad_1228 (
        .y(_WTEMP_115),
        .in(15'h707F)
    );
    BITWISEAND #(.width(32)) bitwiseand_1229 (
        .y(_T_56),
        .a(io_inst),
        .b(_WTEMP_115)
    );
    wire _T_57;
    wire [31:0] _WTEMP_116;
    PAD_UNSIGNED #(.width(15), .n(32)) u_pad_1230 (
        .y(_WTEMP_116),
        .in(15'h4063)
    );
    EQ_UNSIGNED #(.width(32)) u_eq_1231 (
        .y(_T_57),
        .a(_WTEMP_116),
        .b(_T_56)
    );
    wire [31:0] _T_60;
    wire [31:0] _WTEMP_117;
    PAD_UNSIGNED #(.width(15), .n(32)) u_pad_1232 (
        .y(_WTEMP_117),
        .in(15'h707F)
    );
    BITWISEAND #(.width(32)) bitwiseand_1233 (
        .y(_T_60),
        .a(io_inst),
        .b(_WTEMP_117)
    );
    wire _T_61;
    wire [31:0] _WTEMP_118;
    PAD_UNSIGNED #(.width(15), .n(32)) u_pad_1234 (
        .y(_WTEMP_118),
        .in(15'h5063)
    );
    EQ_UNSIGNED #(.width(32)) u_eq_1235 (
        .y(_T_61),
        .a(_WTEMP_118),
        .b(_T_60)
    );
    wire [31:0] _T_64;
    wire [31:0] _WTEMP_119;
    PAD_UNSIGNED #(.width(15), .n(32)) u_pad_1236 (
        .y(_WTEMP_119),
        .in(15'h707F)
    );
    BITWISEAND #(.width(32)) bitwiseand_1237 (
        .y(_T_64),
        .a(io_inst),
        .b(_WTEMP_119)
    );
    wire _T_65;
    wire [31:0] _WTEMP_120;
    PAD_UNSIGNED #(.width(15), .n(32)) u_pad_1238 (
        .y(_WTEMP_120),
        .in(15'h6063)
    );
    EQ_UNSIGNED #(.width(32)) u_eq_1239 (
        .y(_T_65),
        .a(_WTEMP_120),
        .b(_T_64)
    );
    wire [31:0] _T_68;
    wire [31:0] _WTEMP_121;
    PAD_UNSIGNED #(.width(15), .n(32)) u_pad_1240 (
        .y(_WTEMP_121),
        .in(15'h707F)
    );
    BITWISEAND #(.width(32)) bitwiseand_1241 (
        .y(_T_68),
        .a(io_inst),
        .b(_WTEMP_121)
    );
    wire _T_69;
    wire [31:0] _WTEMP_122;
    PAD_UNSIGNED #(.width(15), .n(32)) u_pad_1242 (
        .y(_WTEMP_122),
        .in(15'h7063)
    );
    EQ_UNSIGNED #(.width(32)) u_eq_1243 (
        .y(_T_69),
        .a(_WTEMP_122),
        .b(_T_68)
    );
    wire [31:0] _T_72;
    wire [31:0] _WTEMP_123;
    PAD_UNSIGNED #(.width(15), .n(32)) u_pad_1244 (
        .y(_WTEMP_123),
        .in(15'h707F)
    );
    BITWISEAND #(.width(32)) bitwiseand_1245 (
        .y(_T_72),
        .a(io_inst),
        .b(_WTEMP_123)
    );
    wire _T_73;
    wire [31:0] _WTEMP_124;
    PAD_UNSIGNED #(.width(2), .n(32)) u_pad_1246 (
        .y(_WTEMP_124),
        .in(2'h3)
    );
    EQ_UNSIGNED #(.width(32)) u_eq_1247 (
        .y(_T_73),
        .a(_WTEMP_124),
        .b(_T_72)
    );
    wire [31:0] _T_76;
    wire [31:0] _WTEMP_125;
    PAD_UNSIGNED #(.width(15), .n(32)) u_pad_1248 (
        .y(_WTEMP_125),
        .in(15'h707F)
    );
    BITWISEAND #(.width(32)) bitwiseand_1249 (
        .y(_T_76),
        .a(io_inst),
        .b(_WTEMP_125)
    );
    wire _T_77;
    wire [31:0] _WTEMP_126;
    PAD_UNSIGNED #(.width(13), .n(32)) u_pad_1250 (
        .y(_WTEMP_126),
        .in(13'h1003)
    );
    EQ_UNSIGNED #(.width(32)) u_eq_1251 (
        .y(_T_77),
        .a(_WTEMP_126),
        .b(_T_76)
    );
    wire [31:0] _T_80;
    wire [31:0] _WTEMP_127;
    PAD_UNSIGNED #(.width(15), .n(32)) u_pad_1252 (
        .y(_WTEMP_127),
        .in(15'h707F)
    );
    BITWISEAND #(.width(32)) bitwiseand_1253 (
        .y(_T_80),
        .a(io_inst),
        .b(_WTEMP_127)
    );
    wire _T_81;
    wire [31:0] _WTEMP_128;
    PAD_UNSIGNED #(.width(14), .n(32)) u_pad_1254 (
        .y(_WTEMP_128),
        .in(14'h2003)
    );
    EQ_UNSIGNED #(.width(32)) u_eq_1255 (
        .y(_T_81),
        .a(_WTEMP_128),
        .b(_T_80)
    );
    wire [31:0] _T_84;
    wire [31:0] _WTEMP_129;
    PAD_UNSIGNED #(.width(15), .n(32)) u_pad_1256 (
        .y(_WTEMP_129),
        .in(15'h707F)
    );
    BITWISEAND #(.width(32)) bitwiseand_1257 (
        .y(_T_84),
        .a(io_inst),
        .b(_WTEMP_129)
    );
    wire _T_85;
    wire [31:0] _WTEMP_130;
    PAD_UNSIGNED #(.width(15), .n(32)) u_pad_1258 (
        .y(_WTEMP_130),
        .in(15'h4003)
    );
    EQ_UNSIGNED #(.width(32)) u_eq_1259 (
        .y(_T_85),
        .a(_WTEMP_130),
        .b(_T_84)
    );
    wire [31:0] _T_88;
    wire [31:0] _WTEMP_131;
    PAD_UNSIGNED #(.width(15), .n(32)) u_pad_1260 (
        .y(_WTEMP_131),
        .in(15'h707F)
    );
    BITWISEAND #(.width(32)) bitwiseand_1261 (
        .y(_T_88),
        .a(io_inst),
        .b(_WTEMP_131)
    );
    wire _T_89;
    wire [31:0] _WTEMP_132;
    PAD_UNSIGNED #(.width(15), .n(32)) u_pad_1262 (
        .y(_WTEMP_132),
        .in(15'h5003)
    );
    EQ_UNSIGNED #(.width(32)) u_eq_1263 (
        .y(_T_89),
        .a(_WTEMP_132),
        .b(_T_88)
    );
    wire [31:0] _T_92;
    wire [31:0] _WTEMP_133;
    PAD_UNSIGNED #(.width(15), .n(32)) u_pad_1264 (
        .y(_WTEMP_133),
        .in(15'h707F)
    );
    BITWISEAND #(.width(32)) bitwiseand_1265 (
        .y(_T_92),
        .a(io_inst),
        .b(_WTEMP_133)
    );
    wire _T_93;
    wire [31:0] _WTEMP_134;
    PAD_UNSIGNED #(.width(6), .n(32)) u_pad_1266 (
        .y(_WTEMP_134),
        .in(6'h23)
    );
    EQ_UNSIGNED #(.width(32)) u_eq_1267 (
        .y(_T_93),
        .a(_WTEMP_134),
        .b(_T_92)
    );
    wire [31:0] _T_96;
    wire [31:0] _WTEMP_135;
    PAD_UNSIGNED #(.width(15), .n(32)) u_pad_1268 (
        .y(_WTEMP_135),
        .in(15'h707F)
    );
    BITWISEAND #(.width(32)) bitwiseand_1269 (
        .y(_T_96),
        .a(io_inst),
        .b(_WTEMP_135)
    );
    wire _T_97;
    wire [31:0] _WTEMP_136;
    PAD_UNSIGNED #(.width(13), .n(32)) u_pad_1270 (
        .y(_WTEMP_136),
        .in(13'h1023)
    );
    EQ_UNSIGNED #(.width(32)) u_eq_1271 (
        .y(_T_97),
        .a(_WTEMP_136),
        .b(_T_96)
    );
    wire [31:0] _T_100;
    wire [31:0] _WTEMP_137;
    PAD_UNSIGNED #(.width(15), .n(32)) u_pad_1272 (
        .y(_WTEMP_137),
        .in(15'h707F)
    );
    BITWISEAND #(.width(32)) bitwiseand_1273 (
        .y(_T_100),
        .a(io_inst),
        .b(_WTEMP_137)
    );
    wire _T_101;
    wire [31:0] _WTEMP_138;
    PAD_UNSIGNED #(.width(14), .n(32)) u_pad_1274 (
        .y(_WTEMP_138),
        .in(14'h2023)
    );
    EQ_UNSIGNED #(.width(32)) u_eq_1275 (
        .y(_T_101),
        .a(_WTEMP_138),
        .b(_T_100)
    );
    wire [31:0] _T_104;
    wire [31:0] _WTEMP_139;
    PAD_UNSIGNED #(.width(15), .n(32)) u_pad_1276 (
        .y(_WTEMP_139),
        .in(15'h707F)
    );
    BITWISEAND #(.width(32)) bitwiseand_1277 (
        .y(_T_104),
        .a(io_inst),
        .b(_WTEMP_139)
    );
    wire _T_105;
    wire [31:0] _WTEMP_140;
    PAD_UNSIGNED #(.width(5), .n(32)) u_pad_1278 (
        .y(_WTEMP_140),
        .in(5'h13)
    );
    EQ_UNSIGNED #(.width(32)) u_eq_1279 (
        .y(_T_105),
        .a(_WTEMP_140),
        .b(_T_104)
    );
    wire [31:0] _T_108;
    wire [31:0] _WTEMP_141;
    PAD_UNSIGNED #(.width(15), .n(32)) u_pad_1280 (
        .y(_WTEMP_141),
        .in(15'h707F)
    );
    BITWISEAND #(.width(32)) bitwiseand_1281 (
        .y(_T_108),
        .a(io_inst),
        .b(_WTEMP_141)
    );
    wire _T_109;
    wire [31:0] _WTEMP_142;
    PAD_UNSIGNED #(.width(14), .n(32)) u_pad_1282 (
        .y(_WTEMP_142),
        .in(14'h2013)
    );
    EQ_UNSIGNED #(.width(32)) u_eq_1283 (
        .y(_T_109),
        .a(_WTEMP_142),
        .b(_T_108)
    );
    wire [31:0] _T_112;
    wire [31:0] _WTEMP_143;
    PAD_UNSIGNED #(.width(15), .n(32)) u_pad_1284 (
        .y(_WTEMP_143),
        .in(15'h707F)
    );
    BITWISEAND #(.width(32)) bitwiseand_1285 (
        .y(_T_112),
        .a(io_inst),
        .b(_WTEMP_143)
    );
    wire _T_113;
    wire [31:0] _WTEMP_144;
    PAD_UNSIGNED #(.width(14), .n(32)) u_pad_1286 (
        .y(_WTEMP_144),
        .in(14'h3013)
    );
    EQ_UNSIGNED #(.width(32)) u_eq_1287 (
        .y(_T_113),
        .a(_WTEMP_144),
        .b(_T_112)
    );
    wire [31:0] _T_116;
    wire [31:0] _WTEMP_145;
    PAD_UNSIGNED #(.width(15), .n(32)) u_pad_1288 (
        .y(_WTEMP_145),
        .in(15'h707F)
    );
    BITWISEAND #(.width(32)) bitwiseand_1289 (
        .y(_T_116),
        .a(io_inst),
        .b(_WTEMP_145)
    );
    wire _T_117;
    wire [31:0] _WTEMP_146;
    PAD_UNSIGNED #(.width(15), .n(32)) u_pad_1290 (
        .y(_WTEMP_146),
        .in(15'h4013)
    );
    EQ_UNSIGNED #(.width(32)) u_eq_1291 (
        .y(_T_117),
        .a(_WTEMP_146),
        .b(_T_116)
    );
    wire [31:0] _T_120;
    wire [31:0] _WTEMP_147;
    PAD_UNSIGNED #(.width(15), .n(32)) u_pad_1292 (
        .y(_WTEMP_147),
        .in(15'h707F)
    );
    BITWISEAND #(.width(32)) bitwiseand_1293 (
        .y(_T_120),
        .a(io_inst),
        .b(_WTEMP_147)
    );
    wire _T_121;
    wire [31:0] _WTEMP_148;
    PAD_UNSIGNED #(.width(15), .n(32)) u_pad_1294 (
        .y(_WTEMP_148),
        .in(15'h6013)
    );
    EQ_UNSIGNED #(.width(32)) u_eq_1295 (
        .y(_T_121),
        .a(_WTEMP_148),
        .b(_T_120)
    );
    wire [31:0] _T_124;
    wire [31:0] _WTEMP_149;
    PAD_UNSIGNED #(.width(15), .n(32)) u_pad_1296 (
        .y(_WTEMP_149),
        .in(15'h707F)
    );
    BITWISEAND #(.width(32)) bitwiseand_1297 (
        .y(_T_124),
        .a(io_inst),
        .b(_WTEMP_149)
    );
    wire _T_125;
    wire [31:0] _WTEMP_150;
    PAD_UNSIGNED #(.width(15), .n(32)) u_pad_1298 (
        .y(_WTEMP_150),
        .in(15'h7013)
    );
    EQ_UNSIGNED #(.width(32)) u_eq_1299 (
        .y(_T_125),
        .a(_WTEMP_150),
        .b(_T_124)
    );
    wire [31:0] _T_128;
    BITWISEAND #(.width(32)) bitwiseand_1300 (
        .y(_T_128),
        .a(io_inst),
        .b(32'hFE00707F)
    );
    wire _T_129;
    wire [31:0] _WTEMP_151;
    PAD_UNSIGNED #(.width(13), .n(32)) u_pad_1301 (
        .y(_WTEMP_151),
        .in(13'h1013)
    );
    EQ_UNSIGNED #(.width(32)) u_eq_1302 (
        .y(_T_129),
        .a(_WTEMP_151),
        .b(_T_128)
    );
    wire [31:0] _T_132;
    BITWISEAND #(.width(32)) bitwiseand_1303 (
        .y(_T_132),
        .a(io_inst),
        .b(32'hFE00707F)
    );
    wire _T_133;
    wire [31:0] _WTEMP_152;
    PAD_UNSIGNED #(.width(15), .n(32)) u_pad_1304 (
        .y(_WTEMP_152),
        .in(15'h5013)
    );
    EQ_UNSIGNED #(.width(32)) u_eq_1305 (
        .y(_T_133),
        .a(_WTEMP_152),
        .b(_T_132)
    );
    wire [31:0] _T_136;
    BITWISEAND #(.width(32)) bitwiseand_1306 (
        .y(_T_136),
        .a(io_inst),
        .b(32'hFE00707F)
    );
    wire _T_137;
    wire [31:0] _WTEMP_153;
    PAD_UNSIGNED #(.width(31), .n(32)) u_pad_1307 (
        .y(_WTEMP_153),
        .in(31'h40005013)
    );
    EQ_UNSIGNED #(.width(32)) u_eq_1308 (
        .y(_T_137),
        .a(_WTEMP_153),
        .b(_T_136)
    );
    wire [31:0] _T_140;
    BITWISEAND #(.width(32)) bitwiseand_1309 (
        .y(_T_140),
        .a(io_inst),
        .b(32'hFE00707F)
    );
    wire _T_141;
    wire [31:0] _WTEMP_154;
    PAD_UNSIGNED #(.width(6), .n(32)) u_pad_1310 (
        .y(_WTEMP_154),
        .in(6'h33)
    );
    EQ_UNSIGNED #(.width(32)) u_eq_1311 (
        .y(_T_141),
        .a(_WTEMP_154),
        .b(_T_140)
    );
    wire [31:0] _T_144;
    BITWISEAND #(.width(32)) bitwiseand_1312 (
        .y(_T_144),
        .a(io_inst),
        .b(32'hFE00707F)
    );
    wire _T_145;
    wire [31:0] _WTEMP_155;
    PAD_UNSIGNED #(.width(31), .n(32)) u_pad_1313 (
        .y(_WTEMP_155),
        .in(31'h40000033)
    );
    EQ_UNSIGNED #(.width(32)) u_eq_1314 (
        .y(_T_145),
        .a(_WTEMP_155),
        .b(_T_144)
    );
    wire [31:0] _T_148;
    BITWISEAND #(.width(32)) bitwiseand_1315 (
        .y(_T_148),
        .a(io_inst),
        .b(32'hFE00707F)
    );
    wire _T_149;
    wire [31:0] _WTEMP_156;
    PAD_UNSIGNED #(.width(13), .n(32)) u_pad_1316 (
        .y(_WTEMP_156),
        .in(13'h1033)
    );
    EQ_UNSIGNED #(.width(32)) u_eq_1317 (
        .y(_T_149),
        .a(_WTEMP_156),
        .b(_T_148)
    );
    wire [31:0] _T_152;
    BITWISEAND #(.width(32)) bitwiseand_1318 (
        .y(_T_152),
        .a(io_inst),
        .b(32'hFE00707F)
    );
    wire _T_153;
    wire [31:0] _WTEMP_157;
    PAD_UNSIGNED #(.width(14), .n(32)) u_pad_1319 (
        .y(_WTEMP_157),
        .in(14'h2033)
    );
    EQ_UNSIGNED #(.width(32)) u_eq_1320 (
        .y(_T_153),
        .a(_WTEMP_157),
        .b(_T_152)
    );
    wire [31:0] _T_156;
    BITWISEAND #(.width(32)) bitwiseand_1321 (
        .y(_T_156),
        .a(io_inst),
        .b(32'hFE00707F)
    );
    wire _T_157;
    wire [31:0] _WTEMP_158;
    PAD_UNSIGNED #(.width(14), .n(32)) u_pad_1322 (
        .y(_WTEMP_158),
        .in(14'h3033)
    );
    EQ_UNSIGNED #(.width(32)) u_eq_1323 (
        .y(_T_157),
        .a(_WTEMP_158),
        .b(_T_156)
    );
    wire [31:0] _T_160;
    BITWISEAND #(.width(32)) bitwiseand_1324 (
        .y(_T_160),
        .a(io_inst),
        .b(32'hFE00707F)
    );
    wire _T_161;
    wire [31:0] _WTEMP_159;
    PAD_UNSIGNED #(.width(15), .n(32)) u_pad_1325 (
        .y(_WTEMP_159),
        .in(15'h4033)
    );
    EQ_UNSIGNED #(.width(32)) u_eq_1326 (
        .y(_T_161),
        .a(_WTEMP_159),
        .b(_T_160)
    );
    wire [31:0] _T_164;
    BITWISEAND #(.width(32)) bitwiseand_1327 (
        .y(_T_164),
        .a(io_inst),
        .b(32'hFE00707F)
    );
    wire _T_165;
    wire [31:0] _WTEMP_160;
    PAD_UNSIGNED #(.width(15), .n(32)) u_pad_1328 (
        .y(_WTEMP_160),
        .in(15'h5033)
    );
    EQ_UNSIGNED #(.width(32)) u_eq_1329 (
        .y(_T_165),
        .a(_WTEMP_160),
        .b(_T_164)
    );
    wire [31:0] _T_168;
    BITWISEAND #(.width(32)) bitwiseand_1330 (
        .y(_T_168),
        .a(io_inst),
        .b(32'hFE00707F)
    );
    wire _T_169;
    wire [31:0] _WTEMP_161;
    PAD_UNSIGNED #(.width(31), .n(32)) u_pad_1331 (
        .y(_WTEMP_161),
        .in(31'h40005033)
    );
    EQ_UNSIGNED #(.width(32)) u_eq_1332 (
        .y(_T_169),
        .a(_WTEMP_161),
        .b(_T_168)
    );
    wire [31:0] _T_172;
    BITWISEAND #(.width(32)) bitwiseand_1333 (
        .y(_T_172),
        .a(io_inst),
        .b(32'hFE00707F)
    );
    wire _T_173;
    wire [31:0] _WTEMP_162;
    PAD_UNSIGNED #(.width(15), .n(32)) u_pad_1334 (
        .y(_WTEMP_162),
        .in(15'h6033)
    );
    EQ_UNSIGNED #(.width(32)) u_eq_1335 (
        .y(_T_173),
        .a(_WTEMP_162),
        .b(_T_172)
    );
    wire [31:0] _T_176;
    BITWISEAND #(.width(32)) bitwiseand_1336 (
        .y(_T_176),
        .a(io_inst),
        .b(32'hFE00707F)
    );
    wire _T_177;
    wire [31:0] _WTEMP_163;
    PAD_UNSIGNED #(.width(15), .n(32)) u_pad_1337 (
        .y(_WTEMP_163),
        .in(15'h7033)
    );
    EQ_UNSIGNED #(.width(32)) u_eq_1338 (
        .y(_T_177),
        .a(_WTEMP_163),
        .b(_T_176)
    );
    wire [31:0] _T_180;
    BITWISEAND #(.width(32)) bitwiseand_1339 (
        .y(_T_180),
        .a(io_inst),
        .b(32'hF00FFFFF)
    );
    wire _T_181;
    wire [31:0] _WTEMP_164;
    PAD_UNSIGNED #(.width(4), .n(32)) u_pad_1340 (
        .y(_WTEMP_164),
        .in(4'hF)
    );
    EQ_UNSIGNED #(.width(32)) u_eq_1341 (
        .y(_T_181),
        .a(_WTEMP_164),
        .b(_T_180)
    );
    wire [31:0] _T_184;
    BITWISEAND #(.width(32)) bitwiseand_1342 (
        .y(_T_184),
        .a(io_inst),
        .b(32'hFFFFFFFF)
    );
    wire _T_185;
    wire [31:0] _WTEMP_165;
    PAD_UNSIGNED #(.width(13), .n(32)) u_pad_1343 (
        .y(_WTEMP_165),
        .in(13'h100F)
    );
    EQ_UNSIGNED #(.width(32)) u_eq_1344 (
        .y(_T_185),
        .a(_WTEMP_165),
        .b(_T_184)
    );
    wire [31:0] _T_188;
    wire [31:0] _WTEMP_166;
    PAD_UNSIGNED #(.width(15), .n(32)) u_pad_1345 (
        .y(_WTEMP_166),
        .in(15'h707F)
    );
    BITWISEAND #(.width(32)) bitwiseand_1346 (
        .y(_T_188),
        .a(io_inst),
        .b(_WTEMP_166)
    );
    wire _T_189;
    wire [31:0] _WTEMP_167;
    PAD_UNSIGNED #(.width(13), .n(32)) u_pad_1347 (
        .y(_WTEMP_167),
        .in(13'h1073)
    );
    EQ_UNSIGNED #(.width(32)) u_eq_1348 (
        .y(_T_189),
        .a(_WTEMP_167),
        .b(_T_188)
    );
    wire [31:0] _T_192;
    wire [31:0] _WTEMP_168;
    PAD_UNSIGNED #(.width(15), .n(32)) u_pad_1349 (
        .y(_WTEMP_168),
        .in(15'h707F)
    );
    BITWISEAND #(.width(32)) bitwiseand_1350 (
        .y(_T_192),
        .a(io_inst),
        .b(_WTEMP_168)
    );
    wire _T_193;
    wire [31:0] _WTEMP_169;
    PAD_UNSIGNED #(.width(14), .n(32)) u_pad_1351 (
        .y(_WTEMP_169),
        .in(14'h2073)
    );
    EQ_UNSIGNED #(.width(32)) u_eq_1352 (
        .y(_T_193),
        .a(_WTEMP_169),
        .b(_T_192)
    );
    wire [31:0] _T_196;
    wire [31:0] _WTEMP_170;
    PAD_UNSIGNED #(.width(15), .n(32)) u_pad_1353 (
        .y(_WTEMP_170),
        .in(15'h707F)
    );
    BITWISEAND #(.width(32)) bitwiseand_1354 (
        .y(_T_196),
        .a(io_inst),
        .b(_WTEMP_170)
    );
    wire _T_197;
    wire [31:0] _WTEMP_171;
    PAD_UNSIGNED #(.width(14), .n(32)) u_pad_1355 (
        .y(_WTEMP_171),
        .in(14'h3073)
    );
    EQ_UNSIGNED #(.width(32)) u_eq_1356 (
        .y(_T_197),
        .a(_WTEMP_171),
        .b(_T_196)
    );
    wire [31:0] _T_200;
    wire [31:0] _WTEMP_172;
    PAD_UNSIGNED #(.width(15), .n(32)) u_pad_1357 (
        .y(_WTEMP_172),
        .in(15'h707F)
    );
    BITWISEAND #(.width(32)) bitwiseand_1358 (
        .y(_T_200),
        .a(io_inst),
        .b(_WTEMP_172)
    );
    wire _T_201;
    wire [31:0] _WTEMP_173;
    PAD_UNSIGNED #(.width(15), .n(32)) u_pad_1359 (
        .y(_WTEMP_173),
        .in(15'h5073)
    );
    EQ_UNSIGNED #(.width(32)) u_eq_1360 (
        .y(_T_201),
        .a(_WTEMP_173),
        .b(_T_200)
    );
    wire [31:0] _T_204;
    wire [31:0] _WTEMP_174;
    PAD_UNSIGNED #(.width(15), .n(32)) u_pad_1361 (
        .y(_WTEMP_174),
        .in(15'h707F)
    );
    BITWISEAND #(.width(32)) bitwiseand_1362 (
        .y(_T_204),
        .a(io_inst),
        .b(_WTEMP_174)
    );
    wire _T_205;
    wire [31:0] _WTEMP_175;
    PAD_UNSIGNED #(.width(15), .n(32)) u_pad_1363 (
        .y(_WTEMP_175),
        .in(15'h6073)
    );
    EQ_UNSIGNED #(.width(32)) u_eq_1364 (
        .y(_T_205),
        .a(_WTEMP_175),
        .b(_T_204)
    );
    wire [31:0] _T_208;
    wire [31:0] _WTEMP_176;
    PAD_UNSIGNED #(.width(15), .n(32)) u_pad_1365 (
        .y(_WTEMP_176),
        .in(15'h707F)
    );
    BITWISEAND #(.width(32)) bitwiseand_1366 (
        .y(_T_208),
        .a(io_inst),
        .b(_WTEMP_176)
    );
    wire _T_209;
    wire [31:0] _WTEMP_177;
    PAD_UNSIGNED #(.width(15), .n(32)) u_pad_1367 (
        .y(_WTEMP_177),
        .in(15'h7073)
    );
    EQ_UNSIGNED #(.width(32)) u_eq_1368 (
        .y(_T_209),
        .a(_WTEMP_177),
        .b(_T_208)
    );
    wire [31:0] _T_212;
    BITWISEAND #(.width(32)) bitwiseand_1369 (
        .y(_T_212),
        .a(io_inst),
        .b(32'hFFFFFFFF)
    );
    wire _T_213;
    wire [31:0] _WTEMP_178;
    PAD_UNSIGNED #(.width(7), .n(32)) u_pad_1370 (
        .y(_WTEMP_178),
        .in(7'h73)
    );
    EQ_UNSIGNED #(.width(32)) u_eq_1371 (
        .y(_T_213),
        .a(_WTEMP_178),
        .b(_T_212)
    );
    wire [31:0] _T_216;
    BITWISEAND #(.width(32)) bitwiseand_1372 (
        .y(_T_216),
        .a(io_inst),
        .b(32'hFFFFFFFF)
    );
    wire _T_217;
    wire [31:0] _WTEMP_179;
    PAD_UNSIGNED #(.width(21), .n(32)) u_pad_1373 (
        .y(_WTEMP_179),
        .in(21'h100073)
    );
    EQ_UNSIGNED #(.width(32)) u_eq_1374 (
        .y(_T_217),
        .a(_WTEMP_179),
        .b(_T_216)
    );
    wire [31:0] _T_220;
    BITWISEAND #(.width(32)) bitwiseand_1375 (
        .y(_T_220),
        .a(io_inst),
        .b(32'hFFFFFFFF)
    );
    wire _T_221;
    wire [31:0] _WTEMP_180;
    PAD_UNSIGNED #(.width(29), .n(32)) u_pad_1376 (
        .y(_WTEMP_180),
        .in(29'h10000073)
    );
    EQ_UNSIGNED #(.width(32)) u_eq_1377 (
        .y(_T_221),
        .a(_WTEMP_180),
        .b(_T_220)
    );
    wire [31:0] _T_224;
    BITWISEAND #(.width(32)) bitwiseand_1378 (
        .y(_T_224),
        .a(io_inst),
        .b(32'hFFFFFFFF)
    );
    wire _T_225;
    wire [31:0] _WTEMP_181;
    PAD_UNSIGNED #(.width(29), .n(32)) u_pad_1379 (
        .y(_WTEMP_181),
        .in(29'h10200073)
    );
    EQ_UNSIGNED #(.width(32)) u_eq_1380 (
        .y(_T_225),
        .a(_WTEMP_181),
        .b(_T_224)
    );
    wire [1:0] _T_226;
    assign _T_226 = 2'h0;
    wire [1:0] _T_227;
    MUX_UNSIGNED #(.width(2)) u_mux_1381 (
        .y(_T_227),
        .sel(_T_221),
        .a(2'h3),
        .b(_T_226)
    );
    wire [1:0] _T_228;
    MUX_UNSIGNED #(.width(2)) u_mux_1382 (
        .y(_T_228),
        .sel(_T_217),
        .a(2'h0),
        .b(_T_227)
    );
    wire [1:0] _T_229;
    MUX_UNSIGNED #(.width(2)) u_mux_1383 (
        .y(_T_229),
        .sel(_T_213),
        .a(2'h0),
        .b(_T_228)
    );
    wire [1:0] _T_230;
    MUX_UNSIGNED #(.width(2)) u_mux_1384 (
        .y(_T_230),
        .sel(_T_209),
        .a(2'h2),
        .b(_T_229)
    );
    wire [1:0] _T_231;
    MUX_UNSIGNED #(.width(2)) u_mux_1385 (
        .y(_T_231),
        .sel(_T_205),
        .a(2'h2),
        .b(_T_230)
    );
    wire [1:0] _T_232;
    MUX_UNSIGNED #(.width(2)) u_mux_1386 (
        .y(_T_232),
        .sel(_T_201),
        .a(2'h2),
        .b(_T_231)
    );
    wire [1:0] _T_233;
    MUX_UNSIGNED #(.width(2)) u_mux_1387 (
        .y(_T_233),
        .sel(_T_197),
        .a(2'h2),
        .b(_T_232)
    );
    wire [1:0] _T_234;
    MUX_UNSIGNED #(.width(2)) u_mux_1388 (
        .y(_T_234),
        .sel(_T_193),
        .a(2'h2),
        .b(_T_233)
    );
    wire [1:0] _T_235;
    MUX_UNSIGNED #(.width(2)) u_mux_1389 (
        .y(_T_235),
        .sel(_T_189),
        .a(2'h2),
        .b(_T_234)
    );
    wire [1:0] _T_236;
    MUX_UNSIGNED #(.width(2)) u_mux_1390 (
        .y(_T_236),
        .sel(_T_185),
        .a(2'h2),
        .b(_T_235)
    );
    wire [1:0] _T_237;
    MUX_UNSIGNED #(.width(2)) u_mux_1391 (
        .y(_T_237),
        .sel(_T_181),
        .a(2'h0),
        .b(_T_236)
    );
    wire [1:0] _T_238;
    MUX_UNSIGNED #(.width(2)) u_mux_1392 (
        .y(_T_238),
        .sel(_T_177),
        .a(2'h0),
        .b(_T_237)
    );
    wire [1:0] _T_239;
    MUX_UNSIGNED #(.width(2)) u_mux_1393 (
        .y(_T_239),
        .sel(_T_173),
        .a(2'h0),
        .b(_T_238)
    );
    wire [1:0] _T_240;
    MUX_UNSIGNED #(.width(2)) u_mux_1394 (
        .y(_T_240),
        .sel(_T_169),
        .a(2'h0),
        .b(_T_239)
    );
    wire [1:0] _T_241;
    MUX_UNSIGNED #(.width(2)) u_mux_1395 (
        .y(_T_241),
        .sel(_T_165),
        .a(2'h0),
        .b(_T_240)
    );
    wire [1:0] _T_242;
    MUX_UNSIGNED #(.width(2)) u_mux_1396 (
        .y(_T_242),
        .sel(_T_161),
        .a(2'h0),
        .b(_T_241)
    );
    wire [1:0] _T_243;
    MUX_UNSIGNED #(.width(2)) u_mux_1397 (
        .y(_T_243),
        .sel(_T_157),
        .a(2'h0),
        .b(_T_242)
    );
    wire [1:0] _T_244;
    MUX_UNSIGNED #(.width(2)) u_mux_1398 (
        .y(_T_244),
        .sel(_T_153),
        .a(2'h0),
        .b(_T_243)
    );
    wire [1:0] _T_245;
    MUX_UNSIGNED #(.width(2)) u_mux_1399 (
        .y(_T_245),
        .sel(_T_149),
        .a(2'h0),
        .b(_T_244)
    );
    wire [1:0] _T_246;
    MUX_UNSIGNED #(.width(2)) u_mux_1400 (
        .y(_T_246),
        .sel(_T_145),
        .a(2'h0),
        .b(_T_245)
    );
    wire [1:0] _T_247;
    MUX_UNSIGNED #(.width(2)) u_mux_1401 (
        .y(_T_247),
        .sel(_T_141),
        .a(2'h0),
        .b(_T_246)
    );
    wire [1:0] _T_248;
    MUX_UNSIGNED #(.width(2)) u_mux_1402 (
        .y(_T_248),
        .sel(_T_137),
        .a(2'h0),
        .b(_T_247)
    );
    wire [1:0] _T_249;
    MUX_UNSIGNED #(.width(2)) u_mux_1403 (
        .y(_T_249),
        .sel(_T_133),
        .a(2'h0),
        .b(_T_248)
    );
    wire [1:0] _T_250;
    MUX_UNSIGNED #(.width(2)) u_mux_1404 (
        .y(_T_250),
        .sel(_T_129),
        .a(2'h0),
        .b(_T_249)
    );
    wire [1:0] _T_251;
    MUX_UNSIGNED #(.width(2)) u_mux_1405 (
        .y(_T_251),
        .sel(_T_125),
        .a(2'h0),
        .b(_T_250)
    );
    wire [1:0] _T_252;
    MUX_UNSIGNED #(.width(2)) u_mux_1406 (
        .y(_T_252),
        .sel(_T_121),
        .a(2'h0),
        .b(_T_251)
    );
    wire [1:0] _T_253;
    MUX_UNSIGNED #(.width(2)) u_mux_1407 (
        .y(_T_253),
        .sel(_T_117),
        .a(2'h0),
        .b(_T_252)
    );
    wire [1:0] _T_254;
    MUX_UNSIGNED #(.width(2)) u_mux_1408 (
        .y(_T_254),
        .sel(_T_113),
        .a(2'h0),
        .b(_T_253)
    );
    wire [1:0] _T_255;
    MUX_UNSIGNED #(.width(2)) u_mux_1409 (
        .y(_T_255),
        .sel(_T_109),
        .a(2'h0),
        .b(_T_254)
    );
    wire [1:0] _T_256;
    MUX_UNSIGNED #(.width(2)) u_mux_1410 (
        .y(_T_256),
        .sel(_T_105),
        .a(2'h0),
        .b(_T_255)
    );
    wire [1:0] _T_257;
    MUX_UNSIGNED #(.width(2)) u_mux_1411 (
        .y(_T_257),
        .sel(_T_101),
        .a(2'h0),
        .b(_T_256)
    );
    wire [1:0] _T_258;
    MUX_UNSIGNED #(.width(2)) u_mux_1412 (
        .y(_T_258),
        .sel(_T_97),
        .a(2'h0),
        .b(_T_257)
    );
    wire [1:0] _T_259;
    MUX_UNSIGNED #(.width(2)) u_mux_1413 (
        .y(_T_259),
        .sel(_T_93),
        .a(2'h0),
        .b(_T_258)
    );
    wire [1:0] _T_260;
    MUX_UNSIGNED #(.width(2)) u_mux_1414 (
        .y(_T_260),
        .sel(_T_89),
        .a(2'h2),
        .b(_T_259)
    );
    wire [1:0] _T_261;
    MUX_UNSIGNED #(.width(2)) u_mux_1415 (
        .y(_T_261),
        .sel(_T_85),
        .a(2'h2),
        .b(_T_260)
    );
    wire [1:0] _T_262;
    MUX_UNSIGNED #(.width(2)) u_mux_1416 (
        .y(_T_262),
        .sel(_T_81),
        .a(2'h2),
        .b(_T_261)
    );
    wire [1:0] _T_263;
    MUX_UNSIGNED #(.width(2)) u_mux_1417 (
        .y(_T_263),
        .sel(_T_77),
        .a(2'h2),
        .b(_T_262)
    );
    wire [1:0] _T_264;
    MUX_UNSIGNED #(.width(2)) u_mux_1418 (
        .y(_T_264),
        .sel(_T_73),
        .a(2'h2),
        .b(_T_263)
    );
    wire [1:0] _T_265;
    MUX_UNSIGNED #(.width(2)) u_mux_1419 (
        .y(_T_265),
        .sel(_T_69),
        .a(2'h0),
        .b(_T_264)
    );
    wire [1:0] _T_266;
    MUX_UNSIGNED #(.width(2)) u_mux_1420 (
        .y(_T_266),
        .sel(_T_65),
        .a(2'h0),
        .b(_T_265)
    );
    wire [1:0] _T_267;
    MUX_UNSIGNED #(.width(2)) u_mux_1421 (
        .y(_T_267),
        .sel(_T_61),
        .a(2'h0),
        .b(_T_266)
    );
    wire [1:0] _T_268;
    MUX_UNSIGNED #(.width(2)) u_mux_1422 (
        .y(_T_268),
        .sel(_T_57),
        .a(2'h0),
        .b(_T_267)
    );
    wire [1:0] _T_269;
    MUX_UNSIGNED #(.width(2)) u_mux_1423 (
        .y(_T_269),
        .sel(_T_53),
        .a(2'h0),
        .b(_T_268)
    );
    wire [1:0] _T_270;
    MUX_UNSIGNED #(.width(2)) u_mux_1424 (
        .y(_T_270),
        .sel(_T_49),
        .a(2'h0),
        .b(_T_269)
    );
    wire [1:0] _T_271;
    MUX_UNSIGNED #(.width(2)) u_mux_1425 (
        .y(_T_271),
        .sel(_T_45),
        .a(2'h1),
        .b(_T_270)
    );
    wire [1:0] _T_272;
    MUX_UNSIGNED #(.width(2)) u_mux_1426 (
        .y(_T_272),
        .sel(_T_41),
        .a(2'h1),
        .b(_T_271)
    );
    wire [1:0] _T_273;
    MUX_UNSIGNED #(.width(2)) u_mux_1427 (
        .y(_T_273),
        .sel(_T_37),
        .a(2'h0),
        .b(_T_272)
    );
    wire [1:0] ctrlSignals_0;
    MUX_UNSIGNED #(.width(2)) u_mux_1428 (
        .y(ctrlSignals_0),
        .sel(_T_33),
        .a(2'h0),
        .b(_T_273)
    );
    wire _T_274;
    assign _T_274 = 1'h0;
    wire _T_275;
    assign _T_275 = 1'h0;
    wire _T_276;
    assign _T_276 = 1'h0;
    wire _T_277;
    assign _T_277 = 1'h0;
    wire _T_278;
    assign _T_278 = 1'h0;
    wire _T_279;
    assign _T_279 = 1'h0;
    wire _T_280;
    assign _T_280 = 1'h0;
    wire _T_281;
    MUX_UNSIGNED #(.width(1)) u_mux_1429 (
        .y(_T_281),
        .sel(_T_197),
        .a(1'h1),
        .b(_T_280)
    );
    wire _T_282;
    MUX_UNSIGNED #(.width(1)) u_mux_1430 (
        .y(_T_282),
        .sel(_T_193),
        .a(1'h1),
        .b(_T_281)
    );
    wire _T_283;
    MUX_UNSIGNED #(.width(1)) u_mux_1431 (
        .y(_T_283),
        .sel(_T_189),
        .a(1'h1),
        .b(_T_282)
    );
    wire _T_284;
    MUX_UNSIGNED #(.width(1)) u_mux_1432 (
        .y(_T_284),
        .sel(_T_185),
        .a(1'h0),
        .b(_T_283)
    );
    wire _T_285;
    MUX_UNSIGNED #(.width(1)) u_mux_1433 (
        .y(_T_285),
        .sel(_T_181),
        .a(1'h0),
        .b(_T_284)
    );
    wire _T_286;
    MUX_UNSIGNED #(.width(1)) u_mux_1434 (
        .y(_T_286),
        .sel(_T_177),
        .a(1'h1),
        .b(_T_285)
    );
    wire _T_287;
    MUX_UNSIGNED #(.width(1)) u_mux_1435 (
        .y(_T_287),
        .sel(_T_173),
        .a(1'h1),
        .b(_T_286)
    );
    wire _T_288;
    MUX_UNSIGNED #(.width(1)) u_mux_1436 (
        .y(_T_288),
        .sel(_T_169),
        .a(1'h1),
        .b(_T_287)
    );
    wire _T_289;
    MUX_UNSIGNED #(.width(1)) u_mux_1437 (
        .y(_T_289),
        .sel(_T_165),
        .a(1'h1),
        .b(_T_288)
    );
    wire _T_290;
    MUX_UNSIGNED #(.width(1)) u_mux_1438 (
        .y(_T_290),
        .sel(_T_161),
        .a(1'h1),
        .b(_T_289)
    );
    wire _T_291;
    MUX_UNSIGNED #(.width(1)) u_mux_1439 (
        .y(_T_291),
        .sel(_T_157),
        .a(1'h1),
        .b(_T_290)
    );
    wire _T_292;
    MUX_UNSIGNED #(.width(1)) u_mux_1440 (
        .y(_T_292),
        .sel(_T_153),
        .a(1'h1),
        .b(_T_291)
    );
    wire _T_293;
    MUX_UNSIGNED #(.width(1)) u_mux_1441 (
        .y(_T_293),
        .sel(_T_149),
        .a(1'h1),
        .b(_T_292)
    );
    wire _T_294;
    MUX_UNSIGNED #(.width(1)) u_mux_1442 (
        .y(_T_294),
        .sel(_T_145),
        .a(1'h1),
        .b(_T_293)
    );
    wire _T_295;
    MUX_UNSIGNED #(.width(1)) u_mux_1443 (
        .y(_T_295),
        .sel(_T_141),
        .a(1'h1),
        .b(_T_294)
    );
    wire _T_296;
    MUX_UNSIGNED #(.width(1)) u_mux_1444 (
        .y(_T_296),
        .sel(_T_137),
        .a(1'h1),
        .b(_T_295)
    );
    wire _T_297;
    MUX_UNSIGNED #(.width(1)) u_mux_1445 (
        .y(_T_297),
        .sel(_T_133),
        .a(1'h1),
        .b(_T_296)
    );
    wire _T_298;
    MUX_UNSIGNED #(.width(1)) u_mux_1446 (
        .y(_T_298),
        .sel(_T_129),
        .a(1'h1),
        .b(_T_297)
    );
    wire _T_299;
    MUX_UNSIGNED #(.width(1)) u_mux_1447 (
        .y(_T_299),
        .sel(_T_125),
        .a(1'h1),
        .b(_T_298)
    );
    wire _T_300;
    MUX_UNSIGNED #(.width(1)) u_mux_1448 (
        .y(_T_300),
        .sel(_T_121),
        .a(1'h1),
        .b(_T_299)
    );
    wire _T_301;
    MUX_UNSIGNED #(.width(1)) u_mux_1449 (
        .y(_T_301),
        .sel(_T_117),
        .a(1'h1),
        .b(_T_300)
    );
    wire _T_302;
    MUX_UNSIGNED #(.width(1)) u_mux_1450 (
        .y(_T_302),
        .sel(_T_113),
        .a(1'h1),
        .b(_T_301)
    );
    wire _T_303;
    MUX_UNSIGNED #(.width(1)) u_mux_1451 (
        .y(_T_303),
        .sel(_T_109),
        .a(1'h1),
        .b(_T_302)
    );
    wire _T_304;
    MUX_UNSIGNED #(.width(1)) u_mux_1452 (
        .y(_T_304),
        .sel(_T_105),
        .a(1'h1),
        .b(_T_303)
    );
    wire _T_305;
    MUX_UNSIGNED #(.width(1)) u_mux_1453 (
        .y(_T_305),
        .sel(_T_101),
        .a(1'h1),
        .b(_T_304)
    );
    wire _T_306;
    MUX_UNSIGNED #(.width(1)) u_mux_1454 (
        .y(_T_306),
        .sel(_T_97),
        .a(1'h1),
        .b(_T_305)
    );
    wire _T_307;
    MUX_UNSIGNED #(.width(1)) u_mux_1455 (
        .y(_T_307),
        .sel(_T_93),
        .a(1'h1),
        .b(_T_306)
    );
    wire _T_308;
    MUX_UNSIGNED #(.width(1)) u_mux_1456 (
        .y(_T_308),
        .sel(_T_89),
        .a(1'h1),
        .b(_T_307)
    );
    wire _T_309;
    MUX_UNSIGNED #(.width(1)) u_mux_1457 (
        .y(_T_309),
        .sel(_T_85),
        .a(1'h1),
        .b(_T_308)
    );
    wire _T_310;
    MUX_UNSIGNED #(.width(1)) u_mux_1458 (
        .y(_T_310),
        .sel(_T_81),
        .a(1'h1),
        .b(_T_309)
    );
    wire _T_311;
    MUX_UNSIGNED #(.width(1)) u_mux_1459 (
        .y(_T_311),
        .sel(_T_77),
        .a(1'h1),
        .b(_T_310)
    );
    wire _T_312;
    MUX_UNSIGNED #(.width(1)) u_mux_1460 (
        .y(_T_312),
        .sel(_T_73),
        .a(1'h1),
        .b(_T_311)
    );
    wire _T_313;
    MUX_UNSIGNED #(.width(1)) u_mux_1461 (
        .y(_T_313),
        .sel(_T_69),
        .a(1'h0),
        .b(_T_312)
    );
    wire _T_314;
    MUX_UNSIGNED #(.width(1)) u_mux_1462 (
        .y(_T_314),
        .sel(_T_65),
        .a(1'h0),
        .b(_T_313)
    );
    wire _T_315;
    MUX_UNSIGNED #(.width(1)) u_mux_1463 (
        .y(_T_315),
        .sel(_T_61),
        .a(1'h0),
        .b(_T_314)
    );
    wire _T_316;
    MUX_UNSIGNED #(.width(1)) u_mux_1464 (
        .y(_T_316),
        .sel(_T_57),
        .a(1'h0),
        .b(_T_315)
    );
    wire _T_317;
    MUX_UNSIGNED #(.width(1)) u_mux_1465 (
        .y(_T_317),
        .sel(_T_53),
        .a(1'h0),
        .b(_T_316)
    );
    wire _T_318;
    MUX_UNSIGNED #(.width(1)) u_mux_1466 (
        .y(_T_318),
        .sel(_T_49),
        .a(1'h0),
        .b(_T_317)
    );
    wire _T_319;
    MUX_UNSIGNED #(.width(1)) u_mux_1467 (
        .y(_T_319),
        .sel(_T_45),
        .a(1'h1),
        .b(_T_318)
    );
    wire _T_320;
    MUX_UNSIGNED #(.width(1)) u_mux_1468 (
        .y(_T_320),
        .sel(_T_41),
        .a(1'h0),
        .b(_T_319)
    );
    wire _T_321;
    MUX_UNSIGNED #(.width(1)) u_mux_1469 (
        .y(_T_321),
        .sel(_T_37),
        .a(1'h0),
        .b(_T_320)
    );
    wire ctrlSignals_1;
    MUX_UNSIGNED #(.width(1)) u_mux_1470 (
        .y(ctrlSignals_1),
        .sel(_T_33),
        .a(1'h0),
        .b(_T_321)
    );
    wire _T_322;
    assign _T_322 = 1'h0;
    wire _T_323;
    assign _T_323 = 1'h0;
    wire _T_324;
    assign _T_324 = 1'h0;
    wire _T_325;
    assign _T_325 = 1'h0;
    wire _T_326;
    assign _T_326 = 1'h0;
    wire _T_327;
    assign _T_327 = 1'h0;
    wire _T_328;
    assign _T_328 = 1'h0;
    wire _T_329;
    assign _T_329 = 1'h0;
    wire _T_330;
    assign _T_330 = 1'h0;
    wire _T_331;
    assign _T_331 = 1'h0;
    wire _T_332;
    assign _T_332 = 1'h0;
    wire _T_333;
    assign _T_333 = 1'h0;
    wire _T_334;
    MUX_UNSIGNED #(.width(1)) u_mux_1471 (
        .y(_T_334),
        .sel(_T_177),
        .a(1'h1),
        .b(_T_333)
    );
    wire _T_335;
    MUX_UNSIGNED #(.width(1)) u_mux_1472 (
        .y(_T_335),
        .sel(_T_173),
        .a(1'h1),
        .b(_T_334)
    );
    wire _T_336;
    MUX_UNSIGNED #(.width(1)) u_mux_1473 (
        .y(_T_336),
        .sel(_T_169),
        .a(1'h1),
        .b(_T_335)
    );
    wire _T_337;
    MUX_UNSIGNED #(.width(1)) u_mux_1474 (
        .y(_T_337),
        .sel(_T_165),
        .a(1'h1),
        .b(_T_336)
    );
    wire _T_338;
    MUX_UNSIGNED #(.width(1)) u_mux_1475 (
        .y(_T_338),
        .sel(_T_161),
        .a(1'h1),
        .b(_T_337)
    );
    wire _T_339;
    MUX_UNSIGNED #(.width(1)) u_mux_1476 (
        .y(_T_339),
        .sel(_T_157),
        .a(1'h1),
        .b(_T_338)
    );
    wire _T_340;
    MUX_UNSIGNED #(.width(1)) u_mux_1477 (
        .y(_T_340),
        .sel(_T_153),
        .a(1'h1),
        .b(_T_339)
    );
    wire _T_341;
    MUX_UNSIGNED #(.width(1)) u_mux_1478 (
        .y(_T_341),
        .sel(_T_149),
        .a(1'h1),
        .b(_T_340)
    );
    wire _T_342;
    MUX_UNSIGNED #(.width(1)) u_mux_1479 (
        .y(_T_342),
        .sel(_T_145),
        .a(1'h1),
        .b(_T_341)
    );
    wire _T_343;
    MUX_UNSIGNED #(.width(1)) u_mux_1480 (
        .y(_T_343),
        .sel(_T_141),
        .a(1'h1),
        .b(_T_342)
    );
    wire _T_344;
    MUX_UNSIGNED #(.width(1)) u_mux_1481 (
        .y(_T_344),
        .sel(_T_137),
        .a(1'h0),
        .b(_T_343)
    );
    wire _T_345;
    MUX_UNSIGNED #(.width(1)) u_mux_1482 (
        .y(_T_345),
        .sel(_T_133),
        .a(1'h0),
        .b(_T_344)
    );
    wire _T_346;
    MUX_UNSIGNED #(.width(1)) u_mux_1483 (
        .y(_T_346),
        .sel(_T_129),
        .a(1'h0),
        .b(_T_345)
    );
    wire _T_347;
    MUX_UNSIGNED #(.width(1)) u_mux_1484 (
        .y(_T_347),
        .sel(_T_125),
        .a(1'h0),
        .b(_T_346)
    );
    wire _T_348;
    MUX_UNSIGNED #(.width(1)) u_mux_1485 (
        .y(_T_348),
        .sel(_T_121),
        .a(1'h0),
        .b(_T_347)
    );
    wire _T_349;
    MUX_UNSIGNED #(.width(1)) u_mux_1486 (
        .y(_T_349),
        .sel(_T_117),
        .a(1'h0),
        .b(_T_348)
    );
    wire _T_350;
    MUX_UNSIGNED #(.width(1)) u_mux_1487 (
        .y(_T_350),
        .sel(_T_113),
        .a(1'h0),
        .b(_T_349)
    );
    wire _T_351;
    MUX_UNSIGNED #(.width(1)) u_mux_1488 (
        .y(_T_351),
        .sel(_T_109),
        .a(1'h0),
        .b(_T_350)
    );
    wire _T_352;
    MUX_UNSIGNED #(.width(1)) u_mux_1489 (
        .y(_T_352),
        .sel(_T_105),
        .a(1'h0),
        .b(_T_351)
    );
    wire _T_353;
    MUX_UNSIGNED #(.width(1)) u_mux_1490 (
        .y(_T_353),
        .sel(_T_101),
        .a(1'h0),
        .b(_T_352)
    );
    wire _T_354;
    MUX_UNSIGNED #(.width(1)) u_mux_1491 (
        .y(_T_354),
        .sel(_T_97),
        .a(1'h0),
        .b(_T_353)
    );
    wire _T_355;
    MUX_UNSIGNED #(.width(1)) u_mux_1492 (
        .y(_T_355),
        .sel(_T_93),
        .a(1'h0),
        .b(_T_354)
    );
    wire _T_356;
    MUX_UNSIGNED #(.width(1)) u_mux_1493 (
        .y(_T_356),
        .sel(_T_89),
        .a(1'h0),
        .b(_T_355)
    );
    wire _T_357;
    MUX_UNSIGNED #(.width(1)) u_mux_1494 (
        .y(_T_357),
        .sel(_T_85),
        .a(1'h0),
        .b(_T_356)
    );
    wire _T_358;
    MUX_UNSIGNED #(.width(1)) u_mux_1495 (
        .y(_T_358),
        .sel(_T_81),
        .a(1'h0),
        .b(_T_357)
    );
    wire _T_359;
    MUX_UNSIGNED #(.width(1)) u_mux_1496 (
        .y(_T_359),
        .sel(_T_77),
        .a(1'h0),
        .b(_T_358)
    );
    wire _T_360;
    MUX_UNSIGNED #(.width(1)) u_mux_1497 (
        .y(_T_360),
        .sel(_T_73),
        .a(1'h0),
        .b(_T_359)
    );
    wire _T_361;
    MUX_UNSIGNED #(.width(1)) u_mux_1498 (
        .y(_T_361),
        .sel(_T_69),
        .a(1'h0),
        .b(_T_360)
    );
    wire _T_362;
    MUX_UNSIGNED #(.width(1)) u_mux_1499 (
        .y(_T_362),
        .sel(_T_65),
        .a(1'h0),
        .b(_T_361)
    );
    wire _T_363;
    MUX_UNSIGNED #(.width(1)) u_mux_1500 (
        .y(_T_363),
        .sel(_T_61),
        .a(1'h0),
        .b(_T_362)
    );
    wire _T_364;
    MUX_UNSIGNED #(.width(1)) u_mux_1501 (
        .y(_T_364),
        .sel(_T_57),
        .a(1'h0),
        .b(_T_363)
    );
    wire _T_365;
    MUX_UNSIGNED #(.width(1)) u_mux_1502 (
        .y(_T_365),
        .sel(_T_53),
        .a(1'h0),
        .b(_T_364)
    );
    wire _T_366;
    MUX_UNSIGNED #(.width(1)) u_mux_1503 (
        .y(_T_366),
        .sel(_T_49),
        .a(1'h0),
        .b(_T_365)
    );
    wire _T_367;
    MUX_UNSIGNED #(.width(1)) u_mux_1504 (
        .y(_T_367),
        .sel(_T_45),
        .a(1'h0),
        .b(_T_366)
    );
    wire _T_368;
    MUX_UNSIGNED #(.width(1)) u_mux_1505 (
        .y(_T_368),
        .sel(_T_41),
        .a(1'h0),
        .b(_T_367)
    );
    wire _T_369;
    MUX_UNSIGNED #(.width(1)) u_mux_1506 (
        .y(_T_369),
        .sel(_T_37),
        .a(1'h0),
        .b(_T_368)
    );
    wire ctrlSignals_2;
    MUX_UNSIGNED #(.width(1)) u_mux_1507 (
        .y(ctrlSignals_2),
        .sel(_T_33),
        .a(1'h0),
        .b(_T_369)
    );
    wire [2:0] _T_370;
    assign _T_370 = 3'h0;
    wire [2:0] _T_371;
    assign _T_371 = 3'h0;
    wire [2:0] _T_372;
    assign _T_372 = 3'h0;
    wire [2:0] _T_373;
    assign _T_373 = 3'h0;
    wire [2:0] _T_374;
    MUX_UNSIGNED #(.width(3)) u_mux_1508 (
        .y(_T_374),
        .sel(_T_209),
        .a(3'h6),
        .b(_T_373)
    );
    wire [2:0] _T_375;
    MUX_UNSIGNED #(.width(3)) u_mux_1509 (
        .y(_T_375),
        .sel(_T_205),
        .a(3'h6),
        .b(_T_374)
    );
    wire [2:0] _T_376;
    MUX_UNSIGNED #(.width(3)) u_mux_1510 (
        .y(_T_376),
        .sel(_T_201),
        .a(3'h6),
        .b(_T_375)
    );
    wire [2:0] _T_377;
    MUX_UNSIGNED #(.width(3)) u_mux_1511 (
        .y(_T_377),
        .sel(_T_197),
        .a(3'h0),
        .b(_T_376)
    );
    wire [2:0] _T_378;
    MUX_UNSIGNED #(.width(3)) u_mux_1512 (
        .y(_T_378),
        .sel(_T_193),
        .a(3'h0),
        .b(_T_377)
    );
    wire [2:0] _T_379;
    MUX_UNSIGNED #(.width(3)) u_mux_1513 (
        .y(_T_379),
        .sel(_T_189),
        .a(3'h0),
        .b(_T_378)
    );
    wire [2:0] _T_380;
    MUX_UNSIGNED #(.width(3)) u_mux_1514 (
        .y(_T_380),
        .sel(_T_185),
        .a(3'h0),
        .b(_T_379)
    );
    wire [2:0] _T_381;
    MUX_UNSIGNED #(.width(3)) u_mux_1515 (
        .y(_T_381),
        .sel(_T_181),
        .a(3'h0),
        .b(_T_380)
    );
    wire [2:0] _T_382;
    MUX_UNSIGNED #(.width(3)) u_mux_1516 (
        .y(_T_382),
        .sel(_T_177),
        .a(3'h0),
        .b(_T_381)
    );
    wire [2:0] _T_383;
    MUX_UNSIGNED #(.width(3)) u_mux_1517 (
        .y(_T_383),
        .sel(_T_173),
        .a(3'h0),
        .b(_T_382)
    );
    wire [2:0] _T_384;
    MUX_UNSIGNED #(.width(3)) u_mux_1518 (
        .y(_T_384),
        .sel(_T_169),
        .a(3'h0),
        .b(_T_383)
    );
    wire [2:0] _T_385;
    MUX_UNSIGNED #(.width(3)) u_mux_1519 (
        .y(_T_385),
        .sel(_T_165),
        .a(3'h0),
        .b(_T_384)
    );
    wire [2:0] _T_386;
    MUX_UNSIGNED #(.width(3)) u_mux_1520 (
        .y(_T_386),
        .sel(_T_161),
        .a(3'h0),
        .b(_T_385)
    );
    wire [2:0] _T_387;
    MUX_UNSIGNED #(.width(3)) u_mux_1521 (
        .y(_T_387),
        .sel(_T_157),
        .a(3'h0),
        .b(_T_386)
    );
    wire [2:0] _T_388;
    MUX_UNSIGNED #(.width(3)) u_mux_1522 (
        .y(_T_388),
        .sel(_T_153),
        .a(3'h0),
        .b(_T_387)
    );
    wire [2:0] _T_389;
    MUX_UNSIGNED #(.width(3)) u_mux_1523 (
        .y(_T_389),
        .sel(_T_149),
        .a(3'h0),
        .b(_T_388)
    );
    wire [2:0] _T_390;
    MUX_UNSIGNED #(.width(3)) u_mux_1524 (
        .y(_T_390),
        .sel(_T_145),
        .a(3'h0),
        .b(_T_389)
    );
    wire [2:0] _T_391;
    MUX_UNSIGNED #(.width(3)) u_mux_1525 (
        .y(_T_391),
        .sel(_T_141),
        .a(3'h0),
        .b(_T_390)
    );
    wire [2:0] _T_392;
    MUX_UNSIGNED #(.width(3)) u_mux_1526 (
        .y(_T_392),
        .sel(_T_137),
        .a(3'h1),
        .b(_T_391)
    );
    wire [2:0] _T_393;
    MUX_UNSIGNED #(.width(3)) u_mux_1527 (
        .y(_T_393),
        .sel(_T_133),
        .a(3'h1),
        .b(_T_392)
    );
    wire [2:0] _T_394;
    MUX_UNSIGNED #(.width(3)) u_mux_1528 (
        .y(_T_394),
        .sel(_T_129),
        .a(3'h1),
        .b(_T_393)
    );
    wire [2:0] _T_395;
    MUX_UNSIGNED #(.width(3)) u_mux_1529 (
        .y(_T_395),
        .sel(_T_125),
        .a(3'h1),
        .b(_T_394)
    );
    wire [2:0] _T_396;
    MUX_UNSIGNED #(.width(3)) u_mux_1530 (
        .y(_T_396),
        .sel(_T_121),
        .a(3'h1),
        .b(_T_395)
    );
    wire [2:0] _T_397;
    MUX_UNSIGNED #(.width(3)) u_mux_1531 (
        .y(_T_397),
        .sel(_T_117),
        .a(3'h1),
        .b(_T_396)
    );
    wire [2:0] _T_398;
    MUX_UNSIGNED #(.width(3)) u_mux_1532 (
        .y(_T_398),
        .sel(_T_113),
        .a(3'h1),
        .b(_T_397)
    );
    wire [2:0] _T_399;
    MUX_UNSIGNED #(.width(3)) u_mux_1533 (
        .y(_T_399),
        .sel(_T_109),
        .a(3'h1),
        .b(_T_398)
    );
    wire [2:0] _T_400;
    MUX_UNSIGNED #(.width(3)) u_mux_1534 (
        .y(_T_400),
        .sel(_T_105),
        .a(3'h1),
        .b(_T_399)
    );
    wire [2:0] _T_401;
    MUX_UNSIGNED #(.width(3)) u_mux_1535 (
        .y(_T_401),
        .sel(_T_101),
        .a(3'h2),
        .b(_T_400)
    );
    wire [2:0] _T_402;
    MUX_UNSIGNED #(.width(3)) u_mux_1536 (
        .y(_T_402),
        .sel(_T_97),
        .a(3'h2),
        .b(_T_401)
    );
    wire [2:0] _T_403;
    MUX_UNSIGNED #(.width(3)) u_mux_1537 (
        .y(_T_403),
        .sel(_T_93),
        .a(3'h2),
        .b(_T_402)
    );
    wire [2:0] _T_404;
    MUX_UNSIGNED #(.width(3)) u_mux_1538 (
        .y(_T_404),
        .sel(_T_89),
        .a(3'h1),
        .b(_T_403)
    );
    wire [2:0] _T_405;
    MUX_UNSIGNED #(.width(3)) u_mux_1539 (
        .y(_T_405),
        .sel(_T_85),
        .a(3'h1),
        .b(_T_404)
    );
    wire [2:0] _T_406;
    MUX_UNSIGNED #(.width(3)) u_mux_1540 (
        .y(_T_406),
        .sel(_T_81),
        .a(3'h1),
        .b(_T_405)
    );
    wire [2:0] _T_407;
    MUX_UNSIGNED #(.width(3)) u_mux_1541 (
        .y(_T_407),
        .sel(_T_77),
        .a(3'h1),
        .b(_T_406)
    );
    wire [2:0] _T_408;
    MUX_UNSIGNED #(.width(3)) u_mux_1542 (
        .y(_T_408),
        .sel(_T_73),
        .a(3'h1),
        .b(_T_407)
    );
    wire [2:0] _T_409;
    MUX_UNSIGNED #(.width(3)) u_mux_1543 (
        .y(_T_409),
        .sel(_T_69),
        .a(3'h5),
        .b(_T_408)
    );
    wire [2:0] _T_410;
    MUX_UNSIGNED #(.width(3)) u_mux_1544 (
        .y(_T_410),
        .sel(_T_65),
        .a(3'h5),
        .b(_T_409)
    );
    wire [2:0] _T_411;
    MUX_UNSIGNED #(.width(3)) u_mux_1545 (
        .y(_T_411),
        .sel(_T_61),
        .a(3'h5),
        .b(_T_410)
    );
    wire [2:0] _T_412;
    MUX_UNSIGNED #(.width(3)) u_mux_1546 (
        .y(_T_412),
        .sel(_T_57),
        .a(3'h5),
        .b(_T_411)
    );
    wire [2:0] _T_413;
    MUX_UNSIGNED #(.width(3)) u_mux_1547 (
        .y(_T_413),
        .sel(_T_53),
        .a(3'h5),
        .b(_T_412)
    );
    wire [2:0] _T_414;
    MUX_UNSIGNED #(.width(3)) u_mux_1548 (
        .y(_T_414),
        .sel(_T_49),
        .a(3'h5),
        .b(_T_413)
    );
    wire [2:0] _T_415;
    MUX_UNSIGNED #(.width(3)) u_mux_1549 (
        .y(_T_415),
        .sel(_T_45),
        .a(3'h1),
        .b(_T_414)
    );
    wire [2:0] _T_416;
    MUX_UNSIGNED #(.width(3)) u_mux_1550 (
        .y(_T_416),
        .sel(_T_41),
        .a(3'h4),
        .b(_T_415)
    );
    wire [2:0] _T_417;
    MUX_UNSIGNED #(.width(3)) u_mux_1551 (
        .y(_T_417),
        .sel(_T_37),
        .a(3'h3),
        .b(_T_416)
    );
    wire [2:0] ctrlSignals_3;
    MUX_UNSIGNED #(.width(3)) u_mux_1552 (
        .y(ctrlSignals_3),
        .sel(_T_33),
        .a(3'h3),
        .b(_T_417)
    );
    wire [3:0] _T_418;
    assign _T_418 = 4'hF;
    wire [3:0] _T_419;
    assign _T_419 = 4'hF;
    wire [3:0] _T_420;
    assign _T_420 = 4'hF;
    wire [3:0] _T_421;
    assign _T_421 = 4'hF;
    wire [3:0] _T_422;
    assign _T_422 = 4'hF;
    wire [3:0] _T_423;
    assign _T_423 = 4'hF;
    wire [3:0] _T_424;
    assign _T_424 = 4'hF;
    wire [3:0] _T_425;
    MUX_UNSIGNED #(.width(4)) u_mux_1553 (
        .y(_T_425),
        .sel(_T_197),
        .a(4'hA),
        .b(_T_424)
    );
    wire [3:0] _T_426;
    MUX_UNSIGNED #(.width(4)) u_mux_1554 (
        .y(_T_426),
        .sel(_T_193),
        .a(4'hA),
        .b(_T_425)
    );
    wire [3:0] _T_427;
    MUX_UNSIGNED #(.width(4)) u_mux_1555 (
        .y(_T_427),
        .sel(_T_189),
        .a(4'hA),
        .b(_T_426)
    );
    wire [3:0] _T_428;
    MUX_UNSIGNED #(.width(4)) u_mux_1556 (
        .y(_T_428),
        .sel(_T_185),
        .a(4'hF),
        .b(_T_427)
    );
    wire [3:0] _T_429;
    MUX_UNSIGNED #(.width(4)) u_mux_1557 (
        .y(_T_429),
        .sel(_T_181),
        .a(4'hF),
        .b(_T_428)
    );
    wire [3:0] _T_430;
    MUX_UNSIGNED #(.width(4)) u_mux_1558 (
        .y(_T_430),
        .sel(_T_177),
        .a(4'h2),
        .b(_T_429)
    );
    wire [3:0] _T_431;
    MUX_UNSIGNED #(.width(4)) u_mux_1559 (
        .y(_T_431),
        .sel(_T_173),
        .a(4'h3),
        .b(_T_430)
    );
    wire [3:0] _T_432;
    MUX_UNSIGNED #(.width(4)) u_mux_1560 (
        .y(_T_432),
        .sel(_T_169),
        .a(4'h9),
        .b(_T_431)
    );
    wire [3:0] _T_433;
    MUX_UNSIGNED #(.width(4)) u_mux_1561 (
        .y(_T_433),
        .sel(_T_165),
        .a(4'h8),
        .b(_T_432)
    );
    wire [3:0] _T_434;
    MUX_UNSIGNED #(.width(4)) u_mux_1562 (
        .y(_T_434),
        .sel(_T_161),
        .a(4'h4),
        .b(_T_433)
    );
    wire [3:0] _T_435;
    MUX_UNSIGNED #(.width(4)) u_mux_1563 (
        .y(_T_435),
        .sel(_T_157),
        .a(4'h7),
        .b(_T_434)
    );
    wire [3:0] _T_436;
    MUX_UNSIGNED #(.width(4)) u_mux_1564 (
        .y(_T_436),
        .sel(_T_153),
        .a(4'h5),
        .b(_T_435)
    );
    wire [3:0] _T_437;
    MUX_UNSIGNED #(.width(4)) u_mux_1565 (
        .y(_T_437),
        .sel(_T_149),
        .a(4'h6),
        .b(_T_436)
    );
    wire [3:0] _T_438;
    MUX_UNSIGNED #(.width(4)) u_mux_1566 (
        .y(_T_438),
        .sel(_T_145),
        .a(4'h1),
        .b(_T_437)
    );
    wire [3:0] _T_439;
    MUX_UNSIGNED #(.width(4)) u_mux_1567 (
        .y(_T_439),
        .sel(_T_141),
        .a(4'h0),
        .b(_T_438)
    );
    wire [3:0] _T_440;
    MUX_UNSIGNED #(.width(4)) u_mux_1568 (
        .y(_T_440),
        .sel(_T_137),
        .a(4'h9),
        .b(_T_439)
    );
    wire [3:0] _T_441;
    MUX_UNSIGNED #(.width(4)) u_mux_1569 (
        .y(_T_441),
        .sel(_T_133),
        .a(4'h8),
        .b(_T_440)
    );
    wire [3:0] _T_442;
    MUX_UNSIGNED #(.width(4)) u_mux_1570 (
        .y(_T_442),
        .sel(_T_129),
        .a(4'h6),
        .b(_T_441)
    );
    wire [3:0] _T_443;
    MUX_UNSIGNED #(.width(4)) u_mux_1571 (
        .y(_T_443),
        .sel(_T_125),
        .a(4'h2),
        .b(_T_442)
    );
    wire [3:0] _T_444;
    MUX_UNSIGNED #(.width(4)) u_mux_1572 (
        .y(_T_444),
        .sel(_T_121),
        .a(4'h3),
        .b(_T_443)
    );
    wire [3:0] _T_445;
    MUX_UNSIGNED #(.width(4)) u_mux_1573 (
        .y(_T_445),
        .sel(_T_117),
        .a(4'h4),
        .b(_T_444)
    );
    wire [3:0] _T_446;
    MUX_UNSIGNED #(.width(4)) u_mux_1574 (
        .y(_T_446),
        .sel(_T_113),
        .a(4'h7),
        .b(_T_445)
    );
    wire [3:0] _T_447;
    MUX_UNSIGNED #(.width(4)) u_mux_1575 (
        .y(_T_447),
        .sel(_T_109),
        .a(4'h5),
        .b(_T_446)
    );
    wire [3:0] _T_448;
    MUX_UNSIGNED #(.width(4)) u_mux_1576 (
        .y(_T_448),
        .sel(_T_105),
        .a(4'h0),
        .b(_T_447)
    );
    wire [3:0] _T_449;
    MUX_UNSIGNED #(.width(4)) u_mux_1577 (
        .y(_T_449),
        .sel(_T_101),
        .a(4'h0),
        .b(_T_448)
    );
    wire [3:0] _T_450;
    MUX_UNSIGNED #(.width(4)) u_mux_1578 (
        .y(_T_450),
        .sel(_T_97),
        .a(4'h0),
        .b(_T_449)
    );
    wire [3:0] _T_451;
    MUX_UNSIGNED #(.width(4)) u_mux_1579 (
        .y(_T_451),
        .sel(_T_93),
        .a(4'h0),
        .b(_T_450)
    );
    wire [3:0] _T_452;
    MUX_UNSIGNED #(.width(4)) u_mux_1580 (
        .y(_T_452),
        .sel(_T_89),
        .a(4'h0),
        .b(_T_451)
    );
    wire [3:0] _T_453;
    MUX_UNSIGNED #(.width(4)) u_mux_1581 (
        .y(_T_453),
        .sel(_T_85),
        .a(4'h0),
        .b(_T_452)
    );
    wire [3:0] _T_454;
    MUX_UNSIGNED #(.width(4)) u_mux_1582 (
        .y(_T_454),
        .sel(_T_81),
        .a(4'h0),
        .b(_T_453)
    );
    wire [3:0] _T_455;
    MUX_UNSIGNED #(.width(4)) u_mux_1583 (
        .y(_T_455),
        .sel(_T_77),
        .a(4'h0),
        .b(_T_454)
    );
    wire [3:0] _T_456;
    MUX_UNSIGNED #(.width(4)) u_mux_1584 (
        .y(_T_456),
        .sel(_T_73),
        .a(4'h0),
        .b(_T_455)
    );
    wire [3:0] _T_457;
    MUX_UNSIGNED #(.width(4)) u_mux_1585 (
        .y(_T_457),
        .sel(_T_69),
        .a(4'h0),
        .b(_T_456)
    );
    wire [3:0] _T_458;
    MUX_UNSIGNED #(.width(4)) u_mux_1586 (
        .y(_T_458),
        .sel(_T_65),
        .a(4'h0),
        .b(_T_457)
    );
    wire [3:0] _T_459;
    MUX_UNSIGNED #(.width(4)) u_mux_1587 (
        .y(_T_459),
        .sel(_T_61),
        .a(4'h0),
        .b(_T_458)
    );
    wire [3:0] _T_460;
    MUX_UNSIGNED #(.width(4)) u_mux_1588 (
        .y(_T_460),
        .sel(_T_57),
        .a(4'h0),
        .b(_T_459)
    );
    wire [3:0] _T_461;
    MUX_UNSIGNED #(.width(4)) u_mux_1589 (
        .y(_T_461),
        .sel(_T_53),
        .a(4'h0),
        .b(_T_460)
    );
    wire [3:0] _T_462;
    MUX_UNSIGNED #(.width(4)) u_mux_1590 (
        .y(_T_462),
        .sel(_T_49),
        .a(4'h0),
        .b(_T_461)
    );
    wire [3:0] _T_463;
    MUX_UNSIGNED #(.width(4)) u_mux_1591 (
        .y(_T_463),
        .sel(_T_45),
        .a(4'h0),
        .b(_T_462)
    );
    wire [3:0] _T_464;
    MUX_UNSIGNED #(.width(4)) u_mux_1592 (
        .y(_T_464),
        .sel(_T_41),
        .a(4'h0),
        .b(_T_463)
    );
    wire [3:0] _T_465;
    MUX_UNSIGNED #(.width(4)) u_mux_1593 (
        .y(_T_465),
        .sel(_T_37),
        .a(4'h0),
        .b(_T_464)
    );
    wire [3:0] ctrlSignals_4;
    MUX_UNSIGNED #(.width(4)) u_mux_1594 (
        .y(ctrlSignals_4),
        .sel(_T_33),
        .a(4'hB),
        .b(_T_465)
    );
    wire [2:0] _T_466;
    assign _T_466 = 3'h0;
    wire [2:0] _T_467;
    assign _T_467 = 3'h0;
    wire [2:0] _T_468;
    assign _T_468 = 3'h0;
    wire [2:0] _T_469;
    assign _T_469 = 3'h0;
    wire [2:0] _T_470;
    assign _T_470 = 3'h0;
    wire [2:0] _T_471;
    assign _T_471 = 3'h0;
    wire [2:0] _T_472;
    assign _T_472 = 3'h0;
    wire [2:0] _T_473;
    assign _T_473 = 3'h0;
    wire [2:0] _T_474;
    assign _T_474 = 3'h0;
    wire [2:0] _T_475;
    assign _T_475 = 3'h0;
    wire [2:0] _T_476;
    assign _T_476 = 3'h0;
    wire [2:0] _T_477;
    assign _T_477 = 3'h0;
    wire [2:0] _T_478;
    assign _T_478 = 3'h0;
    wire [2:0] _T_479;
    assign _T_479 = 3'h0;
    wire [2:0] _T_480;
    assign _T_480 = 3'h0;
    wire [2:0] _T_481;
    assign _T_481 = 3'h0;
    wire [2:0] _T_482;
    assign _T_482 = 3'h0;
    wire [2:0] _T_483;
    assign _T_483 = 3'h0;
    wire [2:0] _T_484;
    assign _T_484 = 3'h0;
    wire [2:0] _T_485;
    assign _T_485 = 3'h0;
    wire [2:0] _T_486;
    assign _T_486 = 3'h0;
    wire [2:0] _T_487;
    assign _T_487 = 3'h0;
    wire [2:0] _T_488;
    assign _T_488 = 3'h0;
    wire [2:0] _T_489;
    assign _T_489 = 3'h0;
    wire [2:0] _T_490;
    assign _T_490 = 3'h0;
    wire [2:0] _T_491;
    assign _T_491 = 3'h0;
    wire [2:0] _T_492;
    assign _T_492 = 3'h0;
    wire [2:0] _T_493;
    assign _T_493 = 3'h0;
    wire [2:0] _T_494;
    assign _T_494 = 3'h0;
    wire [2:0] _T_495;
    assign _T_495 = 3'h0;
    wire [2:0] _T_496;
    assign _T_496 = 3'h0;
    wire [2:0] _T_497;
    assign _T_497 = 3'h0;
    wire [2:0] _T_498;
    assign _T_498 = 3'h0;
    wire [2:0] _T_499;
    assign _T_499 = 3'h0;
    wire [2:0] _T_500;
    assign _T_500 = 3'h0;
    wire [2:0] _T_501;
    assign _T_501 = 3'h0;
    wire [2:0] _T_502;
    assign _T_502 = 3'h0;
    wire [2:0] _T_503;
    assign _T_503 = 3'h0;
    wire [2:0] _T_504;
    assign _T_504 = 3'h0;
    wire [2:0] _T_505;
    MUX_UNSIGNED #(.width(3)) u_mux_1595 (
        .y(_T_505),
        .sel(_T_69),
        .a(3'h4),
        .b(_T_504)
    );
    wire [2:0] _T_506;
    MUX_UNSIGNED #(.width(3)) u_mux_1596 (
        .y(_T_506),
        .sel(_T_65),
        .a(3'h1),
        .b(_T_505)
    );
    wire [2:0] _T_507;
    MUX_UNSIGNED #(.width(3)) u_mux_1597 (
        .y(_T_507),
        .sel(_T_61),
        .a(3'h5),
        .b(_T_506)
    );
    wire [2:0] _T_508;
    MUX_UNSIGNED #(.width(3)) u_mux_1598 (
        .y(_T_508),
        .sel(_T_57),
        .a(3'h2),
        .b(_T_507)
    );
    wire [2:0] _T_509;
    MUX_UNSIGNED #(.width(3)) u_mux_1599 (
        .y(_T_509),
        .sel(_T_53),
        .a(3'h6),
        .b(_T_508)
    );
    wire [2:0] _T_510;
    MUX_UNSIGNED #(.width(3)) u_mux_1600 (
        .y(_T_510),
        .sel(_T_49),
        .a(3'h3),
        .b(_T_509)
    );
    wire [2:0] _T_511;
    MUX_UNSIGNED #(.width(3)) u_mux_1601 (
        .y(_T_511),
        .sel(_T_45),
        .a(3'h0),
        .b(_T_510)
    );
    wire [2:0] _T_512;
    MUX_UNSIGNED #(.width(3)) u_mux_1602 (
        .y(_T_512),
        .sel(_T_41),
        .a(3'h0),
        .b(_T_511)
    );
    wire [2:0] _T_513;
    MUX_UNSIGNED #(.width(3)) u_mux_1603 (
        .y(_T_513),
        .sel(_T_37),
        .a(3'h0),
        .b(_T_512)
    );
    wire [2:0] ctrlSignals_5;
    MUX_UNSIGNED #(.width(3)) u_mux_1604 (
        .y(ctrlSignals_5),
        .sel(_T_33),
        .a(3'h0),
        .b(_T_513)
    );
    wire _T_514;
    assign _T_514 = 1'h0;
    wire _T_515;
    MUX_UNSIGNED #(.width(1)) u_mux_1605 (
        .y(_T_515),
        .sel(_T_221),
        .a(1'h1),
        .b(_T_514)
    );
    wire _T_516;
    MUX_UNSIGNED #(.width(1)) u_mux_1606 (
        .y(_T_516),
        .sel(_T_217),
        .a(1'h0),
        .b(_T_515)
    );
    wire _T_517;
    MUX_UNSIGNED #(.width(1)) u_mux_1607 (
        .y(_T_517),
        .sel(_T_213),
        .a(1'h0),
        .b(_T_516)
    );
    wire _T_518;
    MUX_UNSIGNED #(.width(1)) u_mux_1608 (
        .y(_T_518),
        .sel(_T_209),
        .a(1'h1),
        .b(_T_517)
    );
    wire _T_519;
    MUX_UNSIGNED #(.width(1)) u_mux_1609 (
        .y(_T_519),
        .sel(_T_205),
        .a(1'h1),
        .b(_T_518)
    );
    wire _T_520;
    MUX_UNSIGNED #(.width(1)) u_mux_1610 (
        .y(_T_520),
        .sel(_T_201),
        .a(1'h1),
        .b(_T_519)
    );
    wire _T_521;
    MUX_UNSIGNED #(.width(1)) u_mux_1611 (
        .y(_T_521),
        .sel(_T_197),
        .a(1'h1),
        .b(_T_520)
    );
    wire _T_522;
    MUX_UNSIGNED #(.width(1)) u_mux_1612 (
        .y(_T_522),
        .sel(_T_193),
        .a(1'h1),
        .b(_T_521)
    );
    wire _T_523;
    MUX_UNSIGNED #(.width(1)) u_mux_1613 (
        .y(_T_523),
        .sel(_T_189),
        .a(1'h1),
        .b(_T_522)
    );
    wire _T_524;
    MUX_UNSIGNED #(.width(1)) u_mux_1614 (
        .y(_T_524),
        .sel(_T_185),
        .a(1'h1),
        .b(_T_523)
    );
    wire _T_525;
    MUX_UNSIGNED #(.width(1)) u_mux_1615 (
        .y(_T_525),
        .sel(_T_181),
        .a(1'h0),
        .b(_T_524)
    );
    wire _T_526;
    MUX_UNSIGNED #(.width(1)) u_mux_1616 (
        .y(_T_526),
        .sel(_T_177),
        .a(1'h0),
        .b(_T_525)
    );
    wire _T_527;
    MUX_UNSIGNED #(.width(1)) u_mux_1617 (
        .y(_T_527),
        .sel(_T_173),
        .a(1'h0),
        .b(_T_526)
    );
    wire _T_528;
    MUX_UNSIGNED #(.width(1)) u_mux_1618 (
        .y(_T_528),
        .sel(_T_169),
        .a(1'h0),
        .b(_T_527)
    );
    wire _T_529;
    MUX_UNSIGNED #(.width(1)) u_mux_1619 (
        .y(_T_529),
        .sel(_T_165),
        .a(1'h0),
        .b(_T_528)
    );
    wire _T_530;
    MUX_UNSIGNED #(.width(1)) u_mux_1620 (
        .y(_T_530),
        .sel(_T_161),
        .a(1'h0),
        .b(_T_529)
    );
    wire _T_531;
    MUX_UNSIGNED #(.width(1)) u_mux_1621 (
        .y(_T_531),
        .sel(_T_157),
        .a(1'h0),
        .b(_T_530)
    );
    wire _T_532;
    MUX_UNSIGNED #(.width(1)) u_mux_1622 (
        .y(_T_532),
        .sel(_T_153),
        .a(1'h0),
        .b(_T_531)
    );
    wire _T_533;
    MUX_UNSIGNED #(.width(1)) u_mux_1623 (
        .y(_T_533),
        .sel(_T_149),
        .a(1'h0),
        .b(_T_532)
    );
    wire _T_534;
    MUX_UNSIGNED #(.width(1)) u_mux_1624 (
        .y(_T_534),
        .sel(_T_145),
        .a(1'h0),
        .b(_T_533)
    );
    wire _T_535;
    MUX_UNSIGNED #(.width(1)) u_mux_1625 (
        .y(_T_535),
        .sel(_T_141),
        .a(1'h0),
        .b(_T_534)
    );
    wire _T_536;
    MUX_UNSIGNED #(.width(1)) u_mux_1626 (
        .y(_T_536),
        .sel(_T_137),
        .a(1'h0),
        .b(_T_535)
    );
    wire _T_537;
    MUX_UNSIGNED #(.width(1)) u_mux_1627 (
        .y(_T_537),
        .sel(_T_133),
        .a(1'h0),
        .b(_T_536)
    );
    wire _T_538;
    MUX_UNSIGNED #(.width(1)) u_mux_1628 (
        .y(_T_538),
        .sel(_T_129),
        .a(1'h0),
        .b(_T_537)
    );
    wire _T_539;
    MUX_UNSIGNED #(.width(1)) u_mux_1629 (
        .y(_T_539),
        .sel(_T_125),
        .a(1'h0),
        .b(_T_538)
    );
    wire _T_540;
    MUX_UNSIGNED #(.width(1)) u_mux_1630 (
        .y(_T_540),
        .sel(_T_121),
        .a(1'h0),
        .b(_T_539)
    );
    wire _T_541;
    MUX_UNSIGNED #(.width(1)) u_mux_1631 (
        .y(_T_541),
        .sel(_T_117),
        .a(1'h0),
        .b(_T_540)
    );
    wire _T_542;
    MUX_UNSIGNED #(.width(1)) u_mux_1632 (
        .y(_T_542),
        .sel(_T_113),
        .a(1'h0),
        .b(_T_541)
    );
    wire _T_543;
    MUX_UNSIGNED #(.width(1)) u_mux_1633 (
        .y(_T_543),
        .sel(_T_109),
        .a(1'h0),
        .b(_T_542)
    );
    wire _T_544;
    MUX_UNSIGNED #(.width(1)) u_mux_1634 (
        .y(_T_544),
        .sel(_T_105),
        .a(1'h0),
        .b(_T_543)
    );
    wire _T_545;
    MUX_UNSIGNED #(.width(1)) u_mux_1635 (
        .y(_T_545),
        .sel(_T_101),
        .a(1'h0),
        .b(_T_544)
    );
    wire _T_546;
    MUX_UNSIGNED #(.width(1)) u_mux_1636 (
        .y(_T_546),
        .sel(_T_97),
        .a(1'h0),
        .b(_T_545)
    );
    wire _T_547;
    MUX_UNSIGNED #(.width(1)) u_mux_1637 (
        .y(_T_547),
        .sel(_T_93),
        .a(1'h0),
        .b(_T_546)
    );
    wire _T_548;
    MUX_UNSIGNED #(.width(1)) u_mux_1638 (
        .y(_T_548),
        .sel(_T_89),
        .a(1'h1),
        .b(_T_547)
    );
    wire _T_549;
    MUX_UNSIGNED #(.width(1)) u_mux_1639 (
        .y(_T_549),
        .sel(_T_85),
        .a(1'h1),
        .b(_T_548)
    );
    wire _T_550;
    MUX_UNSIGNED #(.width(1)) u_mux_1640 (
        .y(_T_550),
        .sel(_T_81),
        .a(1'h1),
        .b(_T_549)
    );
    wire _T_551;
    MUX_UNSIGNED #(.width(1)) u_mux_1641 (
        .y(_T_551),
        .sel(_T_77),
        .a(1'h1),
        .b(_T_550)
    );
    wire _T_552;
    MUX_UNSIGNED #(.width(1)) u_mux_1642 (
        .y(_T_552),
        .sel(_T_73),
        .a(1'h1),
        .b(_T_551)
    );
    wire _T_553;
    MUX_UNSIGNED #(.width(1)) u_mux_1643 (
        .y(_T_553),
        .sel(_T_69),
        .a(1'h0),
        .b(_T_552)
    );
    wire _T_554;
    MUX_UNSIGNED #(.width(1)) u_mux_1644 (
        .y(_T_554),
        .sel(_T_65),
        .a(1'h0),
        .b(_T_553)
    );
    wire _T_555;
    MUX_UNSIGNED #(.width(1)) u_mux_1645 (
        .y(_T_555),
        .sel(_T_61),
        .a(1'h0),
        .b(_T_554)
    );
    wire _T_556;
    MUX_UNSIGNED #(.width(1)) u_mux_1646 (
        .y(_T_556),
        .sel(_T_57),
        .a(1'h0),
        .b(_T_555)
    );
    wire _T_557;
    MUX_UNSIGNED #(.width(1)) u_mux_1647 (
        .y(_T_557),
        .sel(_T_53),
        .a(1'h0),
        .b(_T_556)
    );
    wire _T_558;
    MUX_UNSIGNED #(.width(1)) u_mux_1648 (
        .y(_T_558),
        .sel(_T_49),
        .a(1'h0),
        .b(_T_557)
    );
    wire _T_559;
    MUX_UNSIGNED #(.width(1)) u_mux_1649 (
        .y(_T_559),
        .sel(_T_45),
        .a(1'h1),
        .b(_T_558)
    );
    wire _T_560;
    MUX_UNSIGNED #(.width(1)) u_mux_1650 (
        .y(_T_560),
        .sel(_T_41),
        .a(1'h1),
        .b(_T_559)
    );
    wire _T_561;
    MUX_UNSIGNED #(.width(1)) u_mux_1651 (
        .y(_T_561),
        .sel(_T_37),
        .a(1'h0),
        .b(_T_560)
    );
    wire ctrlSignals_6;
    MUX_UNSIGNED #(.width(1)) u_mux_1652 (
        .y(ctrlSignals_6),
        .sel(_T_33),
        .a(1'h0),
        .b(_T_561)
    );
    wire [1:0] _T_562;
    assign _T_562 = 2'h0;
    wire [1:0] _T_563;
    assign _T_563 = 2'h0;
    wire [1:0] _T_564;
    assign _T_564 = 2'h0;
    wire [1:0] _T_565;
    assign _T_565 = 2'h0;
    wire [1:0] _T_566;
    assign _T_566 = 2'h0;
    wire [1:0] _T_567;
    assign _T_567 = 2'h0;
    wire [1:0] _T_568;
    assign _T_568 = 2'h0;
    wire [1:0] _T_569;
    assign _T_569 = 2'h0;
    wire [1:0] _T_570;
    assign _T_570 = 2'h0;
    wire [1:0] _T_571;
    assign _T_571 = 2'h0;
    wire [1:0] _T_572;
    assign _T_572 = 2'h0;
    wire [1:0] _T_573;
    assign _T_573 = 2'h0;
    wire [1:0] _T_574;
    assign _T_574 = 2'h0;
    wire [1:0] _T_575;
    assign _T_575 = 2'h0;
    wire [1:0] _T_576;
    assign _T_576 = 2'h0;
    wire [1:0] _T_577;
    assign _T_577 = 2'h0;
    wire [1:0] _T_578;
    assign _T_578 = 2'h0;
    wire [1:0] _T_579;
    assign _T_579 = 2'h0;
    wire [1:0] _T_580;
    assign _T_580 = 2'h0;
    wire [1:0] _T_581;
    assign _T_581 = 2'h0;
    wire [1:0] _T_582;
    assign _T_582 = 2'h0;
    wire [1:0] _T_583;
    assign _T_583 = 2'h0;
    wire [1:0] _T_584;
    assign _T_584 = 2'h0;
    wire [1:0] _T_585;
    assign _T_585 = 2'h0;
    wire [1:0] _T_586;
    assign _T_586 = 2'h0;
    wire [1:0] _T_587;
    assign _T_587 = 2'h0;
    wire [1:0] _T_588;
    assign _T_588 = 2'h0;
    wire [1:0] _T_589;
    assign _T_589 = 2'h0;
    wire [1:0] _T_590;
    assign _T_590 = 2'h0;
    wire [1:0] _T_591;
    assign _T_591 = 2'h0;
    wire [1:0] _T_592;
    assign _T_592 = 2'h0;
    wire [1:0] _T_593;
    MUX_UNSIGNED #(.width(2)) u_mux_1653 (
        .y(_T_593),
        .sel(_T_101),
        .a(2'h1),
        .b(_T_592)
    );
    wire [1:0] _T_594;
    MUX_UNSIGNED #(.width(2)) u_mux_1654 (
        .y(_T_594),
        .sel(_T_97),
        .a(2'h2),
        .b(_T_593)
    );
    wire [1:0] _T_595;
    MUX_UNSIGNED #(.width(2)) u_mux_1655 (
        .y(_T_595),
        .sel(_T_93),
        .a(2'h3),
        .b(_T_594)
    );
    wire [1:0] _T_596;
    MUX_UNSIGNED #(.width(2)) u_mux_1656 (
        .y(_T_596),
        .sel(_T_89),
        .a(2'h0),
        .b(_T_595)
    );
    wire [1:0] _T_597;
    MUX_UNSIGNED #(.width(2)) u_mux_1657 (
        .y(_T_597),
        .sel(_T_85),
        .a(2'h0),
        .b(_T_596)
    );
    wire [1:0] _T_598;
    MUX_UNSIGNED #(.width(2)) u_mux_1658 (
        .y(_T_598),
        .sel(_T_81),
        .a(2'h0),
        .b(_T_597)
    );
    wire [1:0] _T_599;
    MUX_UNSIGNED #(.width(2)) u_mux_1659 (
        .y(_T_599),
        .sel(_T_77),
        .a(2'h0),
        .b(_T_598)
    );
    wire [1:0] _T_600;
    MUX_UNSIGNED #(.width(2)) u_mux_1660 (
        .y(_T_600),
        .sel(_T_73),
        .a(2'h0),
        .b(_T_599)
    );
    wire [1:0] _T_601;
    MUX_UNSIGNED #(.width(2)) u_mux_1661 (
        .y(_T_601),
        .sel(_T_69),
        .a(2'h0),
        .b(_T_600)
    );
    wire [1:0] _T_602;
    MUX_UNSIGNED #(.width(2)) u_mux_1662 (
        .y(_T_602),
        .sel(_T_65),
        .a(2'h0),
        .b(_T_601)
    );
    wire [1:0] _T_603;
    MUX_UNSIGNED #(.width(2)) u_mux_1663 (
        .y(_T_603),
        .sel(_T_61),
        .a(2'h0),
        .b(_T_602)
    );
    wire [1:0] _T_604;
    MUX_UNSIGNED #(.width(2)) u_mux_1664 (
        .y(_T_604),
        .sel(_T_57),
        .a(2'h0),
        .b(_T_603)
    );
    wire [1:0] _T_605;
    MUX_UNSIGNED #(.width(2)) u_mux_1665 (
        .y(_T_605),
        .sel(_T_53),
        .a(2'h0),
        .b(_T_604)
    );
    wire [1:0] _T_606;
    MUX_UNSIGNED #(.width(2)) u_mux_1666 (
        .y(_T_606),
        .sel(_T_49),
        .a(2'h0),
        .b(_T_605)
    );
    wire [1:0] _T_607;
    MUX_UNSIGNED #(.width(2)) u_mux_1667 (
        .y(_T_607),
        .sel(_T_45),
        .a(2'h0),
        .b(_T_606)
    );
    wire [1:0] _T_608;
    MUX_UNSIGNED #(.width(2)) u_mux_1668 (
        .y(_T_608),
        .sel(_T_41),
        .a(2'h0),
        .b(_T_607)
    );
    wire [1:0] _T_609;
    MUX_UNSIGNED #(.width(2)) u_mux_1669 (
        .y(_T_609),
        .sel(_T_37),
        .a(2'h0),
        .b(_T_608)
    );
    wire [1:0] ctrlSignals_7;
    MUX_UNSIGNED #(.width(2)) u_mux_1670 (
        .y(ctrlSignals_7),
        .sel(_T_33),
        .a(2'h0),
        .b(_T_609)
    );
    wire [2:0] _T_610;
    assign _T_610 = 3'h0;
    wire [2:0] _T_611;
    assign _T_611 = 3'h0;
    wire [2:0] _T_612;
    assign _T_612 = 3'h0;
    wire [2:0] _T_613;
    assign _T_613 = 3'h0;
    wire [2:0] _T_614;
    assign _T_614 = 3'h0;
    wire [2:0] _T_615;
    assign _T_615 = 3'h0;
    wire [2:0] _T_616;
    assign _T_616 = 3'h0;
    wire [2:0] _T_617;
    assign _T_617 = 3'h0;
    wire [2:0] _T_618;
    assign _T_618 = 3'h0;
    wire [2:0] _T_619;
    assign _T_619 = 3'h0;
    wire [2:0] _T_620;
    assign _T_620 = 3'h0;
    wire [2:0] _T_621;
    assign _T_621 = 3'h0;
    wire [2:0] _T_622;
    assign _T_622 = 3'h0;
    wire [2:0] _T_623;
    assign _T_623 = 3'h0;
    wire [2:0] _T_624;
    assign _T_624 = 3'h0;
    wire [2:0] _T_625;
    assign _T_625 = 3'h0;
    wire [2:0] _T_626;
    assign _T_626 = 3'h0;
    wire [2:0] _T_627;
    assign _T_627 = 3'h0;
    wire [2:0] _T_628;
    assign _T_628 = 3'h0;
    wire [2:0] _T_629;
    assign _T_629 = 3'h0;
    wire [2:0] _T_630;
    assign _T_630 = 3'h0;
    wire [2:0] _T_631;
    assign _T_631 = 3'h0;
    wire [2:0] _T_632;
    assign _T_632 = 3'h0;
    wire [2:0] _T_633;
    assign _T_633 = 3'h0;
    wire [2:0] _T_634;
    assign _T_634 = 3'h0;
    wire [2:0] _T_635;
    assign _T_635 = 3'h0;
    wire [2:0] _T_636;
    assign _T_636 = 3'h0;
    wire [2:0] _T_637;
    assign _T_637 = 3'h0;
    wire [2:0] _T_638;
    assign _T_638 = 3'h0;
    wire [2:0] _T_639;
    assign _T_639 = 3'h0;
    wire [2:0] _T_640;
    assign _T_640 = 3'h0;
    wire [2:0] _T_641;
    assign _T_641 = 3'h0;
    wire [2:0] _T_642;
    assign _T_642 = 3'h0;
    wire [2:0] _T_643;
    assign _T_643 = 3'h0;
    wire [2:0] _T_644;
    MUX_UNSIGNED #(.width(3)) u_mux_1671 (
        .y(_T_644),
        .sel(_T_89),
        .a(3'h4),
        .b(_T_643)
    );
    wire [2:0] _T_645;
    MUX_UNSIGNED #(.width(3)) u_mux_1672 (
        .y(_T_645),
        .sel(_T_85),
        .a(3'h5),
        .b(_T_644)
    );
    wire [2:0] _T_646;
    MUX_UNSIGNED #(.width(3)) u_mux_1673 (
        .y(_T_646),
        .sel(_T_81),
        .a(3'h1),
        .b(_T_645)
    );
    wire [2:0] _T_647;
    MUX_UNSIGNED #(.width(3)) u_mux_1674 (
        .y(_T_647),
        .sel(_T_77),
        .a(3'h2),
        .b(_T_646)
    );
    wire [2:0] _T_648;
    MUX_UNSIGNED #(.width(3)) u_mux_1675 (
        .y(_T_648),
        .sel(_T_73),
        .a(3'h3),
        .b(_T_647)
    );
    wire [2:0] _T_649;
    MUX_UNSIGNED #(.width(3)) u_mux_1676 (
        .y(_T_649),
        .sel(_T_69),
        .a(3'h0),
        .b(_T_648)
    );
    wire [2:0] _T_650;
    MUX_UNSIGNED #(.width(3)) u_mux_1677 (
        .y(_T_650),
        .sel(_T_65),
        .a(3'h0),
        .b(_T_649)
    );
    wire [2:0] _T_651;
    MUX_UNSIGNED #(.width(3)) u_mux_1678 (
        .y(_T_651),
        .sel(_T_61),
        .a(3'h0),
        .b(_T_650)
    );
    wire [2:0] _T_652;
    MUX_UNSIGNED #(.width(3)) u_mux_1679 (
        .y(_T_652),
        .sel(_T_57),
        .a(3'h0),
        .b(_T_651)
    );
    wire [2:0] _T_653;
    MUX_UNSIGNED #(.width(3)) u_mux_1680 (
        .y(_T_653),
        .sel(_T_53),
        .a(3'h0),
        .b(_T_652)
    );
    wire [2:0] _T_654;
    MUX_UNSIGNED #(.width(3)) u_mux_1681 (
        .y(_T_654),
        .sel(_T_49),
        .a(3'h0),
        .b(_T_653)
    );
    wire [2:0] _T_655;
    MUX_UNSIGNED #(.width(3)) u_mux_1682 (
        .y(_T_655),
        .sel(_T_45),
        .a(3'h0),
        .b(_T_654)
    );
    wire [2:0] _T_656;
    MUX_UNSIGNED #(.width(3)) u_mux_1683 (
        .y(_T_656),
        .sel(_T_41),
        .a(3'h0),
        .b(_T_655)
    );
    wire [2:0] _T_657;
    MUX_UNSIGNED #(.width(3)) u_mux_1684 (
        .y(_T_657),
        .sel(_T_37),
        .a(3'h0),
        .b(_T_656)
    );
    wire [2:0] ctrlSignals_8;
    MUX_UNSIGNED #(.width(3)) u_mux_1685 (
        .y(ctrlSignals_8),
        .sel(_T_33),
        .a(3'h0),
        .b(_T_657)
    );
    wire [1:0] _T_658;
    assign _T_658 = 2'h0;
    wire [1:0] _T_659;
    MUX_UNSIGNED #(.width(2)) u_mux_1686 (
        .y(_T_659),
        .sel(_T_221),
        .a(2'h3),
        .b(_T_658)
    );
    wire [1:0] _T_660;
    MUX_UNSIGNED #(.width(2)) u_mux_1687 (
        .y(_T_660),
        .sel(_T_217),
        .a(2'h3),
        .b(_T_659)
    );
    wire [1:0] _T_661;
    MUX_UNSIGNED #(.width(2)) u_mux_1688 (
        .y(_T_661),
        .sel(_T_213),
        .a(2'h3),
        .b(_T_660)
    );
    wire [1:0] _T_662;
    MUX_UNSIGNED #(.width(2)) u_mux_1689 (
        .y(_T_662),
        .sel(_T_209),
        .a(2'h3),
        .b(_T_661)
    );
    wire [1:0] _T_663;
    MUX_UNSIGNED #(.width(2)) u_mux_1690 (
        .y(_T_663),
        .sel(_T_205),
        .a(2'h3),
        .b(_T_662)
    );
    wire [1:0] _T_664;
    MUX_UNSIGNED #(.width(2)) u_mux_1691 (
        .y(_T_664),
        .sel(_T_201),
        .a(2'h3),
        .b(_T_663)
    );
    wire [1:0] _T_665;
    MUX_UNSIGNED #(.width(2)) u_mux_1692 (
        .y(_T_665),
        .sel(_T_197),
        .a(2'h3),
        .b(_T_664)
    );
    wire [1:0] _T_666;
    MUX_UNSIGNED #(.width(2)) u_mux_1693 (
        .y(_T_666),
        .sel(_T_193),
        .a(2'h3),
        .b(_T_665)
    );
    wire [1:0] _T_667;
    MUX_UNSIGNED #(.width(2)) u_mux_1694 (
        .y(_T_667),
        .sel(_T_189),
        .a(2'h3),
        .b(_T_666)
    );
    wire [1:0] _T_668;
    MUX_UNSIGNED #(.width(2)) u_mux_1695 (
        .y(_T_668),
        .sel(_T_185),
        .a(2'h0),
        .b(_T_667)
    );
    wire [1:0] _T_669;
    MUX_UNSIGNED #(.width(2)) u_mux_1696 (
        .y(_T_669),
        .sel(_T_181),
        .a(2'h0),
        .b(_T_668)
    );
    wire [1:0] _T_670;
    MUX_UNSIGNED #(.width(2)) u_mux_1697 (
        .y(_T_670),
        .sel(_T_177),
        .a(2'h0),
        .b(_T_669)
    );
    wire [1:0] _T_671;
    MUX_UNSIGNED #(.width(2)) u_mux_1698 (
        .y(_T_671),
        .sel(_T_173),
        .a(2'h0),
        .b(_T_670)
    );
    wire [1:0] _T_672;
    MUX_UNSIGNED #(.width(2)) u_mux_1699 (
        .y(_T_672),
        .sel(_T_169),
        .a(2'h0),
        .b(_T_671)
    );
    wire [1:0] _T_673;
    MUX_UNSIGNED #(.width(2)) u_mux_1700 (
        .y(_T_673),
        .sel(_T_165),
        .a(2'h0),
        .b(_T_672)
    );
    wire [1:0] _T_674;
    MUX_UNSIGNED #(.width(2)) u_mux_1701 (
        .y(_T_674),
        .sel(_T_161),
        .a(2'h0),
        .b(_T_673)
    );
    wire [1:0] _T_675;
    MUX_UNSIGNED #(.width(2)) u_mux_1702 (
        .y(_T_675),
        .sel(_T_157),
        .a(2'h0),
        .b(_T_674)
    );
    wire [1:0] _T_676;
    MUX_UNSIGNED #(.width(2)) u_mux_1703 (
        .y(_T_676),
        .sel(_T_153),
        .a(2'h0),
        .b(_T_675)
    );
    wire [1:0] _T_677;
    MUX_UNSIGNED #(.width(2)) u_mux_1704 (
        .y(_T_677),
        .sel(_T_149),
        .a(2'h0),
        .b(_T_676)
    );
    wire [1:0] _T_678;
    MUX_UNSIGNED #(.width(2)) u_mux_1705 (
        .y(_T_678),
        .sel(_T_145),
        .a(2'h0),
        .b(_T_677)
    );
    wire [1:0] _T_679;
    MUX_UNSIGNED #(.width(2)) u_mux_1706 (
        .y(_T_679),
        .sel(_T_141),
        .a(2'h0),
        .b(_T_678)
    );
    wire [1:0] _T_680;
    MUX_UNSIGNED #(.width(2)) u_mux_1707 (
        .y(_T_680),
        .sel(_T_137),
        .a(2'h0),
        .b(_T_679)
    );
    wire [1:0] _T_681;
    MUX_UNSIGNED #(.width(2)) u_mux_1708 (
        .y(_T_681),
        .sel(_T_133),
        .a(2'h0),
        .b(_T_680)
    );
    wire [1:0] _T_682;
    MUX_UNSIGNED #(.width(2)) u_mux_1709 (
        .y(_T_682),
        .sel(_T_129),
        .a(2'h0),
        .b(_T_681)
    );
    wire [1:0] _T_683;
    MUX_UNSIGNED #(.width(2)) u_mux_1710 (
        .y(_T_683),
        .sel(_T_125),
        .a(2'h0),
        .b(_T_682)
    );
    wire [1:0] _T_684;
    MUX_UNSIGNED #(.width(2)) u_mux_1711 (
        .y(_T_684),
        .sel(_T_121),
        .a(2'h0),
        .b(_T_683)
    );
    wire [1:0] _T_685;
    MUX_UNSIGNED #(.width(2)) u_mux_1712 (
        .y(_T_685),
        .sel(_T_117),
        .a(2'h0),
        .b(_T_684)
    );
    wire [1:0] _T_686;
    MUX_UNSIGNED #(.width(2)) u_mux_1713 (
        .y(_T_686),
        .sel(_T_113),
        .a(2'h0),
        .b(_T_685)
    );
    wire [1:0] _T_687;
    MUX_UNSIGNED #(.width(2)) u_mux_1714 (
        .y(_T_687),
        .sel(_T_109),
        .a(2'h0),
        .b(_T_686)
    );
    wire [1:0] _T_688;
    MUX_UNSIGNED #(.width(2)) u_mux_1715 (
        .y(_T_688),
        .sel(_T_105),
        .a(2'h0),
        .b(_T_687)
    );
    wire [1:0] _T_689;
    MUX_UNSIGNED #(.width(2)) u_mux_1716 (
        .y(_T_689),
        .sel(_T_101),
        .a(2'h0),
        .b(_T_688)
    );
    wire [1:0] _T_690;
    MUX_UNSIGNED #(.width(2)) u_mux_1717 (
        .y(_T_690),
        .sel(_T_97),
        .a(2'h0),
        .b(_T_689)
    );
    wire [1:0] _T_691;
    MUX_UNSIGNED #(.width(2)) u_mux_1718 (
        .y(_T_691),
        .sel(_T_93),
        .a(2'h0),
        .b(_T_690)
    );
    wire [1:0] _T_692;
    MUX_UNSIGNED #(.width(2)) u_mux_1719 (
        .y(_T_692),
        .sel(_T_89),
        .a(2'h1),
        .b(_T_691)
    );
    wire [1:0] _T_693;
    MUX_UNSIGNED #(.width(2)) u_mux_1720 (
        .y(_T_693),
        .sel(_T_85),
        .a(2'h1),
        .b(_T_692)
    );
    wire [1:0] _T_694;
    MUX_UNSIGNED #(.width(2)) u_mux_1721 (
        .y(_T_694),
        .sel(_T_81),
        .a(2'h1),
        .b(_T_693)
    );
    wire [1:0] _T_695;
    MUX_UNSIGNED #(.width(2)) u_mux_1722 (
        .y(_T_695),
        .sel(_T_77),
        .a(2'h1),
        .b(_T_694)
    );
    wire [1:0] _T_696;
    MUX_UNSIGNED #(.width(2)) u_mux_1723 (
        .y(_T_696),
        .sel(_T_73),
        .a(2'h1),
        .b(_T_695)
    );
    wire [1:0] _T_697;
    MUX_UNSIGNED #(.width(2)) u_mux_1724 (
        .y(_T_697),
        .sel(_T_69),
        .a(2'h0),
        .b(_T_696)
    );
    wire [1:0] _T_698;
    MUX_UNSIGNED #(.width(2)) u_mux_1725 (
        .y(_T_698),
        .sel(_T_65),
        .a(2'h0),
        .b(_T_697)
    );
    wire [1:0] _T_699;
    MUX_UNSIGNED #(.width(2)) u_mux_1726 (
        .y(_T_699),
        .sel(_T_61),
        .a(2'h0),
        .b(_T_698)
    );
    wire [1:0] _T_700;
    MUX_UNSIGNED #(.width(2)) u_mux_1727 (
        .y(_T_700),
        .sel(_T_57),
        .a(2'h0),
        .b(_T_699)
    );
    wire [1:0] _T_701;
    MUX_UNSIGNED #(.width(2)) u_mux_1728 (
        .y(_T_701),
        .sel(_T_53),
        .a(2'h0),
        .b(_T_700)
    );
    wire [1:0] _T_702;
    MUX_UNSIGNED #(.width(2)) u_mux_1729 (
        .y(_T_702),
        .sel(_T_49),
        .a(2'h0),
        .b(_T_701)
    );
    wire [1:0] _T_703;
    MUX_UNSIGNED #(.width(2)) u_mux_1730 (
        .y(_T_703),
        .sel(_T_45),
        .a(2'h2),
        .b(_T_702)
    );
    wire [1:0] _T_704;
    MUX_UNSIGNED #(.width(2)) u_mux_1731 (
        .y(_T_704),
        .sel(_T_41),
        .a(2'h2),
        .b(_T_703)
    );
    wire [1:0] _T_705;
    MUX_UNSIGNED #(.width(2)) u_mux_1732 (
        .y(_T_705),
        .sel(_T_37),
        .a(2'h0),
        .b(_T_704)
    );
    wire [1:0] ctrlSignals_9;
    MUX_UNSIGNED #(.width(2)) u_mux_1733 (
        .y(ctrlSignals_9),
        .sel(_T_33),
        .a(2'h0),
        .b(_T_705)
    );
    wire _T_706;
    assign _T_706 = 1'h0;
    wire _T_707;
    assign _T_707 = 1'h0;
    wire _T_708;
    assign _T_708 = 1'h0;
    wire _T_709;
    assign _T_709 = 1'h0;
    wire _T_710;
    MUX_UNSIGNED #(.width(1)) u_mux_1734 (
        .y(_T_710),
        .sel(_T_209),
        .a(1'h1),
        .b(_T_709)
    );
    wire _T_711;
    MUX_UNSIGNED #(.width(1)) u_mux_1735 (
        .y(_T_711),
        .sel(_T_205),
        .a(1'h1),
        .b(_T_710)
    );
    wire _T_712;
    MUX_UNSIGNED #(.width(1)) u_mux_1736 (
        .y(_T_712),
        .sel(_T_201),
        .a(1'h1),
        .b(_T_711)
    );
    wire _T_713;
    MUX_UNSIGNED #(.width(1)) u_mux_1737 (
        .y(_T_713),
        .sel(_T_197),
        .a(1'h1),
        .b(_T_712)
    );
    wire _T_714;
    MUX_UNSIGNED #(.width(1)) u_mux_1738 (
        .y(_T_714),
        .sel(_T_193),
        .a(1'h1),
        .b(_T_713)
    );
    wire _T_715;
    MUX_UNSIGNED #(.width(1)) u_mux_1739 (
        .y(_T_715),
        .sel(_T_189),
        .a(1'h1),
        .b(_T_714)
    );
    wire _T_716;
    MUX_UNSIGNED #(.width(1)) u_mux_1740 (
        .y(_T_716),
        .sel(_T_185),
        .a(1'h0),
        .b(_T_715)
    );
    wire _T_717;
    MUX_UNSIGNED #(.width(1)) u_mux_1741 (
        .y(_T_717),
        .sel(_T_181),
        .a(1'h0),
        .b(_T_716)
    );
    wire _T_718;
    MUX_UNSIGNED #(.width(1)) u_mux_1742 (
        .y(_T_718),
        .sel(_T_177),
        .a(1'h1),
        .b(_T_717)
    );
    wire _T_719;
    MUX_UNSIGNED #(.width(1)) u_mux_1743 (
        .y(_T_719),
        .sel(_T_173),
        .a(1'h1),
        .b(_T_718)
    );
    wire _T_720;
    MUX_UNSIGNED #(.width(1)) u_mux_1744 (
        .y(_T_720),
        .sel(_T_169),
        .a(1'h1),
        .b(_T_719)
    );
    wire _T_721;
    MUX_UNSIGNED #(.width(1)) u_mux_1745 (
        .y(_T_721),
        .sel(_T_165),
        .a(1'h1),
        .b(_T_720)
    );
    wire _T_722;
    MUX_UNSIGNED #(.width(1)) u_mux_1746 (
        .y(_T_722),
        .sel(_T_161),
        .a(1'h1),
        .b(_T_721)
    );
    wire _T_723;
    MUX_UNSIGNED #(.width(1)) u_mux_1747 (
        .y(_T_723),
        .sel(_T_157),
        .a(1'h1),
        .b(_T_722)
    );
    wire _T_724;
    MUX_UNSIGNED #(.width(1)) u_mux_1748 (
        .y(_T_724),
        .sel(_T_153),
        .a(1'h1),
        .b(_T_723)
    );
    wire _T_725;
    MUX_UNSIGNED #(.width(1)) u_mux_1749 (
        .y(_T_725),
        .sel(_T_149),
        .a(1'h1),
        .b(_T_724)
    );
    wire _T_726;
    MUX_UNSIGNED #(.width(1)) u_mux_1750 (
        .y(_T_726),
        .sel(_T_145),
        .a(1'h1),
        .b(_T_725)
    );
    wire _T_727;
    MUX_UNSIGNED #(.width(1)) u_mux_1751 (
        .y(_T_727),
        .sel(_T_141),
        .a(1'h1),
        .b(_T_726)
    );
    wire _T_728;
    MUX_UNSIGNED #(.width(1)) u_mux_1752 (
        .y(_T_728),
        .sel(_T_137),
        .a(1'h1),
        .b(_T_727)
    );
    wire _T_729;
    MUX_UNSIGNED #(.width(1)) u_mux_1753 (
        .y(_T_729),
        .sel(_T_133),
        .a(1'h1),
        .b(_T_728)
    );
    wire _T_730;
    MUX_UNSIGNED #(.width(1)) u_mux_1754 (
        .y(_T_730),
        .sel(_T_129),
        .a(1'h1),
        .b(_T_729)
    );
    wire _T_731;
    MUX_UNSIGNED #(.width(1)) u_mux_1755 (
        .y(_T_731),
        .sel(_T_125),
        .a(1'h1),
        .b(_T_730)
    );
    wire _T_732;
    MUX_UNSIGNED #(.width(1)) u_mux_1756 (
        .y(_T_732),
        .sel(_T_121),
        .a(1'h1),
        .b(_T_731)
    );
    wire _T_733;
    MUX_UNSIGNED #(.width(1)) u_mux_1757 (
        .y(_T_733),
        .sel(_T_117),
        .a(1'h1),
        .b(_T_732)
    );
    wire _T_734;
    MUX_UNSIGNED #(.width(1)) u_mux_1758 (
        .y(_T_734),
        .sel(_T_113),
        .a(1'h1),
        .b(_T_733)
    );
    wire _T_735;
    MUX_UNSIGNED #(.width(1)) u_mux_1759 (
        .y(_T_735),
        .sel(_T_109),
        .a(1'h1),
        .b(_T_734)
    );
    wire _T_736;
    MUX_UNSIGNED #(.width(1)) u_mux_1760 (
        .y(_T_736),
        .sel(_T_105),
        .a(1'h1),
        .b(_T_735)
    );
    wire _T_737;
    MUX_UNSIGNED #(.width(1)) u_mux_1761 (
        .y(_T_737),
        .sel(_T_101),
        .a(1'h0),
        .b(_T_736)
    );
    wire _T_738;
    MUX_UNSIGNED #(.width(1)) u_mux_1762 (
        .y(_T_738),
        .sel(_T_97),
        .a(1'h0),
        .b(_T_737)
    );
    wire _T_739;
    MUX_UNSIGNED #(.width(1)) u_mux_1763 (
        .y(_T_739),
        .sel(_T_93),
        .a(1'h0),
        .b(_T_738)
    );
    wire _T_740;
    MUX_UNSIGNED #(.width(1)) u_mux_1764 (
        .y(_T_740),
        .sel(_T_89),
        .a(1'h1),
        .b(_T_739)
    );
    wire _T_741;
    MUX_UNSIGNED #(.width(1)) u_mux_1765 (
        .y(_T_741),
        .sel(_T_85),
        .a(1'h1),
        .b(_T_740)
    );
    wire _T_742;
    MUX_UNSIGNED #(.width(1)) u_mux_1766 (
        .y(_T_742),
        .sel(_T_81),
        .a(1'h1),
        .b(_T_741)
    );
    wire _T_743;
    MUX_UNSIGNED #(.width(1)) u_mux_1767 (
        .y(_T_743),
        .sel(_T_77),
        .a(1'h1),
        .b(_T_742)
    );
    wire _T_744;
    MUX_UNSIGNED #(.width(1)) u_mux_1768 (
        .y(_T_744),
        .sel(_T_73),
        .a(1'h1),
        .b(_T_743)
    );
    wire _T_745;
    MUX_UNSIGNED #(.width(1)) u_mux_1769 (
        .y(_T_745),
        .sel(_T_69),
        .a(1'h0),
        .b(_T_744)
    );
    wire _T_746;
    MUX_UNSIGNED #(.width(1)) u_mux_1770 (
        .y(_T_746),
        .sel(_T_65),
        .a(1'h0),
        .b(_T_745)
    );
    wire _T_747;
    MUX_UNSIGNED #(.width(1)) u_mux_1771 (
        .y(_T_747),
        .sel(_T_61),
        .a(1'h0),
        .b(_T_746)
    );
    wire _T_748;
    MUX_UNSIGNED #(.width(1)) u_mux_1772 (
        .y(_T_748),
        .sel(_T_57),
        .a(1'h0),
        .b(_T_747)
    );
    wire _T_749;
    MUX_UNSIGNED #(.width(1)) u_mux_1773 (
        .y(_T_749),
        .sel(_T_53),
        .a(1'h0),
        .b(_T_748)
    );
    wire _T_750;
    MUX_UNSIGNED #(.width(1)) u_mux_1774 (
        .y(_T_750),
        .sel(_T_49),
        .a(1'h0),
        .b(_T_749)
    );
    wire _T_751;
    MUX_UNSIGNED #(.width(1)) u_mux_1775 (
        .y(_T_751),
        .sel(_T_45),
        .a(1'h1),
        .b(_T_750)
    );
    wire _T_752;
    MUX_UNSIGNED #(.width(1)) u_mux_1776 (
        .y(_T_752),
        .sel(_T_41),
        .a(1'h1),
        .b(_T_751)
    );
    wire _T_753;
    MUX_UNSIGNED #(.width(1)) u_mux_1777 (
        .y(_T_753),
        .sel(_T_37),
        .a(1'h1),
        .b(_T_752)
    );
    wire ctrlSignals_10;
    MUX_UNSIGNED #(.width(1)) u_mux_1778 (
        .y(ctrlSignals_10),
        .sel(_T_33),
        .a(1'h1),
        .b(_T_753)
    );
    wire [2:0] _T_754;
    assign _T_754 = 3'h0;
    wire [2:0] _T_755;
    MUX_UNSIGNED #(.width(3)) u_mux_1779 (
        .y(_T_755),
        .sel(_T_221),
        .a(3'h4),
        .b(_T_754)
    );
    wire [2:0] _T_756;
    MUX_UNSIGNED #(.width(3)) u_mux_1780 (
        .y(_T_756),
        .sel(_T_217),
        .a(3'h4),
        .b(_T_755)
    );
    wire [2:0] _T_757;
    MUX_UNSIGNED #(.width(3)) u_mux_1781 (
        .y(_T_757),
        .sel(_T_213),
        .a(3'h4),
        .b(_T_756)
    );
    wire [2:0] _T_758;
    MUX_UNSIGNED #(.width(3)) u_mux_1782 (
        .y(_T_758),
        .sel(_T_209),
        .a(3'h3),
        .b(_T_757)
    );
    wire [2:0] _T_759;
    MUX_UNSIGNED #(.width(3)) u_mux_1783 (
        .y(_T_759),
        .sel(_T_205),
        .a(3'h2),
        .b(_T_758)
    );
    wire [2:0] _T_760;
    MUX_UNSIGNED #(.width(3)) u_mux_1784 (
        .y(_T_760),
        .sel(_T_201),
        .a(3'h1),
        .b(_T_759)
    );
    wire [2:0] _T_761;
    MUX_UNSIGNED #(.width(3)) u_mux_1785 (
        .y(_T_761),
        .sel(_T_197),
        .a(3'h3),
        .b(_T_760)
    );
    wire [2:0] _T_762;
    MUX_UNSIGNED #(.width(3)) u_mux_1786 (
        .y(_T_762),
        .sel(_T_193),
        .a(3'h2),
        .b(_T_761)
    );
    wire [2:0] _T_763;
    MUX_UNSIGNED #(.width(3)) u_mux_1787 (
        .y(_T_763),
        .sel(_T_189),
        .a(3'h1),
        .b(_T_762)
    );
    wire [2:0] _T_764;
    MUX_UNSIGNED #(.width(3)) u_mux_1788 (
        .y(_T_764),
        .sel(_T_185),
        .a(3'h0),
        .b(_T_763)
    );
    wire [2:0] _T_765;
    MUX_UNSIGNED #(.width(3)) u_mux_1789 (
        .y(_T_765),
        .sel(_T_181),
        .a(3'h0),
        .b(_T_764)
    );
    wire [2:0] _T_766;
    MUX_UNSIGNED #(.width(3)) u_mux_1790 (
        .y(_T_766),
        .sel(_T_177),
        .a(3'h0),
        .b(_T_765)
    );
    wire [2:0] _T_767;
    MUX_UNSIGNED #(.width(3)) u_mux_1791 (
        .y(_T_767),
        .sel(_T_173),
        .a(3'h0),
        .b(_T_766)
    );
    wire [2:0] _T_768;
    MUX_UNSIGNED #(.width(3)) u_mux_1792 (
        .y(_T_768),
        .sel(_T_169),
        .a(3'h0),
        .b(_T_767)
    );
    wire [2:0] _T_769;
    MUX_UNSIGNED #(.width(3)) u_mux_1793 (
        .y(_T_769),
        .sel(_T_165),
        .a(3'h0),
        .b(_T_768)
    );
    wire [2:0] _T_770;
    MUX_UNSIGNED #(.width(3)) u_mux_1794 (
        .y(_T_770),
        .sel(_T_161),
        .a(3'h0),
        .b(_T_769)
    );
    wire [2:0] _T_771;
    MUX_UNSIGNED #(.width(3)) u_mux_1795 (
        .y(_T_771),
        .sel(_T_157),
        .a(3'h0),
        .b(_T_770)
    );
    wire [2:0] _T_772;
    MUX_UNSIGNED #(.width(3)) u_mux_1796 (
        .y(_T_772),
        .sel(_T_153),
        .a(3'h0),
        .b(_T_771)
    );
    wire [2:0] _T_773;
    MUX_UNSIGNED #(.width(3)) u_mux_1797 (
        .y(_T_773),
        .sel(_T_149),
        .a(3'h0),
        .b(_T_772)
    );
    wire [2:0] _T_774;
    MUX_UNSIGNED #(.width(3)) u_mux_1798 (
        .y(_T_774),
        .sel(_T_145),
        .a(3'h0),
        .b(_T_773)
    );
    wire [2:0] _T_775;
    MUX_UNSIGNED #(.width(3)) u_mux_1799 (
        .y(_T_775),
        .sel(_T_141),
        .a(3'h0),
        .b(_T_774)
    );
    wire [2:0] _T_776;
    MUX_UNSIGNED #(.width(3)) u_mux_1800 (
        .y(_T_776),
        .sel(_T_137),
        .a(3'h0),
        .b(_T_775)
    );
    wire [2:0] _T_777;
    MUX_UNSIGNED #(.width(3)) u_mux_1801 (
        .y(_T_777),
        .sel(_T_133),
        .a(3'h0),
        .b(_T_776)
    );
    wire [2:0] _T_778;
    MUX_UNSIGNED #(.width(3)) u_mux_1802 (
        .y(_T_778),
        .sel(_T_129),
        .a(3'h0),
        .b(_T_777)
    );
    wire [2:0] _T_779;
    MUX_UNSIGNED #(.width(3)) u_mux_1803 (
        .y(_T_779),
        .sel(_T_125),
        .a(3'h0),
        .b(_T_778)
    );
    wire [2:0] _T_780;
    MUX_UNSIGNED #(.width(3)) u_mux_1804 (
        .y(_T_780),
        .sel(_T_121),
        .a(3'h0),
        .b(_T_779)
    );
    wire [2:0] _T_781;
    MUX_UNSIGNED #(.width(3)) u_mux_1805 (
        .y(_T_781),
        .sel(_T_117),
        .a(3'h0),
        .b(_T_780)
    );
    wire [2:0] _T_782;
    MUX_UNSIGNED #(.width(3)) u_mux_1806 (
        .y(_T_782),
        .sel(_T_113),
        .a(3'h0),
        .b(_T_781)
    );
    wire [2:0] _T_783;
    MUX_UNSIGNED #(.width(3)) u_mux_1807 (
        .y(_T_783),
        .sel(_T_109),
        .a(3'h0),
        .b(_T_782)
    );
    wire [2:0] _T_784;
    MUX_UNSIGNED #(.width(3)) u_mux_1808 (
        .y(_T_784),
        .sel(_T_105),
        .a(3'h0),
        .b(_T_783)
    );
    wire [2:0] _T_785;
    MUX_UNSIGNED #(.width(3)) u_mux_1809 (
        .y(_T_785),
        .sel(_T_101),
        .a(3'h0),
        .b(_T_784)
    );
    wire [2:0] _T_786;
    MUX_UNSIGNED #(.width(3)) u_mux_1810 (
        .y(_T_786),
        .sel(_T_97),
        .a(3'h0),
        .b(_T_785)
    );
    wire [2:0] _T_787;
    MUX_UNSIGNED #(.width(3)) u_mux_1811 (
        .y(_T_787),
        .sel(_T_93),
        .a(3'h0),
        .b(_T_786)
    );
    wire [2:0] _T_788;
    MUX_UNSIGNED #(.width(3)) u_mux_1812 (
        .y(_T_788),
        .sel(_T_89),
        .a(3'h0),
        .b(_T_787)
    );
    wire [2:0] _T_789;
    MUX_UNSIGNED #(.width(3)) u_mux_1813 (
        .y(_T_789),
        .sel(_T_85),
        .a(3'h0),
        .b(_T_788)
    );
    wire [2:0] _T_790;
    MUX_UNSIGNED #(.width(3)) u_mux_1814 (
        .y(_T_790),
        .sel(_T_81),
        .a(3'h0),
        .b(_T_789)
    );
    wire [2:0] _T_791;
    MUX_UNSIGNED #(.width(3)) u_mux_1815 (
        .y(_T_791),
        .sel(_T_77),
        .a(3'h0),
        .b(_T_790)
    );
    wire [2:0] _T_792;
    MUX_UNSIGNED #(.width(3)) u_mux_1816 (
        .y(_T_792),
        .sel(_T_73),
        .a(3'h0),
        .b(_T_791)
    );
    wire [2:0] _T_793;
    MUX_UNSIGNED #(.width(3)) u_mux_1817 (
        .y(_T_793),
        .sel(_T_69),
        .a(3'h0),
        .b(_T_792)
    );
    wire [2:0] _T_794;
    MUX_UNSIGNED #(.width(3)) u_mux_1818 (
        .y(_T_794),
        .sel(_T_65),
        .a(3'h0),
        .b(_T_793)
    );
    wire [2:0] _T_795;
    MUX_UNSIGNED #(.width(3)) u_mux_1819 (
        .y(_T_795),
        .sel(_T_61),
        .a(3'h0),
        .b(_T_794)
    );
    wire [2:0] _T_796;
    MUX_UNSIGNED #(.width(3)) u_mux_1820 (
        .y(_T_796),
        .sel(_T_57),
        .a(3'h0),
        .b(_T_795)
    );
    wire [2:0] _T_797;
    MUX_UNSIGNED #(.width(3)) u_mux_1821 (
        .y(_T_797),
        .sel(_T_53),
        .a(3'h0),
        .b(_T_796)
    );
    wire [2:0] _T_798;
    MUX_UNSIGNED #(.width(3)) u_mux_1822 (
        .y(_T_798),
        .sel(_T_49),
        .a(3'h0),
        .b(_T_797)
    );
    wire [2:0] _T_799;
    MUX_UNSIGNED #(.width(3)) u_mux_1823 (
        .y(_T_799),
        .sel(_T_45),
        .a(3'h0),
        .b(_T_798)
    );
    wire [2:0] _T_800;
    MUX_UNSIGNED #(.width(3)) u_mux_1824 (
        .y(_T_800),
        .sel(_T_41),
        .a(3'h0),
        .b(_T_799)
    );
    wire [2:0] _T_801;
    MUX_UNSIGNED #(.width(3)) u_mux_1825 (
        .y(_T_801),
        .sel(_T_37),
        .a(3'h0),
        .b(_T_800)
    );
    wire [2:0] ctrlSignals_11;
    MUX_UNSIGNED #(.width(3)) u_mux_1826 (
        .y(ctrlSignals_11),
        .sel(_T_33),
        .a(3'h0),
        .b(_T_801)
    );
    wire _T_802;
    MUX_UNSIGNED #(.width(1)) u_mux_1827 (
        .y(_T_802),
        .sel(_T_225),
        .a(1'h0),
        .b(1'h1)
    );
    wire _T_803;
    MUX_UNSIGNED #(.width(1)) u_mux_1828 (
        .y(_T_803),
        .sel(_T_221),
        .a(1'h0),
        .b(_T_802)
    );
    wire _T_804;
    MUX_UNSIGNED #(.width(1)) u_mux_1829 (
        .y(_T_804),
        .sel(_T_217),
        .a(1'h0),
        .b(_T_803)
    );
    wire _T_805;
    MUX_UNSIGNED #(.width(1)) u_mux_1830 (
        .y(_T_805),
        .sel(_T_213),
        .a(1'h0),
        .b(_T_804)
    );
    wire _T_806;
    MUX_UNSIGNED #(.width(1)) u_mux_1831 (
        .y(_T_806),
        .sel(_T_209),
        .a(1'h0),
        .b(_T_805)
    );
    wire _T_807;
    MUX_UNSIGNED #(.width(1)) u_mux_1832 (
        .y(_T_807),
        .sel(_T_205),
        .a(1'h0),
        .b(_T_806)
    );
    wire _T_808;
    MUX_UNSIGNED #(.width(1)) u_mux_1833 (
        .y(_T_808),
        .sel(_T_201),
        .a(1'h0),
        .b(_T_807)
    );
    wire _T_809;
    MUX_UNSIGNED #(.width(1)) u_mux_1834 (
        .y(_T_809),
        .sel(_T_197),
        .a(1'h0),
        .b(_T_808)
    );
    wire _T_810;
    MUX_UNSIGNED #(.width(1)) u_mux_1835 (
        .y(_T_810),
        .sel(_T_193),
        .a(1'h0),
        .b(_T_809)
    );
    wire _T_811;
    MUX_UNSIGNED #(.width(1)) u_mux_1836 (
        .y(_T_811),
        .sel(_T_189),
        .a(1'h0),
        .b(_T_810)
    );
    wire _T_812;
    MUX_UNSIGNED #(.width(1)) u_mux_1837 (
        .y(_T_812),
        .sel(_T_185),
        .a(1'h0),
        .b(_T_811)
    );
    wire _T_813;
    MUX_UNSIGNED #(.width(1)) u_mux_1838 (
        .y(_T_813),
        .sel(_T_181),
        .a(1'h0),
        .b(_T_812)
    );
    wire _T_814;
    MUX_UNSIGNED #(.width(1)) u_mux_1839 (
        .y(_T_814),
        .sel(_T_177),
        .a(1'h0),
        .b(_T_813)
    );
    wire _T_815;
    MUX_UNSIGNED #(.width(1)) u_mux_1840 (
        .y(_T_815),
        .sel(_T_173),
        .a(1'h0),
        .b(_T_814)
    );
    wire _T_816;
    MUX_UNSIGNED #(.width(1)) u_mux_1841 (
        .y(_T_816),
        .sel(_T_169),
        .a(1'h0),
        .b(_T_815)
    );
    wire _T_817;
    MUX_UNSIGNED #(.width(1)) u_mux_1842 (
        .y(_T_817),
        .sel(_T_165),
        .a(1'h0),
        .b(_T_816)
    );
    wire _T_818;
    MUX_UNSIGNED #(.width(1)) u_mux_1843 (
        .y(_T_818),
        .sel(_T_161),
        .a(1'h0),
        .b(_T_817)
    );
    wire _T_819;
    MUX_UNSIGNED #(.width(1)) u_mux_1844 (
        .y(_T_819),
        .sel(_T_157),
        .a(1'h0),
        .b(_T_818)
    );
    wire _T_820;
    MUX_UNSIGNED #(.width(1)) u_mux_1845 (
        .y(_T_820),
        .sel(_T_153),
        .a(1'h0),
        .b(_T_819)
    );
    wire _T_821;
    MUX_UNSIGNED #(.width(1)) u_mux_1846 (
        .y(_T_821),
        .sel(_T_149),
        .a(1'h0),
        .b(_T_820)
    );
    wire _T_822;
    MUX_UNSIGNED #(.width(1)) u_mux_1847 (
        .y(_T_822),
        .sel(_T_145),
        .a(1'h0),
        .b(_T_821)
    );
    wire _T_823;
    MUX_UNSIGNED #(.width(1)) u_mux_1848 (
        .y(_T_823),
        .sel(_T_141),
        .a(1'h0),
        .b(_T_822)
    );
    wire _T_824;
    MUX_UNSIGNED #(.width(1)) u_mux_1849 (
        .y(_T_824),
        .sel(_T_137),
        .a(1'h0),
        .b(_T_823)
    );
    wire _T_825;
    MUX_UNSIGNED #(.width(1)) u_mux_1850 (
        .y(_T_825),
        .sel(_T_133),
        .a(1'h0),
        .b(_T_824)
    );
    wire _T_826;
    MUX_UNSIGNED #(.width(1)) u_mux_1851 (
        .y(_T_826),
        .sel(_T_129),
        .a(1'h0),
        .b(_T_825)
    );
    wire _T_827;
    MUX_UNSIGNED #(.width(1)) u_mux_1852 (
        .y(_T_827),
        .sel(_T_125),
        .a(1'h0),
        .b(_T_826)
    );
    wire _T_828;
    MUX_UNSIGNED #(.width(1)) u_mux_1853 (
        .y(_T_828),
        .sel(_T_121),
        .a(1'h0),
        .b(_T_827)
    );
    wire _T_829;
    MUX_UNSIGNED #(.width(1)) u_mux_1854 (
        .y(_T_829),
        .sel(_T_117),
        .a(1'h0),
        .b(_T_828)
    );
    wire _T_830;
    MUX_UNSIGNED #(.width(1)) u_mux_1855 (
        .y(_T_830),
        .sel(_T_113),
        .a(1'h0),
        .b(_T_829)
    );
    wire _T_831;
    MUX_UNSIGNED #(.width(1)) u_mux_1856 (
        .y(_T_831),
        .sel(_T_109),
        .a(1'h0),
        .b(_T_830)
    );
    wire _T_832;
    MUX_UNSIGNED #(.width(1)) u_mux_1857 (
        .y(_T_832),
        .sel(_T_105),
        .a(1'h0),
        .b(_T_831)
    );
    wire _T_833;
    MUX_UNSIGNED #(.width(1)) u_mux_1858 (
        .y(_T_833),
        .sel(_T_101),
        .a(1'h0),
        .b(_T_832)
    );
    wire _T_834;
    MUX_UNSIGNED #(.width(1)) u_mux_1859 (
        .y(_T_834),
        .sel(_T_97),
        .a(1'h0),
        .b(_T_833)
    );
    wire _T_835;
    MUX_UNSIGNED #(.width(1)) u_mux_1860 (
        .y(_T_835),
        .sel(_T_93),
        .a(1'h0),
        .b(_T_834)
    );
    wire _T_836;
    MUX_UNSIGNED #(.width(1)) u_mux_1861 (
        .y(_T_836),
        .sel(_T_89),
        .a(1'h0),
        .b(_T_835)
    );
    wire _T_837;
    MUX_UNSIGNED #(.width(1)) u_mux_1862 (
        .y(_T_837),
        .sel(_T_85),
        .a(1'h0),
        .b(_T_836)
    );
    wire _T_838;
    MUX_UNSIGNED #(.width(1)) u_mux_1863 (
        .y(_T_838),
        .sel(_T_81),
        .a(1'h0),
        .b(_T_837)
    );
    wire _T_839;
    MUX_UNSIGNED #(.width(1)) u_mux_1864 (
        .y(_T_839),
        .sel(_T_77),
        .a(1'h0),
        .b(_T_838)
    );
    wire _T_840;
    MUX_UNSIGNED #(.width(1)) u_mux_1865 (
        .y(_T_840),
        .sel(_T_73),
        .a(1'h0),
        .b(_T_839)
    );
    wire _T_841;
    MUX_UNSIGNED #(.width(1)) u_mux_1866 (
        .y(_T_841),
        .sel(_T_69),
        .a(1'h0),
        .b(_T_840)
    );
    wire _T_842;
    MUX_UNSIGNED #(.width(1)) u_mux_1867 (
        .y(_T_842),
        .sel(_T_65),
        .a(1'h0),
        .b(_T_841)
    );
    wire _T_843;
    MUX_UNSIGNED #(.width(1)) u_mux_1868 (
        .y(_T_843),
        .sel(_T_61),
        .a(1'h0),
        .b(_T_842)
    );
    wire _T_844;
    MUX_UNSIGNED #(.width(1)) u_mux_1869 (
        .y(_T_844),
        .sel(_T_57),
        .a(1'h0),
        .b(_T_843)
    );
    wire _T_845;
    MUX_UNSIGNED #(.width(1)) u_mux_1870 (
        .y(_T_845),
        .sel(_T_53),
        .a(1'h0),
        .b(_T_844)
    );
    wire _T_846;
    MUX_UNSIGNED #(.width(1)) u_mux_1871 (
        .y(_T_846),
        .sel(_T_49),
        .a(1'h0),
        .b(_T_845)
    );
    wire _T_847;
    MUX_UNSIGNED #(.width(1)) u_mux_1872 (
        .y(_T_847),
        .sel(_T_45),
        .a(1'h0),
        .b(_T_846)
    );
    wire _T_848;
    MUX_UNSIGNED #(.width(1)) u_mux_1873 (
        .y(_T_848),
        .sel(_T_41),
        .a(1'h0),
        .b(_T_847)
    );
    wire _T_849;
    MUX_UNSIGNED #(.width(1)) u_mux_1874 (
        .y(_T_849),
        .sel(_T_37),
        .a(1'h0),
        .b(_T_848)
    );
    wire ctrlSignals_12;
    MUX_UNSIGNED #(.width(1)) u_mux_1875 (
        .y(ctrlSignals_12),
        .sel(_T_33),
        .a(1'h0),
        .b(_T_849)
    );
    wire _T_850;
    BITS #(.width(1), .high(0), .low(0)) bits_1876 (
        .y(_T_850),
        .in(ctrlSignals_6)
    );
    wire _T_851;
    BITS #(.width(1), .high(0), .low(0)) bits_1877 (
        .y(_T_851),
        .in(ctrlSignals_10)
    );
    assign io_A_sel = ctrlSignals_1;
    assign io_B_sel = ctrlSignals_2;
    assign io_alu_op = ctrlSignals_4;
    assign io_br_type = ctrlSignals_5;
    assign io_csr_cmd = ctrlSignals_11;
    assign io_illegal = ctrlSignals_12;
    assign io_imm_sel = ctrlSignals_3;
    assign io_inst_kill = _T_850;
    assign io_ld_type = ctrlSignals_8;
    assign io_pc_sel = ctrlSignals_0;
    assign io_st_type = ctrlSignals_7;
    assign io_wb_en = _T_851;
    assign io_wb_sel = ctrlSignals_9;
endmodule //Control
module RAMMEM(read_data, read_clk, read_en, read_addr, write_clk, write_en, write_mask, write_addr, write_data);
    parameter depth = 16;
    parameter addrbits = 4;
    parameter width = 32;
    parameter isSyncRead = 0;
    output [width-1:0] read_data;
    input read_clk;
    input read_en;
    input [addrbits-1:0] read_addr;
    input write_clk;
    input write_en;
    input write_mask;
    input [addrbits-1:0] write_addr;
    input [width-1:0] write_data;
    reg [width-1:0] memcore [0:depth-1];
    wire [addrbits-1:0] final_read_addr;
    generate
        if (isSyncRead) begin: raddr_processor
            reg [addrbits-1:0] read_addr_pipe_0;
            always @(posedge read_clk) begin
                if (read_en) begin
                    read_addr_pipe_0 <= read_addr;
                end
            end
            assign final_read_addr = read_addr_pipe_0;
        end else begin: raddr_processor
            assign final_read_addr = read_addr;
        end
    endgenerate
    assign read_data = memcore[final_read_addr];
    always @(posedge write_clk) begin
        if (write_en & write_mask) begin
            memcore[write_addr] <= write_data;
        end
    end
endmodule // RAMMEM
module DIV_UNSIGNED(y, num, den);
    parameter width_num = 4;
    parameter width_den = 4;
    output [width_num-1:0] y;
    input [width_num-1:0] num;
    input [width_den-1:0] den;
    assign y = num / den;
endmodule // DIV_UNSIGNED
module MUL2_UNSIGNED(y, a, b);
    parameter width_a = 4;
    parameter width_b = 4;
    output [width_a+width_b-1:0] y;
    input [width_a-1:0] a;
    input [width_b-1:0] b;
    assign y = a * b;
endmodule // MUL2_UNSIGNED
module LT_UNSIGNED(y, a, b);
    parameter width = 4;
    output y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a < b;
endmodule // LT_UNSIGNED
