module RocketCore(
    input clock,
    input reset,
    input io_interrupts_debug,
    input io_interrupts_mtip,
    input io_interrupts_msip,
    input io_interrupts_meip,
    input io_interrupts_seip,
    input [63:0] io_hartid,
    output io_imem_req_valid,
    output [39:0] io_imem_req_bits_pc,
    output io_imem_req_bits_speculative,
    output io_imem_resp_ready,
    input io_imem_resp_valid,
    input io_imem_resp_bits_btb_valid,
    input io_imem_resp_bits_btb_bits_taken,
    input [1:0] io_imem_resp_bits_btb_bits_mask,
    input io_imem_resp_bits_btb_bits_bridx,
    input [38:0] io_imem_resp_bits_btb_bits_target,
    input [5:0] io_imem_resp_bits_btb_bits_entry,
    input [6:0] io_imem_resp_bits_btb_bits_bht_history,
    input [1:0] io_imem_resp_bits_btb_bits_bht_value,
    input [39:0] io_imem_resp_bits_pc,
    input [31:0] io_imem_resp_bits_data,
    input [1:0] io_imem_resp_bits_mask,
    input io_imem_resp_bits_xcpt_if,
    input io_imem_resp_bits_replay,
    output io_imem_btb_update_valid,
    output io_imem_btb_update_bits_prediction_valid,
    output io_imem_btb_update_bits_prediction_bits_taken,
    output [1:0] io_imem_btb_update_bits_prediction_bits_mask,
    output io_imem_btb_update_bits_prediction_bits_bridx,
    output [38:0] io_imem_btb_update_bits_prediction_bits_target,
    output [5:0] io_imem_btb_update_bits_prediction_bits_entry,
    output [6:0] io_imem_btb_update_bits_prediction_bits_bht_history,
    output [1:0] io_imem_btb_update_bits_prediction_bits_bht_value,
    output [38:0] io_imem_btb_update_bits_pc,
    output [38:0] io_imem_btb_update_bits_target,
    output io_imem_btb_update_bits_taken,
    output io_imem_btb_update_bits_isValid,
    output io_imem_btb_update_bits_isJump,
    output io_imem_btb_update_bits_isReturn,
    output [38:0] io_imem_btb_update_bits_br_pc,
    output io_imem_bht_update_valid,
    output io_imem_bht_update_bits_prediction_valid,
    output io_imem_bht_update_bits_prediction_bits_taken,
    output [1:0] io_imem_bht_update_bits_prediction_bits_mask,
    output io_imem_bht_update_bits_prediction_bits_bridx,
    output [38:0] io_imem_bht_update_bits_prediction_bits_target,
    output [5:0] io_imem_bht_update_bits_prediction_bits_entry,
    output [6:0] io_imem_bht_update_bits_prediction_bits_bht_history,
    output [1:0] io_imem_bht_update_bits_prediction_bits_bht_value,
    output [38:0] io_imem_bht_update_bits_pc,
    output io_imem_bht_update_bits_taken,
    output io_imem_bht_update_bits_mispredict,
    output io_imem_ras_update_valid,
    output io_imem_ras_update_bits_isCall,
    output io_imem_ras_update_bits_isReturn,
    output [38:0] io_imem_ras_update_bits_returnAddr,
    output io_imem_ras_update_bits_prediction_valid,
    output io_imem_ras_update_bits_prediction_bits_taken,
    output [1:0] io_imem_ras_update_bits_prediction_bits_mask,
    output io_imem_ras_update_bits_prediction_bits_bridx,
    output [38:0] io_imem_ras_update_bits_prediction_bits_target,
    output [5:0] io_imem_ras_update_bits_prediction_bits_entry,
    output [6:0] io_imem_ras_update_bits_prediction_bits_bht_history,
    output [1:0] io_imem_ras_update_bits_prediction_bits_bht_value,
    output io_imem_flush_icache,
    output io_imem_flush_tlb,
    input [39:0] io_imem_npc,
    input io_imem_acquire,
    input io_dmem_req_ready,
    output io_dmem_req_valid,
    output [39:0] io_dmem_req_bits_addr,
    output [6:0] io_dmem_req_bits_tag,
    output [4:0] io_dmem_req_bits_cmd,
    output [2:0] io_dmem_req_bits_typ,
    output io_dmem_req_bits_phys,
    output [63:0] io_dmem_req_bits_data,
    output io_dmem_s1_kill,
    output [63:0] io_dmem_s1_data,
    input io_dmem_s2_nack,
    input io_dmem_acquire,
    input io_dmem_release,
    input io_dmem_resp_valid,
    input [39:0] io_dmem_resp_bits_addr,
    input [6:0] io_dmem_resp_bits_tag,
    input [4:0] io_dmem_resp_bits_cmd,
    input [2:0] io_dmem_resp_bits_typ,
    input [63:0] io_dmem_resp_bits_data,
    input io_dmem_resp_bits_replay,
    input io_dmem_resp_bits_has_data,
    input [63:0] io_dmem_resp_bits_data_word_bypass,
    input [63:0] io_dmem_resp_bits_store_data,
    input io_dmem_replay_next,
    input io_dmem_xcpt_ma_ld,
    input io_dmem_xcpt_ma_st,
    input io_dmem_xcpt_pf_ld,
    input io_dmem_xcpt_pf_st,
    output io_dmem_invalidate_lr,
    input io_dmem_ordered,
    output [3:0] io_ptw_ptbr_mode,
    output [15:0] io_ptw_ptbr_asid,
    output [43:0] io_ptw_ptbr_ppn,
    output io_ptw_invalidate,
    output io_ptw_status_debug,
    output [31:0] io_ptw_status_isa,
    output [1:0] io_ptw_status_prv,
    output io_ptw_status_sd,
    output [26:0] io_ptw_status_zero2,
    output [1:0] io_ptw_status_sxl,
    output [1:0] io_ptw_status_uxl,
    output io_ptw_status_sd_rv32,
    output [7:0] io_ptw_status_zero1,
    output io_ptw_status_tsr,
    output io_ptw_status_tw,
    output io_ptw_status_tvm,
    output io_ptw_status_mxr,
    output io_ptw_status_pum,
    output io_ptw_status_mprv,
    output [1:0] io_ptw_status_xs,
    output [1:0] io_ptw_status_fs,
    output [1:0] io_ptw_status_mpp,
    output [1:0] io_ptw_status_hpp,
    output io_ptw_status_spp,
    output io_ptw_status_mpie,
    output io_ptw_status_hpie,
    output io_ptw_status_spie,
    output io_ptw_status_upie,
    output io_ptw_status_mie,
    output io_ptw_status_hie,
    output io_ptw_status_sie,
    output io_ptw_status_uie,
    output [31:0] io_fpu_inst,
    output [63:0] io_fpu_fromint_data,
    output [2:0] io_fpu_fcsr_rm,
    input io_fpu_fcsr_flags_valid,
    input [4:0] io_fpu_fcsr_flags_bits,
    input [63:0] io_fpu_store_data,
    input [63:0] io_fpu_toint_data,
    output io_fpu_dmem_resp_val,
    output [2:0] io_fpu_dmem_resp_type,
    output [4:0] io_fpu_dmem_resp_tag,
    output [63:0] io_fpu_dmem_resp_data,
    output io_fpu_valid,
    input io_fpu_fcsr_rdy,
    input io_fpu_nack_mem,
    input io_fpu_illegal_rm,
    output io_fpu_killx,
    output io_fpu_killm,
    input [4:0] io_fpu_dec_cmd,
    input io_fpu_dec_ldst,
    input io_fpu_dec_wen,
    input io_fpu_dec_ren1,
    input io_fpu_dec_ren2,
    input io_fpu_dec_ren3,
    input io_fpu_dec_swap12,
    input io_fpu_dec_swap23,
    input io_fpu_dec_single,
    input io_fpu_dec_fromint,
    input io_fpu_dec_toint,
    input io_fpu_dec_fastpipe,
    input io_fpu_dec_fma,
    input io_fpu_dec_div,
    input io_fpu_dec_sqrt,
    input io_fpu_dec_wflags,
    input io_fpu_sboard_set,
    input io_fpu_sboard_clr,
    input [4:0] io_fpu_sboard_clra,
    input io_rocc_cmd_ready,
    output io_rocc_cmd_valid,
    output [6:0] io_rocc_cmd_bits_inst_funct,
    output [4:0] io_rocc_cmd_bits_inst_rs2,
    output [4:0] io_rocc_cmd_bits_inst_rs1,
    output io_rocc_cmd_bits_inst_xd,
    output io_rocc_cmd_bits_inst_xs1,
    output io_rocc_cmd_bits_inst_xs2,
    output [4:0] io_rocc_cmd_bits_inst_rd,
    output [6:0] io_rocc_cmd_bits_inst_opcode,
    output [63:0] io_rocc_cmd_bits_rs1,
    output [63:0] io_rocc_cmd_bits_rs2,
    output io_rocc_cmd_bits_status_debug,
    output [31:0] io_rocc_cmd_bits_status_isa,
    output [1:0] io_rocc_cmd_bits_status_prv,
    output io_rocc_cmd_bits_status_sd,
    output [26:0] io_rocc_cmd_bits_status_zero2,
    output [1:0] io_rocc_cmd_bits_status_sxl,
    output [1:0] io_rocc_cmd_bits_status_uxl,
    output io_rocc_cmd_bits_status_sd_rv32,
    output [7:0] io_rocc_cmd_bits_status_zero1,
    output io_rocc_cmd_bits_status_tsr,
    output io_rocc_cmd_bits_status_tw,
    output io_rocc_cmd_bits_status_tvm,
    output io_rocc_cmd_bits_status_mxr,
    output io_rocc_cmd_bits_status_pum,
    output io_rocc_cmd_bits_status_mprv,
    output [1:0] io_rocc_cmd_bits_status_xs,
    output [1:0] io_rocc_cmd_bits_status_fs,
    output [1:0] io_rocc_cmd_bits_status_mpp,
    output [1:0] io_rocc_cmd_bits_status_hpp,
    output io_rocc_cmd_bits_status_spp,
    output io_rocc_cmd_bits_status_mpie,
    output io_rocc_cmd_bits_status_hpie,
    output io_rocc_cmd_bits_status_spie,
    output io_rocc_cmd_bits_status_upie,
    output io_rocc_cmd_bits_status_mie,
    output io_rocc_cmd_bits_status_hie,
    output io_rocc_cmd_bits_status_sie,
    output io_rocc_cmd_bits_status_uie,
    output io_rocc_resp_ready,
    input io_rocc_resp_valid,
    input [4:0] io_rocc_resp_bits_rd,
    input [63:0] io_rocc_resp_bits_data,
    output io_rocc_mem_req_ready,
    input io_rocc_mem_req_valid,
    input [39:0] io_rocc_mem_req_bits_addr,
    input [6:0] io_rocc_mem_req_bits_tag,
    input [4:0] io_rocc_mem_req_bits_cmd,
    input [2:0] io_rocc_mem_req_bits_typ,
    input io_rocc_mem_req_bits_phys,
    input [63:0] io_rocc_mem_req_bits_data,
    input io_rocc_mem_s1_kill,
    input [63:0] io_rocc_mem_s1_data,
    output io_rocc_mem_s2_nack,
    output io_rocc_mem_acquire,
    output io_rocc_mem_release,
    output io_rocc_mem_resp_valid,
    output [39:0] io_rocc_mem_resp_bits_addr,
    output [6:0] io_rocc_mem_resp_bits_tag,
    output [4:0] io_rocc_mem_resp_bits_cmd,
    output [2:0] io_rocc_mem_resp_bits_typ,
    output [63:0] io_rocc_mem_resp_bits_data,
    output io_rocc_mem_resp_bits_replay,
    output io_rocc_mem_resp_bits_has_data,
    output [63:0] io_rocc_mem_resp_bits_data_word_bypass,
    output [63:0] io_rocc_mem_resp_bits_store_data,
    output io_rocc_mem_replay_next,
    output io_rocc_mem_xcpt_ma_ld,
    output io_rocc_mem_xcpt_ma_st,
    output io_rocc_mem_xcpt_pf_ld,
    output io_rocc_mem_xcpt_pf_st,
    input io_rocc_mem_invalidate_lr,
    output io_rocc_mem_ordered,
    input io_rocc_busy,
    input io_rocc_interrupt,
    output io_rocc_exception
);
    wire _ex_ctrl_fp__q;
    wire _ex_ctrl_fp__d;
    DFF_POSCLK #(.width(1)) ex_ctrl_fp (
        .q(_ex_ctrl_fp__q),
        .d(_ex_ctrl_fp__d),
        .clk(clock)
    );
    wire _ex_ctrl_branch__q;
    wire _ex_ctrl_branch__d;
    DFF_POSCLK #(.width(1)) ex_ctrl_branch (
        .q(_ex_ctrl_branch__q),
        .d(_ex_ctrl_branch__d),
        .clk(clock)
    );
    wire _ex_ctrl_jal__q;
    wire _ex_ctrl_jal__d;
    DFF_POSCLK #(.width(1)) ex_ctrl_jal (
        .q(_ex_ctrl_jal__q),
        .d(_ex_ctrl_jal__d),
        .clk(clock)
    );
    wire _ex_ctrl_jalr__q;
    wire _ex_ctrl_jalr__d;
    DFF_POSCLK #(.width(1)) ex_ctrl_jalr (
        .q(_ex_ctrl_jalr__q),
        .d(_ex_ctrl_jalr__d),
        .clk(clock)
    );
    wire _ex_ctrl_rxs2__q;
    wire _ex_ctrl_rxs2__d;
    DFF_POSCLK #(.width(1)) ex_ctrl_rxs2 (
        .q(_ex_ctrl_rxs2__q),
        .d(_ex_ctrl_rxs2__d),
        .clk(clock)
    );
    wire [1:0] _ex_ctrl_sel_alu2__q;
    wire [1:0] _ex_ctrl_sel_alu2__d;
    DFF_POSCLK #(.width(2)) ex_ctrl_sel_alu2 (
        .q(_ex_ctrl_sel_alu2__q),
        .d(_ex_ctrl_sel_alu2__d),
        .clk(clock)
    );
    wire [1:0] _ex_ctrl_sel_alu1__q;
    wire [1:0] _ex_ctrl_sel_alu1__d;
    DFF_POSCLK #(.width(2)) ex_ctrl_sel_alu1 (
        .q(_ex_ctrl_sel_alu1__q),
        .d(_ex_ctrl_sel_alu1__d),
        .clk(clock)
    );
    wire [2:0] _ex_ctrl_sel_imm__q;
    wire [2:0] _ex_ctrl_sel_imm__d;
    DFF_POSCLK #(.width(3)) ex_ctrl_sel_imm (
        .q(_ex_ctrl_sel_imm__q),
        .d(_ex_ctrl_sel_imm__d),
        .clk(clock)
    );
    wire _ex_ctrl_alu_dw__q;
    wire _ex_ctrl_alu_dw__d;
    DFF_POSCLK #(.width(1)) ex_ctrl_alu_dw (
        .q(_ex_ctrl_alu_dw__q),
        .d(_ex_ctrl_alu_dw__d),
        .clk(clock)
    );
    wire [3:0] _ex_ctrl_alu_fn__q;
    wire [3:0] _ex_ctrl_alu_fn__d;
    DFF_POSCLK #(.width(4)) ex_ctrl_alu_fn (
        .q(_ex_ctrl_alu_fn__q),
        .d(_ex_ctrl_alu_fn__d),
        .clk(clock)
    );
    wire _ex_ctrl_mem__q;
    wire _ex_ctrl_mem__d;
    DFF_POSCLK #(.width(1)) ex_ctrl_mem (
        .q(_ex_ctrl_mem__q),
        .d(_ex_ctrl_mem__d),
        .clk(clock)
    );
    wire [4:0] _ex_ctrl_mem_cmd__q;
    wire [4:0] _ex_ctrl_mem_cmd__d;
    DFF_POSCLK #(.width(5)) ex_ctrl_mem_cmd (
        .q(_ex_ctrl_mem_cmd__q),
        .d(_ex_ctrl_mem_cmd__d),
        .clk(clock)
    );
    wire [2:0] _ex_ctrl_mem_type__q;
    wire [2:0] _ex_ctrl_mem_type__d;
    DFF_POSCLK #(.width(3)) ex_ctrl_mem_type (
        .q(_ex_ctrl_mem_type__q),
        .d(_ex_ctrl_mem_type__d),
        .clk(clock)
    );
    wire _ex_ctrl_wfd__q;
    wire _ex_ctrl_wfd__d;
    DFF_POSCLK #(.width(1)) ex_ctrl_wfd (
        .q(_ex_ctrl_wfd__q),
        .d(_ex_ctrl_wfd__d),
        .clk(clock)
    );
    wire _ex_ctrl_div__q;
    wire _ex_ctrl_div__d;
    DFF_POSCLK #(.width(1)) ex_ctrl_div (
        .q(_ex_ctrl_div__q),
        .d(_ex_ctrl_div__d),
        .clk(clock)
    );
    wire _ex_ctrl_wxd__q;
    wire _ex_ctrl_wxd__d;
    DFF_POSCLK #(.width(1)) ex_ctrl_wxd (
        .q(_ex_ctrl_wxd__q),
        .d(_ex_ctrl_wxd__d),
        .clk(clock)
    );
    wire [2:0] _ex_ctrl_csr__q;
    wire [2:0] _ex_ctrl_csr__d;
    DFF_POSCLK #(.width(3)) ex_ctrl_csr (
        .q(_ex_ctrl_csr__q),
        .d(_ex_ctrl_csr__d),
        .clk(clock)
    );
    wire _ex_ctrl_fence_i__q;
    wire _ex_ctrl_fence_i__d;
    DFF_POSCLK #(.width(1)) ex_ctrl_fence_i (
        .q(_ex_ctrl_fence_i__q),
        .d(_ex_ctrl_fence_i__d),
        .clk(clock)
    );
    wire _mem_ctrl_fp__q;
    wire _mem_ctrl_fp__d;
    DFF_POSCLK #(.width(1)) mem_ctrl_fp (
        .q(_mem_ctrl_fp__q),
        .d(_mem_ctrl_fp__d),
        .clk(clock)
    );
    wire _mem_ctrl_branch__q;
    wire _mem_ctrl_branch__d;
    DFF_POSCLK #(.width(1)) mem_ctrl_branch (
        .q(_mem_ctrl_branch__q),
        .d(_mem_ctrl_branch__d),
        .clk(clock)
    );
    wire _mem_ctrl_jal__q;
    wire _mem_ctrl_jal__d;
    DFF_POSCLK #(.width(1)) mem_ctrl_jal (
        .q(_mem_ctrl_jal__q),
        .d(_mem_ctrl_jal__d),
        .clk(clock)
    );
    wire _mem_ctrl_jalr__q;
    wire _mem_ctrl_jalr__d;
    DFF_POSCLK #(.width(1)) mem_ctrl_jalr (
        .q(_mem_ctrl_jalr__q),
        .d(_mem_ctrl_jalr__d),
        .clk(clock)
    );
    wire _mem_ctrl_mem__q;
    wire _mem_ctrl_mem__d;
    DFF_POSCLK #(.width(1)) mem_ctrl_mem (
        .q(_mem_ctrl_mem__q),
        .d(_mem_ctrl_mem__d),
        .clk(clock)
    );
    wire _mem_ctrl_wfd__q;
    wire _mem_ctrl_wfd__d;
    DFF_POSCLK #(.width(1)) mem_ctrl_wfd (
        .q(_mem_ctrl_wfd__q),
        .d(_mem_ctrl_wfd__d),
        .clk(clock)
    );
    wire _mem_ctrl_div__q;
    wire _mem_ctrl_div__d;
    DFF_POSCLK #(.width(1)) mem_ctrl_div (
        .q(_mem_ctrl_div__q),
        .d(_mem_ctrl_div__d),
        .clk(clock)
    );
    wire _mem_ctrl_wxd__q;
    wire _mem_ctrl_wxd__d;
    DFF_POSCLK #(.width(1)) mem_ctrl_wxd (
        .q(_mem_ctrl_wxd__q),
        .d(_mem_ctrl_wxd__d),
        .clk(clock)
    );
    wire [2:0] _mem_ctrl_csr__q;
    wire [2:0] _mem_ctrl_csr__d;
    DFF_POSCLK #(.width(3)) mem_ctrl_csr (
        .q(_mem_ctrl_csr__q),
        .d(_mem_ctrl_csr__d),
        .clk(clock)
    );
    wire _mem_ctrl_fence_i__q;
    wire _mem_ctrl_fence_i__d;
    DFF_POSCLK #(.width(1)) mem_ctrl_fence_i (
        .q(_mem_ctrl_fence_i__q),
        .d(_mem_ctrl_fence_i__d),
        .clk(clock)
    );
    wire _wb_ctrl_mem__q;
    wire _wb_ctrl_mem__d;
    DFF_POSCLK #(.width(1)) wb_ctrl_mem (
        .q(_wb_ctrl_mem__q),
        .d(_wb_ctrl_mem__d),
        .clk(clock)
    );
    wire _wb_ctrl_wfd__q;
    wire _wb_ctrl_wfd__d;
    DFF_POSCLK #(.width(1)) wb_ctrl_wfd (
        .q(_wb_ctrl_wfd__q),
        .d(_wb_ctrl_wfd__d),
        .clk(clock)
    );
    wire _wb_ctrl_div__q;
    wire _wb_ctrl_div__d;
    DFF_POSCLK #(.width(1)) wb_ctrl_div (
        .q(_wb_ctrl_div__q),
        .d(_wb_ctrl_div__d),
        .clk(clock)
    );
    wire _wb_ctrl_wxd__q;
    wire _wb_ctrl_wxd__d;
    DFF_POSCLK #(.width(1)) wb_ctrl_wxd (
        .q(_wb_ctrl_wxd__q),
        .d(_wb_ctrl_wxd__d),
        .clk(clock)
    );
    wire [2:0] _wb_ctrl_csr__q;
    wire [2:0] _wb_ctrl_csr__d;
    DFF_POSCLK #(.width(3)) wb_ctrl_csr (
        .q(_wb_ctrl_csr__q),
        .d(_wb_ctrl_csr__d),
        .clk(clock)
    );
    wire _wb_ctrl_fence_i__q;
    wire _wb_ctrl_fence_i__d;
    DFF_POSCLK #(.width(1)) wb_ctrl_fence_i (
        .q(_wb_ctrl_fence_i__q),
        .d(_wb_ctrl_fence_i__d),
        .clk(clock)
    );
    wire _ex_reg_xcpt_interrupt__q;
    wire _ex_reg_xcpt_interrupt__d;
    DFF_POSCLK #(.width(1)) ex_reg_xcpt_interrupt (
        .q(_ex_reg_xcpt_interrupt__q),
        .d(_ex_reg_xcpt_interrupt__d),
        .clk(clock)
    );
    wire _ex_reg_valid__q;
    wire _ex_reg_valid__d;
    DFF_POSCLK #(.width(1)) ex_reg_valid (
        .q(_ex_reg_valid__q),
        .d(_ex_reg_valid__d),
        .clk(clock)
    );
    wire _ex_reg_rvc__q;
    wire _ex_reg_rvc__d;
    DFF_POSCLK #(.width(1)) ex_reg_rvc (
        .q(_ex_reg_rvc__q),
        .d(_ex_reg_rvc__d),
        .clk(clock)
    );
    wire _ex_reg_btb_hit__q;
    wire _ex_reg_btb_hit__d;
    DFF_POSCLK #(.width(1)) ex_reg_btb_hit (
        .q(_ex_reg_btb_hit__q),
        .d(_ex_reg_btb_hit__d),
        .clk(clock)
    );
    wire _ex_reg_btb_resp_taken__q;
    wire _ex_reg_btb_resp_taken__d;
    DFF_POSCLK #(.width(1)) ex_reg_btb_resp_taken (
        .q(_ex_reg_btb_resp_taken__q),
        .d(_ex_reg_btb_resp_taken__d),
        .clk(clock)
    );
    wire [1:0] _ex_reg_btb_resp_mask__q;
    wire [1:0] _ex_reg_btb_resp_mask__d;
    DFF_POSCLK #(.width(2)) ex_reg_btb_resp_mask (
        .q(_ex_reg_btb_resp_mask__q),
        .d(_ex_reg_btb_resp_mask__d),
        .clk(clock)
    );
    wire _ex_reg_btb_resp_bridx__q;
    wire _ex_reg_btb_resp_bridx__d;
    DFF_POSCLK #(.width(1)) ex_reg_btb_resp_bridx (
        .q(_ex_reg_btb_resp_bridx__q),
        .d(_ex_reg_btb_resp_bridx__d),
        .clk(clock)
    );
    wire [38:0] _ex_reg_btb_resp_target__q;
    wire [38:0] _ex_reg_btb_resp_target__d;
    DFF_POSCLK #(.width(39)) ex_reg_btb_resp_target (
        .q(_ex_reg_btb_resp_target__q),
        .d(_ex_reg_btb_resp_target__d),
        .clk(clock)
    );
    wire [5:0] _ex_reg_btb_resp_entry__q;
    wire [5:0] _ex_reg_btb_resp_entry__d;
    DFF_POSCLK #(.width(6)) ex_reg_btb_resp_entry (
        .q(_ex_reg_btb_resp_entry__q),
        .d(_ex_reg_btb_resp_entry__d),
        .clk(clock)
    );
    wire [6:0] _ex_reg_btb_resp_bht_history__q;
    wire [6:0] _ex_reg_btb_resp_bht_history__d;
    DFF_POSCLK #(.width(7)) ex_reg_btb_resp_bht_history (
        .q(_ex_reg_btb_resp_bht_history__q),
        .d(_ex_reg_btb_resp_bht_history__d),
        .clk(clock)
    );
    wire [1:0] _ex_reg_btb_resp_bht_value__q;
    wire [1:0] _ex_reg_btb_resp_bht_value__d;
    DFF_POSCLK #(.width(2)) ex_reg_btb_resp_bht_value (
        .q(_ex_reg_btb_resp_bht_value__q),
        .d(_ex_reg_btb_resp_bht_value__d),
        .clk(clock)
    );
    wire _ex_reg_xcpt__q;
    wire _ex_reg_xcpt__d;
    DFF_POSCLK #(.width(1)) ex_reg_xcpt (
        .q(_ex_reg_xcpt__q),
        .d(_ex_reg_xcpt__d),
        .clk(clock)
    );
    wire _ex_reg_flush_pipe__q;
    wire _ex_reg_flush_pipe__d;
    DFF_POSCLK #(.width(1)) ex_reg_flush_pipe (
        .q(_ex_reg_flush_pipe__q),
        .d(_ex_reg_flush_pipe__d),
        .clk(clock)
    );
    wire _ex_reg_load_use__q;
    wire _ex_reg_load_use__d;
    DFF_POSCLK #(.width(1)) ex_reg_load_use (
        .q(_ex_reg_load_use__q),
        .d(_ex_reg_load_use__d),
        .clk(clock)
    );
    wire [63:0] _ex_cause__q;
    wire [63:0] _ex_cause__d;
    DFF_POSCLK #(.width(64)) ex_cause (
        .q(_ex_cause__q),
        .d(_ex_cause__d),
        .clk(clock)
    );
    wire _ex_reg_replay__q;
    wire _ex_reg_replay__d;
    DFF_POSCLK #(.width(1)) ex_reg_replay (
        .q(_ex_reg_replay__q),
        .d(_ex_reg_replay__d),
        .clk(clock)
    );
    wire [39:0] _ex_reg_pc__q;
    wire [39:0] _ex_reg_pc__d;
    DFF_POSCLK #(.width(40)) ex_reg_pc (
        .q(_ex_reg_pc__q),
        .d(_ex_reg_pc__d),
        .clk(clock)
    );
    wire [31:0] _ex_reg_inst__q;
    wire [31:0] _ex_reg_inst__d;
    DFF_POSCLK #(.width(32)) ex_reg_inst (
        .q(_ex_reg_inst__q),
        .d(_ex_reg_inst__d),
        .clk(clock)
    );
    wire _mem_reg_xcpt_interrupt__q;
    wire _mem_reg_xcpt_interrupt__d;
    DFF_POSCLK #(.width(1)) mem_reg_xcpt_interrupt (
        .q(_mem_reg_xcpt_interrupt__q),
        .d(_mem_reg_xcpt_interrupt__d),
        .clk(clock)
    );
    wire _mem_reg_valid__q;
    wire _mem_reg_valid__d;
    DFF_POSCLK #(.width(1)) mem_reg_valid (
        .q(_mem_reg_valid__q),
        .d(_mem_reg_valid__d),
        .clk(clock)
    );
    wire _mem_reg_rvc__q;
    wire _mem_reg_rvc__d;
    DFF_POSCLK #(.width(1)) mem_reg_rvc (
        .q(_mem_reg_rvc__q),
        .d(_mem_reg_rvc__d),
        .clk(clock)
    );
    wire _mem_reg_btb_hit__q;
    wire _mem_reg_btb_hit__d;
    DFF_POSCLK #(.width(1)) mem_reg_btb_hit (
        .q(_mem_reg_btb_hit__q),
        .d(_mem_reg_btb_hit__d),
        .clk(clock)
    );
    wire _mem_reg_btb_resp_taken__q;
    wire _mem_reg_btb_resp_taken__d;
    DFF_POSCLK #(.width(1)) mem_reg_btb_resp_taken (
        .q(_mem_reg_btb_resp_taken__q),
        .d(_mem_reg_btb_resp_taken__d),
        .clk(clock)
    );
    wire [1:0] _mem_reg_btb_resp_mask__q;
    wire [1:0] _mem_reg_btb_resp_mask__d;
    DFF_POSCLK #(.width(2)) mem_reg_btb_resp_mask (
        .q(_mem_reg_btb_resp_mask__q),
        .d(_mem_reg_btb_resp_mask__d),
        .clk(clock)
    );
    wire _mem_reg_btb_resp_bridx__q;
    wire _mem_reg_btb_resp_bridx__d;
    DFF_POSCLK #(.width(1)) mem_reg_btb_resp_bridx (
        .q(_mem_reg_btb_resp_bridx__q),
        .d(_mem_reg_btb_resp_bridx__d),
        .clk(clock)
    );
    wire [38:0] _mem_reg_btb_resp_target__q;
    wire [38:0] _mem_reg_btb_resp_target__d;
    DFF_POSCLK #(.width(39)) mem_reg_btb_resp_target (
        .q(_mem_reg_btb_resp_target__q),
        .d(_mem_reg_btb_resp_target__d),
        .clk(clock)
    );
    wire [5:0] _mem_reg_btb_resp_entry__q;
    wire [5:0] _mem_reg_btb_resp_entry__d;
    DFF_POSCLK #(.width(6)) mem_reg_btb_resp_entry (
        .q(_mem_reg_btb_resp_entry__q),
        .d(_mem_reg_btb_resp_entry__d),
        .clk(clock)
    );
    wire [6:0] _mem_reg_btb_resp_bht_history__q;
    wire [6:0] _mem_reg_btb_resp_bht_history__d;
    DFF_POSCLK #(.width(7)) mem_reg_btb_resp_bht_history (
        .q(_mem_reg_btb_resp_bht_history__q),
        .d(_mem_reg_btb_resp_bht_history__d),
        .clk(clock)
    );
    wire [1:0] _mem_reg_btb_resp_bht_value__q;
    wire [1:0] _mem_reg_btb_resp_bht_value__d;
    DFF_POSCLK #(.width(2)) mem_reg_btb_resp_bht_value (
        .q(_mem_reg_btb_resp_bht_value__q),
        .d(_mem_reg_btb_resp_bht_value__d),
        .clk(clock)
    );
    wire _mem_reg_xcpt__q;
    wire _mem_reg_xcpt__d;
    DFF_POSCLK #(.width(1)) mem_reg_xcpt (
        .q(_mem_reg_xcpt__q),
        .d(_mem_reg_xcpt__d),
        .clk(clock)
    );
    wire _mem_reg_replay__q;
    wire _mem_reg_replay__d;
    DFF_POSCLK #(.width(1)) mem_reg_replay (
        .q(_mem_reg_replay__q),
        .d(_mem_reg_replay__d),
        .clk(clock)
    );
    wire _mem_reg_flush_pipe__q;
    wire _mem_reg_flush_pipe__d;
    DFF_POSCLK #(.width(1)) mem_reg_flush_pipe (
        .q(_mem_reg_flush_pipe__q),
        .d(_mem_reg_flush_pipe__d),
        .clk(clock)
    );
    wire [63:0] _mem_reg_cause__q;
    wire [63:0] _mem_reg_cause__d;
    DFF_POSCLK #(.width(64)) mem_reg_cause (
        .q(_mem_reg_cause__q),
        .d(_mem_reg_cause__d),
        .clk(clock)
    );
    wire _mem_reg_slow_bypass__q;
    wire _mem_reg_slow_bypass__d;
    DFF_POSCLK #(.width(1)) mem_reg_slow_bypass (
        .q(_mem_reg_slow_bypass__q),
        .d(_mem_reg_slow_bypass__d),
        .clk(clock)
    );
    wire _mem_reg_load__q;
    wire _mem_reg_load__d;
    DFF_POSCLK #(.width(1)) mem_reg_load (
        .q(_mem_reg_load__q),
        .d(_mem_reg_load__d),
        .clk(clock)
    );
    wire _mem_reg_store__q;
    wire _mem_reg_store__d;
    DFF_POSCLK #(.width(1)) mem_reg_store (
        .q(_mem_reg_store__q),
        .d(_mem_reg_store__d),
        .clk(clock)
    );
    wire [39:0] _mem_reg_pc__q;
    wire [39:0] _mem_reg_pc__d;
    DFF_POSCLK #(.width(40)) mem_reg_pc (
        .q(_mem_reg_pc__q),
        .d(_mem_reg_pc__d),
        .clk(clock)
    );
    wire [31:0] _mem_reg_inst__q;
    wire [31:0] _mem_reg_inst__d;
    DFF_POSCLK #(.width(32)) mem_reg_inst (
        .q(_mem_reg_inst__q),
        .d(_mem_reg_inst__d),
        .clk(clock)
    );
    wire [63:0] _mem_reg_wdata__q;
    wire [63:0] _mem_reg_wdata__d;
    DFF_POSCLK #(.width(64)) mem_reg_wdata (
        .q(_mem_reg_wdata__q),
        .d(_mem_reg_wdata__d),
        .clk(clock)
    );
    wire [63:0] _mem_reg_rs2__q;
    wire [63:0] _mem_reg_rs2__d;
    DFF_POSCLK #(.width(64)) mem_reg_rs2 (
        .q(_mem_reg_rs2__q),
        .d(_mem_reg_rs2__d),
        .clk(clock)
    );
    wire take_pc_mem;
    wire _wb_reg_valid__q;
    wire _wb_reg_valid__d;
    DFF_POSCLK #(.width(1)) wb_reg_valid (
        .q(_wb_reg_valid__q),
        .d(_wb_reg_valid__d),
        .clk(clock)
    );
    wire _wb_reg_xcpt__q;
    wire _wb_reg_xcpt__d;
    DFF_POSCLK #(.width(1)) wb_reg_xcpt (
        .q(_wb_reg_xcpt__q),
        .d(_wb_reg_xcpt__d),
        .clk(clock)
    );
    wire _wb_reg_replay__q;
    wire _wb_reg_replay__d;
    DFF_POSCLK #(.width(1)) wb_reg_replay (
        .q(_wb_reg_replay__q),
        .d(_wb_reg_replay__d),
        .clk(clock)
    );
    wire [63:0] _wb_reg_cause__q;
    wire [63:0] _wb_reg_cause__d;
    DFF_POSCLK #(.width(64)) wb_reg_cause (
        .q(_wb_reg_cause__q),
        .d(_wb_reg_cause__d),
        .clk(clock)
    );
    wire [39:0] _wb_reg_pc__q;
    wire [39:0] _wb_reg_pc__d;
    DFF_POSCLK #(.width(40)) wb_reg_pc (
        .q(_wb_reg_pc__q),
        .d(_wb_reg_pc__d),
        .clk(clock)
    );
    wire [31:0] _wb_reg_inst__q;
    wire [31:0] _wb_reg_inst__d;
    DFF_POSCLK #(.width(32)) wb_reg_inst (
        .q(_wb_reg_inst__q),
        .d(_wb_reg_inst__d),
        .clk(clock)
    );
    wire [63:0] _wb_reg_wdata__q;
    wire [63:0] _wb_reg_wdata__d;
    DFF_POSCLK #(.width(64)) wb_reg_wdata (
        .q(_wb_reg_wdata__q),
        .d(_wb_reg_wdata__d),
        .clk(clock)
    );
    wire take_pc_wb;
    wire take_pc_id;
    wire take_pc_mem_wb;
    BITWISEOR #(.width(1)) bitwiseor_1 (
        .y(take_pc_mem_wb),
        .a(take_pc_wb),
        .b(take_pc_mem)
    );
    wire take_pc;
    BITWISEOR #(.width(1)) bitwiseor_2 (
        .y(take_pc),
        .a(take_pc_mem_wb),
        .b(take_pc_id)
    );
    wire _ibuf__clock;
    wire _ibuf__reset;
    wire _ibuf__io_imem_ready;
    wire _ibuf__io_imem_valid;
    wire _ibuf__io_imem_bits_btb_valid;
    wire _ibuf__io_imem_bits_btb_bits_taken;
    wire [1:0] _ibuf__io_imem_bits_btb_bits_mask;
    wire _ibuf__io_imem_bits_btb_bits_bridx;
    wire [38:0] _ibuf__io_imem_bits_btb_bits_target;
    wire [5:0] _ibuf__io_imem_bits_btb_bits_entry;
    wire [6:0] _ibuf__io_imem_bits_btb_bits_bht_history;
    wire [1:0] _ibuf__io_imem_bits_btb_bits_bht_value;
    wire [39:0] _ibuf__io_imem_bits_pc;
    wire [31:0] _ibuf__io_imem_bits_data;
    wire [1:0] _ibuf__io_imem_bits_mask;
    wire _ibuf__io_imem_bits_xcpt_if;
    wire _ibuf__io_imem_bits_replay;
    wire _ibuf__io_kill;
    wire [39:0] _ibuf__io_pc;
    wire _ibuf__io_btb_resp_taken;
    wire [1:0] _ibuf__io_btb_resp_mask;
    wire _ibuf__io_btb_resp_bridx;
    wire [38:0] _ibuf__io_btb_resp_target;
    wire [5:0] _ibuf__io_btb_resp_entry;
    wire [6:0] _ibuf__io_btb_resp_bht_history;
    wire [1:0] _ibuf__io_btb_resp_bht_value;
    wire _ibuf__io_inst_0_ready;
    wire _ibuf__io_inst_0_valid;
    wire _ibuf__io_inst_0_bits_pf0;
    wire _ibuf__io_inst_0_bits_pf1;
    wire _ibuf__io_inst_0_bits_replay;
    wire _ibuf__io_inst_0_bits_btb_hit;
    wire _ibuf__io_inst_0_bits_rvc;
    wire [31:0] _ibuf__io_inst_0_bits_inst_bits;
    wire [4:0] _ibuf__io_inst_0_bits_inst_rd;
    wire [4:0] _ibuf__io_inst_0_bits_inst_rs1;
    wire [4:0] _ibuf__io_inst_0_bits_inst_rs2;
    wire [4:0] _ibuf__io_inst_0_bits_inst_rs3;
    wire [31:0] _ibuf__io_inst_0_bits_raw;
    IBuf ibuf (
        .clock(_ibuf__clock),
        .reset(_ibuf__reset),
        .io_imem_ready(_ibuf__io_imem_ready),
        .io_imem_valid(_ibuf__io_imem_valid),
        .io_imem_bits_btb_valid(_ibuf__io_imem_bits_btb_valid),
        .io_imem_bits_btb_bits_taken(_ibuf__io_imem_bits_btb_bits_taken),
        .io_imem_bits_btb_bits_mask(_ibuf__io_imem_bits_btb_bits_mask),
        .io_imem_bits_btb_bits_bridx(_ibuf__io_imem_bits_btb_bits_bridx),
        .io_imem_bits_btb_bits_target(_ibuf__io_imem_bits_btb_bits_target),
        .io_imem_bits_btb_bits_entry(_ibuf__io_imem_bits_btb_bits_entry),
        .io_imem_bits_btb_bits_bht_history(_ibuf__io_imem_bits_btb_bits_bht_history),
        .io_imem_bits_btb_bits_bht_value(_ibuf__io_imem_bits_btb_bits_bht_value),
        .io_imem_bits_pc(_ibuf__io_imem_bits_pc),
        .io_imem_bits_data(_ibuf__io_imem_bits_data),
        .io_imem_bits_mask(_ibuf__io_imem_bits_mask),
        .io_imem_bits_xcpt_if(_ibuf__io_imem_bits_xcpt_if),
        .io_imem_bits_replay(_ibuf__io_imem_bits_replay),
        .io_kill(_ibuf__io_kill),
        .io_pc(_ibuf__io_pc),
        .io_btb_resp_taken(_ibuf__io_btb_resp_taken),
        .io_btb_resp_mask(_ibuf__io_btb_resp_mask),
        .io_btb_resp_bridx(_ibuf__io_btb_resp_bridx),
        .io_btb_resp_target(_ibuf__io_btb_resp_target),
        .io_btb_resp_entry(_ibuf__io_btb_resp_entry),
        .io_btb_resp_bht_history(_ibuf__io_btb_resp_bht_history),
        .io_btb_resp_bht_value(_ibuf__io_btb_resp_bht_value),
        .io_inst_0_ready(_ibuf__io_inst_0_ready),
        .io_inst_0_valid(_ibuf__io_inst_0_valid),
        .io_inst_0_bits_pf0(_ibuf__io_inst_0_bits_pf0),
        .io_inst_0_bits_pf1(_ibuf__io_inst_0_bits_pf1),
        .io_inst_0_bits_replay(_ibuf__io_inst_0_bits_replay),
        .io_inst_0_bits_btb_hit(_ibuf__io_inst_0_bits_btb_hit),
        .io_inst_0_bits_rvc(_ibuf__io_inst_0_bits_rvc),
        .io_inst_0_bits_inst_bits(_ibuf__io_inst_0_bits_inst_bits),
        .io_inst_0_bits_inst_rd(_ibuf__io_inst_0_bits_inst_rd),
        .io_inst_0_bits_inst_rs1(_ibuf__io_inst_0_bits_inst_rs1),
        .io_inst_0_bits_inst_rs2(_ibuf__io_inst_0_bits_inst_rs2),
        .io_inst_0_bits_inst_rs3(_ibuf__io_inst_0_bits_inst_rs3),
        .io_inst_0_bits_raw(_ibuf__io_inst_0_bits_raw)
    );
    wire id_ctrl_legal;
    wire id_ctrl_fp;
    wire id_ctrl_rocc;
    wire id_ctrl_branch;
    wire id_ctrl_jal;
    wire id_ctrl_jalr;
    wire id_ctrl_rxs2;
    wire id_ctrl_rxs1;
    wire [1:0] id_ctrl_sel_alu2;
    wire [1:0] id_ctrl_sel_alu1;
    wire [2:0] id_ctrl_sel_imm;
    wire id_ctrl_alu_dw;
    wire [3:0] id_ctrl_alu_fn;
    wire id_ctrl_mem;
    wire [4:0] id_ctrl_mem_cmd;
    wire [2:0] id_ctrl_mem_type;
    wire id_ctrl_rfs1;
    wire id_ctrl_rfs2;
    wire id_ctrl_rfs3;
    wire id_ctrl_wfd;
    wire id_ctrl_div;
    wire id_ctrl_wxd;
    wire [2:0] id_ctrl_csr;
    wire id_ctrl_fence_i;
    wire id_ctrl_fence;
    wire id_ctrl_amo;
    wire id_ctrl_dp;
    wire [31:0] _T_2603;
    BITWISEAND #(.width(32)) bitwiseand_1353 (
        .y(_T_2603),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h207F)
    );
    wire _T_2605;
    EQ_UNSIGNED #(.width(32)) u_eq_1354 (
        .y(_T_2605),
        .a(_T_2603),
        .b(32'h3)
    );
    wire [31:0] _T_2607;
    BITWISEAND #(.width(32)) bitwiseand_1355 (
        .y(_T_2607),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h106F)
    );
    wire _T_2609;
    EQ_UNSIGNED #(.width(32)) u_eq_1356 (
        .y(_T_2609),
        .a(_T_2607),
        .b(32'h3)
    );
    wire [31:0] _T_2611;
    BITWISEAND #(.width(32)) bitwiseand_1357 (
        .y(_T_2611),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h607F)
    );
    wire _T_2613;
    EQ_UNSIGNED #(.width(32)) u_eq_1358 (
        .y(_T_2613),
        .a(_T_2611),
        .b(32'hF)
    );
    wire [31:0] _T_2615;
    BITWISEAND #(.width(32)) bitwiseand_1359 (
        .y(_T_2615),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h7077)
    );
    wire _T_2617;
    EQ_UNSIGNED #(.width(32)) u_eq_1360 (
        .y(_T_2617),
        .a(_T_2615),
        .b(32'h13)
    );
    wire [31:0] _T_2619;
    BITWISEAND #(.width(32)) bitwiseand_1361 (
        .y(_T_2619),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h5F)
    );
    wire _T_2621;
    EQ_UNSIGNED #(.width(32)) u_eq_1362 (
        .y(_T_2621),
        .a(_T_2619),
        .b(32'h17)
    );
    wire [31:0] _T_2623;
    BITWISEAND #(.width(32)) bitwiseand_1363 (
        .y(_T_2623),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'hFC00007F)
    );
    wire _T_2625;
    EQ_UNSIGNED #(.width(32)) u_eq_1364 (
        .y(_T_2625),
        .a(_T_2623),
        .b(32'h33)
    );
    wire [31:0] _T_2627;
    BITWISEAND #(.width(32)) bitwiseand_1365 (
        .y(_T_2627),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'hBE007077)
    );
    wire _T_2629;
    EQ_UNSIGNED #(.width(32)) u_eq_1366 (
        .y(_T_2629),
        .a(_T_2627),
        .b(32'h33)
    );
    wire [31:0] _T_2631;
    BITWISEAND #(.width(32)) bitwiseand_1367 (
        .y(_T_2631),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h4000073)
    );
    wire _T_2633;
    EQ_UNSIGNED #(.width(32)) u_eq_1368 (
        .y(_T_2633),
        .a(_T_2631),
        .b(32'h43)
    );
    wire [31:0] _T_2635;
    BITWISEAND #(.width(32)) bitwiseand_1369 (
        .y(_T_2635),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'hE400007F)
    );
    wire _T_2637;
    EQ_UNSIGNED #(.width(32)) u_eq_1370 (
        .y(_T_2637),
        .a(_T_2635),
        .b(32'h53)
    );
    wire [31:0] _T_2639;
    BITWISEAND #(.width(32)) bitwiseand_1371 (
        .y(_T_2639),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h707B)
    );
    wire _T_2641;
    EQ_UNSIGNED #(.width(32)) u_eq_1372 (
        .y(_T_2641),
        .a(_T_2639),
        .b(32'h63)
    );
    wire [31:0] _T_2643;
    BITWISEAND #(.width(32)) bitwiseand_1373 (
        .y(_T_2643),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h7F)
    );
    wire _T_2645;
    EQ_UNSIGNED #(.width(32)) u_eq_1374 (
        .y(_T_2645),
        .a(_T_2643),
        .b(32'h6F)
    );
    wire [31:0] _T_2647;
    BITWISEAND #(.width(32)) bitwiseand_1375 (
        .y(_T_2647),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'hFFEFFFFF)
    );
    wire _T_2649;
    EQ_UNSIGNED #(.width(32)) u_eq_1376 (
        .y(_T_2649),
        .a(_T_2647),
        .b(32'h73)
    );
    wire [31:0] _T_2651;
    BITWISEAND #(.width(32)) bitwiseand_1377 (
        .y(_T_2651),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'hFC00305F)
    );
    wire _T_2653;
    EQ_UNSIGNED #(.width(32)) u_eq_1378 (
        .y(_T_2653),
        .a(_T_2651),
        .b(32'h1013)
    );
    wire [31:0] _T_2655;
    BITWISEAND #(.width(32)) bitwiseand_1379 (
        .y(_T_2655),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'hFE00305F)
    );
    wire _T_2657;
    EQ_UNSIGNED #(.width(32)) u_eq_1380 (
        .y(_T_2657),
        .a(_T_2655),
        .b(32'h101B)
    );
    wire [31:0] _T_2659;
    BITWISEAND #(.width(32)) bitwiseand_1381 (
        .y(_T_2659),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h605B)
    );
    wire _T_2661;
    EQ_UNSIGNED #(.width(32)) u_eq_1382 (
        .y(_T_2661),
        .a(_T_2659),
        .b(32'h2003)
    );
    wire [31:0] _T_2663;
    BITWISEAND #(.width(32)) bitwiseand_1383 (
        .y(_T_2663),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h207F)
    );
    wire _T_2665;
    EQ_UNSIGNED #(.width(32)) u_eq_1384 (
        .y(_T_2665),
        .a(_T_2663),
        .b(32'h2013)
    );
    wire [31:0] _T_2667;
    BITWISEAND #(.width(32)) bitwiseand_1385 (
        .y(_T_2667),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h1800607F)
    );
    wire _T_2669;
    EQ_UNSIGNED #(.width(32)) u_eq_1386 (
        .y(_T_2669),
        .a(_T_2667),
        .b(32'h202F)
    );
    wire [31:0] _T_2671;
    BITWISEAND #(.width(32)) bitwiseand_1387 (
        .y(_T_2671),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h207F)
    );
    wire _T_2673;
    EQ_UNSIGNED #(.width(32)) u_eq_1388 (
        .y(_T_2673),
        .a(_T_2671),
        .b(32'h2073)
    );
    wire [31:0] _T_2675;
    BITWISEAND #(.width(32)) bitwiseand_1389 (
        .y(_T_2675),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'hBC00707F)
    );
    wire _T_2677;
    EQ_UNSIGNED #(.width(32)) u_eq_1390 (
        .y(_T_2677),
        .a(_T_2675),
        .b(32'h5013)
    );
    wire [31:0] _T_2679;
    BITWISEAND #(.width(32)) bitwiseand_1391 (
        .y(_T_2679),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'hBE00705F)
    );
    wire _T_2681;
    EQ_UNSIGNED #(.width(32)) u_eq_1392 (
        .y(_T_2681),
        .a(_T_2679),
        .b(32'h501B)
    );
    wire [31:0] _T_2683;
    BITWISEAND #(.width(32)) bitwiseand_1393 (
        .y(_T_2683),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'hBE007077)
    );
    wire _T_2685;
    EQ_UNSIGNED #(.width(32)) u_eq_1394 (
        .y(_T_2685),
        .a(_T_2683),
        .b(32'h5033)
    );
    wire [31:0] _T_2687;
    BITWISEAND #(.width(32)) bitwiseand_1395 (
        .y(_T_2687),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'hFE004077)
    );
    wire _T_2689;
    EQ_UNSIGNED #(.width(32)) u_eq_1396 (
        .y(_T_2689),
        .a(_T_2687),
        .b(32'h2004033)
    );
    wire [31:0] _T_2691;
    BITWISEAND #(.width(32)) bitwiseand_1397 (
        .y(_T_2691),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'hE800607F)
    );
    wire _T_2693;
    EQ_UNSIGNED #(.width(32)) u_eq_1398 (
        .y(_T_2693),
        .a(_T_2691),
        .b(32'h800202F)
    );
    wire [31:0] _T_2695;
    BITWISEAND #(.width(32)) bitwiseand_1399 (
        .y(_T_2695),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'hF9F0607F)
    );
    wire _T_2697;
    EQ_UNSIGNED #(.width(32)) u_eq_1400 (
        .y(_T_2697),
        .a(_T_2695),
        .b(32'h1000202F)
    );
    wire [31:0] _T_2699;
    BITWISEAND #(.width(32)) bitwiseand_1401 (
        .y(_T_2699),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'hDFFFFFFF)
    );
    wire _T_2701;
    EQ_UNSIGNED #(.width(32)) u_eq_1402 (
        .y(_T_2701),
        .a(_T_2699),
        .b(32'h10200073)
    );
    wire _T_2703;
    EQ_UNSIGNED #(.width(32)) u_eq_1403 (
        .y(_T_2703),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h10500073)
    );
    wire [31:0] _T_2705;
    BITWISEAND #(.width(32)) bitwiseand_1404 (
        .y(_T_2705),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'hFE007FFF)
    );
    wire _T_2707;
    EQ_UNSIGNED #(.width(32)) u_eq_1405 (
        .y(_T_2707),
        .a(_T_2705),
        .b(32'h12000073)
    );
    wire [31:0] _T_2709;
    BITWISEAND #(.width(32)) bitwiseand_1406 (
        .y(_T_2709),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'hF400607F)
    );
    wire _T_2711;
    EQ_UNSIGNED #(.width(32)) u_eq_1407 (
        .y(_T_2711),
        .a(_T_2709),
        .b(32'h20000053)
    );
    wire [31:0] _T_2713;
    BITWISEAND #(.width(32)) bitwiseand_1408 (
        .y(_T_2713),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h7C00607F)
    );
    wire _T_2715;
    EQ_UNSIGNED #(.width(32)) u_eq_1409 (
        .y(_T_2715),
        .a(_T_2713),
        .b(32'h20000053)
    );
    wire [31:0] _T_2717;
    BITWISEAND #(.width(32)) bitwiseand_1410 (
        .y(_T_2717),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h7C00507F)
    );
    wire _T_2719;
    EQ_UNSIGNED #(.width(32)) u_eq_1411 (
        .y(_T_2719),
        .a(_T_2717),
        .b(32'h20000053)
    );
    wire [31:0] _T_2721;
    BITWISEAND #(.width(32)) bitwiseand_1412 (
        .y(_T_2721),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h7FF0007F)
    );
    wire _T_2723;
    EQ_UNSIGNED #(.width(32)) u_eq_1413 (
        .y(_T_2723),
        .a(_T_2721),
        .b(32'h40100053)
    );
    wire [31:0] _T_2725;
    BITWISEAND #(.width(32)) bitwiseand_1414 (
        .y(_T_2725),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h7FF0007F)
    );
    wire _T_2727;
    EQ_UNSIGNED #(.width(32)) u_eq_1415 (
        .y(_T_2727),
        .a(_T_2725),
        .b(32'h42000053)
    );
    wire [31:0] _T_2729;
    BITWISEAND #(.width(32)) bitwiseand_1416 (
        .y(_T_2729),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'hFDF0007F)
    );
    wire _T_2731;
    EQ_UNSIGNED #(.width(32)) u_eq_1417 (
        .y(_T_2731),
        .a(_T_2729),
        .b(32'h58000053)
    );
    wire _T_2733;
    EQ_UNSIGNED #(.width(32)) u_eq_1418 (
        .y(_T_2733),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h7B200073)
    );
    wire [31:0] _T_2735;
    BITWISEAND #(.width(32)) bitwiseand_1419 (
        .y(_T_2735),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'hEDC0007F)
    );
    wire _T_2737;
    EQ_UNSIGNED #(.width(32)) u_eq_1420 (
        .y(_T_2737),
        .a(_T_2735),
        .b(32'hC0000053)
    );
    wire [31:0] _T_2739;
    BITWISEAND #(.width(32)) bitwiseand_1421 (
        .y(_T_2739),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'hFDF0607F)
    );
    wire _T_2741;
    EQ_UNSIGNED #(.width(32)) u_eq_1422 (
        .y(_T_2741),
        .a(_T_2739),
        .b(32'hE0000053)
    );
    wire [31:0] _T_2743;
    BITWISEAND #(.width(32)) bitwiseand_1423 (
        .y(_T_2743),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'hEDF0707F)
    );
    wire _T_2745;
    EQ_UNSIGNED #(.width(32)) u_eq_1424 (
        .y(_T_2745),
        .a(_T_2743),
        .b(32'hE0000053)
    );
    wire [31:0] _T_2747;
    BITWISEAND #(.width(32)) bitwiseand_1425 (
        .y(_T_2747),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h603F)
    );
    wire _T_2749;
    EQ_UNSIGNED #(.width(32)) u_eq_1426 (
        .y(_T_2749),
        .a(_T_2747),
        .b(32'h23)
    );
    wire [31:0] _T_2751;
    BITWISEAND #(.width(32)) bitwiseand_1427 (
        .y(_T_2751),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h306F)
    );
    wire _T_2753;
    EQ_UNSIGNED #(.width(32)) u_eq_1428 (
        .y(_T_2753),
        .a(_T_2751),
        .b(32'h1063)
    );
    wire [31:0] _T_2755;
    BITWISEAND #(.width(32)) bitwiseand_1429 (
        .y(_T_2755),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h407F)
    );
    wire _T_2757;
    EQ_UNSIGNED #(.width(32)) u_eq_1430 (
        .y(_T_2757),
        .a(_T_2755),
        .b(32'h4063)
    );
    wire [31:0] _T_2759;
    BITWISEAND #(.width(32)) bitwiseand_1431 (
        .y(_T_2759),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'hFC007077)
    );
    wire _T_2761;
    EQ_UNSIGNED #(.width(32)) u_eq_1432 (
        .y(_T_2761),
        .a(_T_2759),
        .b(32'h33)
    );
    wire _T_2763;
    BITWISEOR #(.width(1)) bitwiseor_1433 (
        .y(_T_2763),
        .a(1'h0),
        .b(_T_2605)
    );
    wire _T_2764;
    BITWISEOR #(.width(1)) bitwiseor_1434 (
        .y(_T_2764),
        .a(_T_2763),
        .b(_T_2609)
    );
    wire _T_2765;
    BITWISEOR #(.width(1)) bitwiseor_1435 (
        .y(_T_2765),
        .a(_T_2764),
        .b(_T_2613)
    );
    wire _T_2766;
    BITWISEOR #(.width(1)) bitwiseor_1436 (
        .y(_T_2766),
        .a(_T_2765),
        .b(_T_2617)
    );
    wire _T_2767;
    BITWISEOR #(.width(1)) bitwiseor_1437 (
        .y(_T_2767),
        .a(_T_2766),
        .b(_T_2621)
    );
    wire _T_2768;
    BITWISEOR #(.width(1)) bitwiseor_1438 (
        .y(_T_2768),
        .a(_T_2767),
        .b(_T_2625)
    );
    wire _T_2769;
    BITWISEOR #(.width(1)) bitwiseor_1439 (
        .y(_T_2769),
        .a(_T_2768),
        .b(_T_2629)
    );
    wire _T_2770;
    BITWISEOR #(.width(1)) bitwiseor_1440 (
        .y(_T_2770),
        .a(_T_2769),
        .b(_T_2633)
    );
    wire _T_2771;
    BITWISEOR #(.width(1)) bitwiseor_1441 (
        .y(_T_2771),
        .a(_T_2770),
        .b(_T_2637)
    );
    wire _T_2772;
    BITWISEOR #(.width(1)) bitwiseor_1442 (
        .y(_T_2772),
        .a(_T_2771),
        .b(_T_2641)
    );
    wire _T_2773;
    BITWISEOR #(.width(1)) bitwiseor_1443 (
        .y(_T_2773),
        .a(_T_2772),
        .b(_T_2645)
    );
    wire _T_2774;
    BITWISEOR #(.width(1)) bitwiseor_1444 (
        .y(_T_2774),
        .a(_T_2773),
        .b(_T_2649)
    );
    wire _T_2775;
    BITWISEOR #(.width(1)) bitwiseor_1445 (
        .y(_T_2775),
        .a(_T_2774),
        .b(_T_2653)
    );
    wire _T_2776;
    BITWISEOR #(.width(1)) bitwiseor_1446 (
        .y(_T_2776),
        .a(_T_2775),
        .b(_T_2657)
    );
    wire _T_2777;
    BITWISEOR #(.width(1)) bitwiseor_1447 (
        .y(_T_2777),
        .a(_T_2776),
        .b(_T_2661)
    );
    wire _T_2778;
    BITWISEOR #(.width(1)) bitwiseor_1448 (
        .y(_T_2778),
        .a(_T_2777),
        .b(_T_2665)
    );
    wire _T_2779;
    BITWISEOR #(.width(1)) bitwiseor_1449 (
        .y(_T_2779),
        .a(_T_2778),
        .b(_T_2669)
    );
    wire _T_2780;
    BITWISEOR #(.width(1)) bitwiseor_1450 (
        .y(_T_2780),
        .a(_T_2779),
        .b(_T_2673)
    );
    wire _T_2781;
    BITWISEOR #(.width(1)) bitwiseor_1451 (
        .y(_T_2781),
        .a(_T_2780),
        .b(_T_2677)
    );
    wire _T_2782;
    BITWISEOR #(.width(1)) bitwiseor_1452 (
        .y(_T_2782),
        .a(_T_2781),
        .b(_T_2681)
    );
    wire _T_2783;
    BITWISEOR #(.width(1)) bitwiseor_1453 (
        .y(_T_2783),
        .a(_T_2782),
        .b(_T_2685)
    );
    wire _T_2784;
    BITWISEOR #(.width(1)) bitwiseor_1454 (
        .y(_T_2784),
        .a(_T_2783),
        .b(_T_2689)
    );
    wire _T_2785;
    BITWISEOR #(.width(1)) bitwiseor_1455 (
        .y(_T_2785),
        .a(_T_2784),
        .b(_T_2693)
    );
    wire _T_2786;
    BITWISEOR #(.width(1)) bitwiseor_1456 (
        .y(_T_2786),
        .a(_T_2785),
        .b(_T_2697)
    );
    wire _T_2787;
    BITWISEOR #(.width(1)) bitwiseor_1457 (
        .y(_T_2787),
        .a(_T_2786),
        .b(_T_2701)
    );
    wire _T_2788;
    BITWISEOR #(.width(1)) bitwiseor_1458 (
        .y(_T_2788),
        .a(_T_2787),
        .b(_T_2703)
    );
    wire _T_2789;
    BITWISEOR #(.width(1)) bitwiseor_1459 (
        .y(_T_2789),
        .a(_T_2788),
        .b(_T_2707)
    );
    wire _T_2790;
    BITWISEOR #(.width(1)) bitwiseor_1460 (
        .y(_T_2790),
        .a(_T_2789),
        .b(_T_2711)
    );
    wire _T_2791;
    BITWISEOR #(.width(1)) bitwiseor_1461 (
        .y(_T_2791),
        .a(_T_2790),
        .b(_T_2715)
    );
    wire _T_2792;
    BITWISEOR #(.width(1)) bitwiseor_1462 (
        .y(_T_2792),
        .a(_T_2791),
        .b(_T_2719)
    );
    wire _T_2793;
    BITWISEOR #(.width(1)) bitwiseor_1463 (
        .y(_T_2793),
        .a(_T_2792),
        .b(_T_2723)
    );
    wire _T_2794;
    BITWISEOR #(.width(1)) bitwiseor_1464 (
        .y(_T_2794),
        .a(_T_2793),
        .b(_T_2727)
    );
    wire _T_2795;
    BITWISEOR #(.width(1)) bitwiseor_1465 (
        .y(_T_2795),
        .a(_T_2794),
        .b(_T_2731)
    );
    wire _T_2796;
    BITWISEOR #(.width(1)) bitwiseor_1466 (
        .y(_T_2796),
        .a(_T_2795),
        .b(_T_2733)
    );
    wire _T_2797;
    BITWISEOR #(.width(1)) bitwiseor_1467 (
        .y(_T_2797),
        .a(_T_2796),
        .b(_T_2737)
    );
    wire _T_2798;
    BITWISEOR #(.width(1)) bitwiseor_1468 (
        .y(_T_2798),
        .a(_T_2797),
        .b(_T_2741)
    );
    wire _T_2799;
    BITWISEOR #(.width(1)) bitwiseor_1469 (
        .y(_T_2799),
        .a(_T_2798),
        .b(_T_2745)
    );
    wire _T_2800;
    BITWISEOR #(.width(1)) bitwiseor_1470 (
        .y(_T_2800),
        .a(_T_2799),
        .b(_T_2749)
    );
    wire _T_2801;
    BITWISEOR #(.width(1)) bitwiseor_1471 (
        .y(_T_2801),
        .a(_T_2800),
        .b(_T_2753)
    );
    wire _T_2802;
    BITWISEOR #(.width(1)) bitwiseor_1472 (
        .y(_T_2802),
        .a(_T_2801),
        .b(_T_2757)
    );
    wire _T_2803;
    BITWISEOR #(.width(1)) bitwiseor_1473 (
        .y(_T_2803),
        .a(_T_2802),
        .b(_T_2761)
    );
    wire [31:0] _T_2805;
    BITWISEAND #(.width(32)) bitwiseand_1474 (
        .y(_T_2805),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h5C)
    );
    wire _T_2807;
    EQ_UNSIGNED #(.width(32)) u_eq_1475 (
        .y(_T_2807),
        .a(_T_2805),
        .b(32'h4)
    );
    wire [31:0] _T_2809;
    BITWISEAND #(.width(32)) bitwiseand_1476 (
        .y(_T_2809),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h60)
    );
    wire _T_2811;
    EQ_UNSIGNED #(.width(32)) u_eq_1477 (
        .y(_T_2811),
        .a(_T_2809),
        .b(32'h40)
    );
    wire _T_2813;
    BITWISEOR #(.width(1)) bitwiseor_1478 (
        .y(_T_2813),
        .a(1'h0),
        .b(_T_2807)
    );
    wire _T_2814;
    BITWISEOR #(.width(1)) bitwiseor_1479 (
        .y(_T_2814),
        .a(_T_2813),
        .b(_T_2811)
    );
    wire [31:0] _T_2817;
    BITWISEAND #(.width(32)) bitwiseand_1480 (
        .y(_T_2817),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h74)
    );
    wire _T_2819;
    EQ_UNSIGNED #(.width(32)) u_eq_1481 (
        .y(_T_2819),
        .a(_T_2817),
        .b(32'h60)
    );
    wire _T_2821;
    BITWISEOR #(.width(1)) bitwiseor_1482 (
        .y(_T_2821),
        .a(1'h0),
        .b(_T_2819)
    );
    wire [31:0] _T_2823;
    BITWISEAND #(.width(32)) bitwiseand_1483 (
        .y(_T_2823),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h68)
    );
    wire _T_2825;
    EQ_UNSIGNED #(.width(32)) u_eq_1484 (
        .y(_T_2825),
        .a(_T_2823),
        .b(32'h68)
    );
    wire _T_2827;
    BITWISEOR #(.width(1)) bitwiseor_1485 (
        .y(_T_2827),
        .a(1'h0),
        .b(_T_2825)
    );
    wire [31:0] _T_2829;
    BITWISEAND #(.width(32)) bitwiseand_1486 (
        .y(_T_2829),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h203C)
    );
    wire _T_2831;
    EQ_UNSIGNED #(.width(32)) u_eq_1487 (
        .y(_T_2831),
        .a(_T_2829),
        .b(32'h24)
    );
    wire _T_2833;
    BITWISEOR #(.width(1)) bitwiseor_1488 (
        .y(_T_2833),
        .a(1'h0),
        .b(_T_2831)
    );
    wire [31:0] _T_2835;
    BITWISEAND #(.width(32)) bitwiseand_1489 (
        .y(_T_2835),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h64)
    );
    wire _T_2837;
    EQ_UNSIGNED #(.width(32)) u_eq_1490 (
        .y(_T_2837),
        .a(_T_2835),
        .b(32'h20)
    );
    wire [31:0] _T_2839;
    BITWISEAND #(.width(32)) bitwiseand_1491 (
        .y(_T_2839),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h34)
    );
    wire _T_2841;
    EQ_UNSIGNED #(.width(32)) u_eq_1492 (
        .y(_T_2841),
        .a(_T_2839),
        .b(32'h20)
    );
    wire [31:0] _T_2843;
    BITWISEAND #(.width(32)) bitwiseand_1493 (
        .y(_T_2843),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h2048)
    );
    wire _T_2845;
    EQ_UNSIGNED #(.width(32)) u_eq_1494 (
        .y(_T_2845),
        .a(_T_2843),
        .b(32'h2008)
    );
    wire [31:0] _T_2847;
    BITWISEAND #(.width(32)) bitwiseand_1495 (
        .y(_T_2847),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h42003024)
    );
    wire _T_2849;
    EQ_UNSIGNED #(.width(32)) u_eq_1496 (
        .y(_T_2849),
        .a(_T_2847),
        .b(32'h2000020)
    );
    wire _T_2851;
    BITWISEOR #(.width(1)) bitwiseor_1497 (
        .y(_T_2851),
        .a(1'h0),
        .b(_T_2837)
    );
    wire _T_2852;
    BITWISEOR #(.width(1)) bitwiseor_1498 (
        .y(_T_2852),
        .a(_T_2851),
        .b(_T_2841)
    );
    wire _T_2853;
    BITWISEOR #(.width(1)) bitwiseor_1499 (
        .y(_T_2853),
        .a(_T_2852),
        .b(_T_2845)
    );
    wire _T_2854;
    BITWISEOR #(.width(1)) bitwiseor_1500 (
        .y(_T_2854),
        .a(_T_2853),
        .b(_T_2849)
    );
    wire [31:0] _T_2856;
    BITWISEAND #(.width(32)) bitwiseand_1501 (
        .y(_T_2856),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h44)
    );
    wire _T_2858;
    EQ_UNSIGNED #(.width(32)) u_eq_1502 (
        .y(_T_2858),
        .a(_T_2856),
        .b(32'h0)
    );
    wire [31:0] _T_2860;
    BITWISEAND #(.width(32)) bitwiseand_1503 (
        .y(_T_2860),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h4024)
    );
    wire _T_2862;
    EQ_UNSIGNED #(.width(32)) u_eq_1504 (
        .y(_T_2862),
        .a(_T_2860),
        .b(32'h20)
    );
    wire [31:0] _T_2864;
    BITWISEAND #(.width(32)) bitwiseand_1505 (
        .y(_T_2864),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h38)
    );
    wire _T_2866;
    EQ_UNSIGNED #(.width(32)) u_eq_1506 (
        .y(_T_2866),
        .a(_T_2864),
        .b(32'h20)
    );
    wire [31:0] _T_2868;
    BITWISEAND #(.width(32)) bitwiseand_1507 (
        .y(_T_2868),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h2050)
    );
    wire _T_2870;
    EQ_UNSIGNED #(.width(32)) u_eq_1508 (
        .y(_T_2870),
        .a(_T_2868),
        .b(32'h2000)
    );
    wire [31:0] _T_2872;
    BITWISEAND #(.width(32)) bitwiseand_1509 (
        .y(_T_2872),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h90000034)
    );
    wire _T_2874;
    EQ_UNSIGNED #(.width(32)) u_eq_1510 (
        .y(_T_2874),
        .a(_T_2872),
        .b(32'h90000010)
    );
    wire _T_2876;
    BITWISEOR #(.width(1)) bitwiseor_1511 (
        .y(_T_2876),
        .a(1'h0),
        .b(_T_2858)
    );
    wire _T_2877;
    BITWISEOR #(.width(1)) bitwiseor_1512 (
        .y(_T_2877),
        .a(_T_2876),
        .b(_T_2862)
    );
    wire _T_2878;
    BITWISEOR #(.width(1)) bitwiseor_1513 (
        .y(_T_2878),
        .a(_T_2877),
        .b(_T_2866)
    );
    wire _T_2879;
    BITWISEOR #(.width(1)) bitwiseor_1514 (
        .y(_T_2879),
        .a(_T_2878),
        .b(_T_2870)
    );
    wire _T_2880;
    BITWISEOR #(.width(1)) bitwiseor_1515 (
        .y(_T_2880),
        .a(_T_2879),
        .b(_T_2874)
    );
    wire [31:0] _T_2882;
    BITWISEAND #(.width(32)) bitwiseand_1516 (
        .y(_T_2882),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h58)
    );
    wire _T_2884;
    EQ_UNSIGNED #(.width(32)) u_eq_1517 (
        .y(_T_2884),
        .a(_T_2882),
        .b(32'h0)
    );
    wire [31:0] _T_2886;
    BITWISEAND #(.width(32)) bitwiseand_1518 (
        .y(_T_2886),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h20)
    );
    wire _T_2888;
    EQ_UNSIGNED #(.width(32)) u_eq_1519 (
        .y(_T_2888),
        .a(_T_2886),
        .b(32'h0)
    );
    wire [31:0] _T_2890;
    BITWISEAND #(.width(32)) bitwiseand_1520 (
        .y(_T_2890),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'hC)
    );
    wire _T_2892;
    EQ_UNSIGNED #(.width(32)) u_eq_1521 (
        .y(_T_2892),
        .a(_T_2890),
        .b(32'h4)
    );
    wire [31:0] _T_2894;
    BITWISEAND #(.width(32)) bitwiseand_1522 (
        .y(_T_2894),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h48)
    );
    wire _T_2896;
    EQ_UNSIGNED #(.width(32)) u_eq_1523 (
        .y(_T_2896),
        .a(_T_2894),
        .b(32'h48)
    );
    wire [31:0] _T_2898;
    BITWISEAND #(.width(32)) bitwiseand_1524 (
        .y(_T_2898),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h4050)
    );
    wire _T_2900;
    EQ_UNSIGNED #(.width(32)) u_eq_1525 (
        .y(_T_2900),
        .a(_T_2898),
        .b(32'h4050)
    );
    wire _T_2902;
    BITWISEOR #(.width(1)) bitwiseor_1526 (
        .y(_T_2902),
        .a(1'h0),
        .b(_T_2884)
    );
    wire _T_2903;
    BITWISEOR #(.width(1)) bitwiseor_1527 (
        .y(_T_2903),
        .a(_T_2902),
        .b(_T_2888)
    );
    wire _T_2904;
    BITWISEOR #(.width(1)) bitwiseor_1528 (
        .y(_T_2904),
        .a(_T_2903),
        .b(_T_2892)
    );
    wire _T_2905;
    BITWISEOR #(.width(1)) bitwiseor_1529 (
        .y(_T_2905),
        .a(_T_2904),
        .b(_T_2896)
    );
    wire _T_2906;
    BITWISEOR #(.width(1)) bitwiseor_1530 (
        .y(_T_2906),
        .a(_T_2905),
        .b(_T_2900)
    );
    wire [31:0] _T_2908;
    BITWISEAND #(.width(32)) bitwiseand_1531 (
        .y(_T_2908),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h48)
    );
    wire _T_2910;
    EQ_UNSIGNED #(.width(32)) u_eq_1532 (
        .y(_T_2910),
        .a(_T_2908),
        .b(32'h0)
    );
    wire [31:0] _T_2912;
    BITWISEAND #(.width(32)) bitwiseand_1533 (
        .y(_T_2912),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h18)
    );
    wire _T_2914;
    EQ_UNSIGNED #(.width(32)) u_eq_1534 (
        .y(_T_2914),
        .a(_T_2912),
        .b(32'h0)
    );
    wire [31:0] _T_2916;
    BITWISEAND #(.width(32)) bitwiseand_1535 (
        .y(_T_2916),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h4008)
    );
    wire _T_2918;
    EQ_UNSIGNED #(.width(32)) u_eq_1536 (
        .y(_T_2918),
        .a(_T_2916),
        .b(32'h4000)
    );
    wire _T_2920;
    BITWISEOR #(.width(1)) bitwiseor_1537 (
        .y(_T_2920),
        .a(1'h0),
        .b(_T_2910)
    );
    wire _T_2921;
    BITWISEOR #(.width(1)) bitwiseor_1538 (
        .y(_T_2921),
        .a(_T_2920),
        .b(_T_2858)
    );
    wire _T_2922;
    BITWISEOR #(.width(1)) bitwiseor_1539 (
        .y(_T_2922),
        .a(_T_2921),
        .b(_T_2914)
    );
    wire _T_2923;
    BITWISEOR #(.width(1)) bitwiseor_1540 (
        .y(_T_2923),
        .a(_T_2922),
        .b(_T_2918)
    );
    wire [1:0] _T_2924;
    CAT #(.width_a(1), .width_b(1)) cat_1541 (
        .y(_T_2924),
        .a(_T_2923),
        .b(_T_2906)
    );
    wire [31:0] _T_2926;
    BITWISEAND #(.width(32)) bitwiseand_1542 (
        .y(_T_2926),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h4004)
    );
    wire _T_2928;
    EQ_UNSIGNED #(.width(32)) u_eq_1543 (
        .y(_T_2928),
        .a(_T_2926),
        .b(32'h0)
    );
    wire [31:0] _T_2930;
    BITWISEAND #(.width(32)) bitwiseand_1544 (
        .y(_T_2930),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h50)
    );
    wire _T_2932;
    EQ_UNSIGNED #(.width(32)) u_eq_1545 (
        .y(_T_2932),
        .a(_T_2930),
        .b(32'h0)
    );
    wire [31:0] _T_2934;
    BITWISEAND #(.width(32)) bitwiseand_1546 (
        .y(_T_2934),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h24)
    );
    wire _T_2936;
    EQ_UNSIGNED #(.width(32)) u_eq_1547 (
        .y(_T_2936),
        .a(_T_2934),
        .b(32'h0)
    );
    wire _T_2938;
    BITWISEOR #(.width(1)) bitwiseor_1548 (
        .y(_T_2938),
        .a(1'h0),
        .b(_T_2928)
    );
    wire _T_2939;
    BITWISEOR #(.width(1)) bitwiseor_1549 (
        .y(_T_2939),
        .a(_T_2938),
        .b(_T_2932)
    );
    wire _T_2940;
    BITWISEOR #(.width(1)) bitwiseor_1550 (
        .y(_T_2940),
        .a(_T_2939),
        .b(_T_2858)
    );
    wire _T_2941;
    BITWISEOR #(.width(1)) bitwiseor_1551 (
        .y(_T_2941),
        .a(_T_2940),
        .b(_T_2936)
    );
    wire _T_2942;
    BITWISEOR #(.width(1)) bitwiseor_1552 (
        .y(_T_2942),
        .a(_T_2941),
        .b(_T_2914)
    );
    wire [31:0] _T_2944;
    BITWISEAND #(.width(32)) bitwiseand_1553 (
        .y(_T_2944),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h34)
    );
    wire _T_2946;
    EQ_UNSIGNED #(.width(32)) u_eq_1554 (
        .y(_T_2946),
        .a(_T_2944),
        .b(32'h14)
    );
    wire _T_2948;
    BITWISEOR #(.width(1)) bitwiseor_1555 (
        .y(_T_2948),
        .a(1'h0),
        .b(_T_2946)
    );
    wire _T_2949;
    BITWISEOR #(.width(1)) bitwiseor_1556 (
        .y(_T_2949),
        .a(_T_2948),
        .b(_T_2896)
    );
    wire [1:0] _T_2950;
    CAT #(.width_a(1), .width_b(1)) cat_1557 (
        .y(_T_2950),
        .a(_T_2949),
        .b(_T_2942)
    );
    wire [31:0] _T_2952;
    BITWISEAND #(.width(32)) bitwiseand_1558 (
        .y(_T_2952),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h18)
    );
    wire _T_2954;
    EQ_UNSIGNED #(.width(32)) u_eq_1559 (
        .y(_T_2954),
        .a(_T_2952),
        .b(32'h8)
    );
    wire [31:0] _T_2956;
    BITWISEAND #(.width(32)) bitwiseand_1560 (
        .y(_T_2956),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h44)
    );
    wire _T_2958;
    EQ_UNSIGNED #(.width(32)) u_eq_1561 (
        .y(_T_2958),
        .a(_T_2956),
        .b(32'h40)
    );
    wire _T_2960;
    BITWISEOR #(.width(1)) bitwiseor_1562 (
        .y(_T_2960),
        .a(1'h0),
        .b(_T_2954)
    );
    wire _T_2961;
    BITWISEOR #(.width(1)) bitwiseor_1563 (
        .y(_T_2961),
        .a(_T_2960),
        .b(_T_2958)
    );
    wire [31:0] _T_2963;
    BITWISEAND #(.width(32)) bitwiseand_1564 (
        .y(_T_2963),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h14)
    );
    wire _T_2965;
    EQ_UNSIGNED #(.width(32)) u_eq_1565 (
        .y(_T_2965),
        .a(_T_2963),
        .b(32'h14)
    );
    wire _T_2967;
    BITWISEOR #(.width(1)) bitwiseor_1566 (
        .y(_T_2967),
        .a(1'h0),
        .b(_T_2954)
    );
    wire _T_2968;
    BITWISEOR #(.width(1)) bitwiseor_1567 (
        .y(_T_2968),
        .a(_T_2967),
        .b(_T_2965)
    );
    wire [31:0] _T_2970;
    BITWISEAND #(.width(32)) bitwiseand_1568 (
        .y(_T_2970),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h30)
    );
    wire _T_2972;
    EQ_UNSIGNED #(.width(32)) u_eq_1569 (
        .y(_T_2972),
        .a(_T_2970),
        .b(32'h0)
    );
    wire [31:0] _T_2974;
    BITWISEAND #(.width(32)) bitwiseand_1570 (
        .y(_T_2974),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h201C)
    );
    wire _T_2976;
    EQ_UNSIGNED #(.width(32)) u_eq_1571 (
        .y(_T_2976),
        .a(_T_2974),
        .b(32'h4)
    );
    wire [31:0] _T_2978;
    BITWISEAND #(.width(32)) bitwiseand_1572 (
        .y(_T_2978),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h14)
    );
    wire _T_2980;
    EQ_UNSIGNED #(.width(32)) u_eq_1573 (
        .y(_T_2980),
        .a(_T_2978),
        .b(32'h10)
    );
    wire _T_2982;
    BITWISEOR #(.width(1)) bitwiseor_1574 (
        .y(_T_2982),
        .a(1'h0),
        .b(_T_2972)
    );
    wire _T_2983;
    BITWISEOR #(.width(1)) bitwiseor_1575 (
        .y(_T_2983),
        .a(_T_2982),
        .b(_T_2976)
    );
    wire _T_2984;
    BITWISEOR #(.width(1)) bitwiseor_1576 (
        .y(_T_2984),
        .a(_T_2983),
        .b(_T_2980)
    );
    wire [1:0] _T_2985;
    CAT #(.width_a(1), .width_b(1)) cat_1577 (
        .y(_T_2985),
        .a(_T_2984),
        .b(_T_2968)
    );
    wire [2:0] _T_2986;
    CAT #(.width_a(2), .width_b(1)) cat_1578 (
        .y(_T_2986),
        .a(_T_2985),
        .b(_T_2961)
    );
    wire [31:0] _T_2988;
    BITWISEAND #(.width(32)) bitwiseand_1579 (
        .y(_T_2988),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h10)
    );
    wire _T_2990;
    EQ_UNSIGNED #(.width(32)) u_eq_1580 (
        .y(_T_2990),
        .a(_T_2988),
        .b(32'h0)
    );
    wire [31:0] _T_2992;
    BITWISEAND #(.width(32)) bitwiseand_1581 (
        .y(_T_2992),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h8)
    );
    wire _T_2994;
    EQ_UNSIGNED #(.width(32)) u_eq_1582 (
        .y(_T_2994),
        .a(_T_2992),
        .b(32'h0)
    );
    wire _T_2996;
    BITWISEOR #(.width(1)) bitwiseor_1583 (
        .y(_T_2996),
        .a(1'h0),
        .b(_T_2990)
    );
    wire _T_2997;
    BITWISEOR #(.width(1)) bitwiseor_1584 (
        .y(_T_2997),
        .a(_T_2996),
        .b(_T_2994)
    );
    wire [31:0] _T_2999;
    BITWISEAND #(.width(32)) bitwiseand_1585 (
        .y(_T_2999),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h3054)
    );
    wire _T_3001;
    EQ_UNSIGNED #(.width(32)) u_eq_1586 (
        .y(_T_3001),
        .a(_T_2999),
        .b(32'h1010)
    );
    wire [31:0] _T_3003;
    BITWISEAND #(.width(32)) bitwiseand_1587 (
        .y(_T_3003),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h1058)
    );
    wire _T_3005;
    EQ_UNSIGNED #(.width(32)) u_eq_1588 (
        .y(_T_3005),
        .a(_T_3003),
        .b(32'h1040)
    );
    wire [31:0] _T_3007;
    BITWISEAND #(.width(32)) bitwiseand_1589 (
        .y(_T_3007),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h7044)
    );
    wire _T_3009;
    EQ_UNSIGNED #(.width(32)) u_eq_1590 (
        .y(_T_3009),
        .a(_T_3007),
        .b(32'h7000)
    );
    wire _T_3011;
    BITWISEOR #(.width(1)) bitwiseor_1591 (
        .y(_T_3011),
        .a(1'h0),
        .b(_T_3001)
    );
    wire _T_3012;
    BITWISEOR #(.width(1)) bitwiseor_1592 (
        .y(_T_3012),
        .a(_T_3011),
        .b(_T_3005)
    );
    wire _T_3013;
    BITWISEOR #(.width(1)) bitwiseor_1593 (
        .y(_T_3013),
        .a(_T_3012),
        .b(_T_3009)
    );
    wire [31:0] _T_3015;
    BITWISEAND #(.width(32)) bitwiseand_1594 (
        .y(_T_3015),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h4054)
    );
    wire _T_3017;
    EQ_UNSIGNED #(.width(32)) u_eq_1595 (
        .y(_T_3017),
        .a(_T_3015),
        .b(32'h40)
    );
    wire [31:0] _T_3019;
    BITWISEAND #(.width(32)) bitwiseand_1596 (
        .y(_T_3019),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h2058)
    );
    wire _T_3021;
    EQ_UNSIGNED #(.width(32)) u_eq_1597 (
        .y(_T_3021),
        .a(_T_3019),
        .b(32'h2040)
    );
    wire [31:0] _T_3023;
    BITWISEAND #(.width(32)) bitwiseand_1598 (
        .y(_T_3023),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h3054)
    );
    wire _T_3025;
    EQ_UNSIGNED #(.width(32)) u_eq_1599 (
        .y(_T_3025),
        .a(_T_3023),
        .b(32'h3010)
    );
    wire [31:0] _T_3027;
    BITWISEAND #(.width(32)) bitwiseand_1600 (
        .y(_T_3027),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h6054)
    );
    wire _T_3029;
    EQ_UNSIGNED #(.width(32)) u_eq_1601 (
        .y(_T_3029),
        .a(_T_3027),
        .b(32'h6010)
    );
    wire [31:0] _T_3031;
    BITWISEAND #(.width(32)) bitwiseand_1602 (
        .y(_T_3031),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h40003034)
    );
    wire _T_3033;
    EQ_UNSIGNED #(.width(32)) u_eq_1603 (
        .y(_T_3033),
        .a(_T_3031),
        .b(32'h40000030)
    );
    wire [31:0] _T_3035;
    BITWISEAND #(.width(32)) bitwiseand_1604 (
        .y(_T_3035),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h40001054)
    );
    wire _T_3037;
    EQ_UNSIGNED #(.width(32)) u_eq_1605 (
        .y(_T_3037),
        .a(_T_3035),
        .b(32'h40001010)
    );
    wire _T_3039;
    BITWISEOR #(.width(1)) bitwiseor_1606 (
        .y(_T_3039),
        .a(1'h0),
        .b(_T_3017)
    );
    wire _T_3040;
    BITWISEOR #(.width(1)) bitwiseor_1607 (
        .y(_T_3040),
        .a(_T_3039),
        .b(_T_3021)
    );
    wire _T_3041;
    BITWISEOR #(.width(1)) bitwiseor_1608 (
        .y(_T_3041),
        .a(_T_3040),
        .b(_T_3025)
    );
    wire _T_3042;
    BITWISEOR #(.width(1)) bitwiseor_1609 (
        .y(_T_3042),
        .a(_T_3041),
        .b(_T_3029)
    );
    wire _T_3043;
    BITWISEOR #(.width(1)) bitwiseor_1610 (
        .y(_T_3043),
        .a(_T_3042),
        .b(_T_3033)
    );
    wire _T_3044;
    BITWISEOR #(.width(1)) bitwiseor_1611 (
        .y(_T_3044),
        .a(_T_3043),
        .b(_T_3037)
    );
    wire [31:0] _T_3046;
    BITWISEAND #(.width(32)) bitwiseand_1612 (
        .y(_T_3046),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h2054)
    );
    wire _T_3048;
    EQ_UNSIGNED #(.width(32)) u_eq_1613 (
        .y(_T_3048),
        .a(_T_3046),
        .b(32'h2010)
    );
    wire [31:0] _T_3050;
    BITWISEAND #(.width(32)) bitwiseand_1614 (
        .y(_T_3050),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h40004054)
    );
    wire _T_3052;
    EQ_UNSIGNED #(.width(32)) u_eq_1615 (
        .y(_T_3052),
        .a(_T_3050),
        .b(32'h4010)
    );
    wire [31:0] _T_3054;
    BITWISEAND #(.width(32)) bitwiseand_1616 (
        .y(_T_3054),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h5054)
    );
    wire _T_3056;
    EQ_UNSIGNED #(.width(32)) u_eq_1617 (
        .y(_T_3056),
        .a(_T_3054),
        .b(32'h4010)
    );
    wire [31:0] _T_3058;
    BITWISEAND #(.width(32)) bitwiseand_1618 (
        .y(_T_3058),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h4058)
    );
    wire _T_3060;
    EQ_UNSIGNED #(.width(32)) u_eq_1619 (
        .y(_T_3060),
        .a(_T_3058),
        .b(32'h4040)
    );
    wire _T_3062;
    BITWISEOR #(.width(1)) bitwiseor_1620 (
        .y(_T_3062),
        .a(1'h0),
        .b(_T_3048)
    );
    wire _T_3063;
    BITWISEOR #(.width(1)) bitwiseor_1621 (
        .y(_T_3063),
        .a(_T_3062),
        .b(_T_3052)
    );
    wire _T_3064;
    BITWISEOR #(.width(1)) bitwiseor_1622 (
        .y(_T_3064),
        .a(_T_3063),
        .b(_T_3056)
    );
    wire _T_3065;
    BITWISEOR #(.width(1)) bitwiseor_1623 (
        .y(_T_3065),
        .a(_T_3064),
        .b(_T_3060)
    );
    wire [31:0] _T_3067;
    BITWISEAND #(.width(32)) bitwiseand_1624 (
        .y(_T_3067),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h6054)
    );
    wire _T_3069;
    EQ_UNSIGNED #(.width(32)) u_eq_1625 (
        .y(_T_3069),
        .a(_T_3067),
        .b(32'h2010)
    );
    wire [31:0] _T_3071;
    BITWISEAND #(.width(32)) bitwiseand_1626 (
        .y(_T_3071),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h40003054)
    );
    wire _T_3073;
    EQ_UNSIGNED #(.width(32)) u_eq_1627 (
        .y(_T_3073),
        .a(_T_3071),
        .b(32'h40001010)
    );
    wire _T_3075;
    BITWISEOR #(.width(1)) bitwiseor_1628 (
        .y(_T_3075),
        .a(1'h0),
        .b(_T_3069)
    );
    wire _T_3076;
    BITWISEOR #(.width(1)) bitwiseor_1629 (
        .y(_T_3076),
        .a(_T_3075),
        .b(_T_3060)
    );
    wire _T_3077;
    BITWISEOR #(.width(1)) bitwiseor_1630 (
        .y(_T_3077),
        .a(_T_3076),
        .b(_T_3033)
    );
    wire _T_3078;
    BITWISEOR #(.width(1)) bitwiseor_1631 (
        .y(_T_3078),
        .a(_T_3077),
        .b(_T_3073)
    );
    wire [1:0] _T_3079;
    CAT #(.width_a(1), .width_b(1)) cat_1632 (
        .y(_T_3079),
        .a(_T_3044),
        .b(_T_3013)
    );
    wire [1:0] _T_3080;
    CAT #(.width_a(1), .width_b(1)) cat_1633 (
        .y(_T_3080),
        .a(_T_3078),
        .b(_T_3065)
    );
    wire [3:0] _T_3081;
    CAT #(.width_a(2), .width_b(2)) cat_1634 (
        .y(_T_3081),
        .a(_T_3080),
        .b(_T_3079)
    );
    wire [31:0] _T_3083;
    BITWISEAND #(.width(32)) bitwiseand_1635 (
        .y(_T_3083),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h405F)
    );
    wire _T_3085;
    EQ_UNSIGNED #(.width(32)) u_eq_1636 (
        .y(_T_3085),
        .a(_T_3083),
        .b(32'h3)
    );
    wire [31:0] _T_3087;
    BITWISEAND #(.width(32)) bitwiseand_1637 (
        .y(_T_3087),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h107F)
    );
    wire _T_3089;
    EQ_UNSIGNED #(.width(32)) u_eq_1638 (
        .y(_T_3089),
        .a(_T_3087),
        .b(32'h3)
    );
    wire [31:0] _T_3091;
    BITWISEAND #(.width(32)) bitwiseand_1639 (
        .y(_T_3091),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h707F)
    );
    wire _T_3093;
    EQ_UNSIGNED #(.width(32)) u_eq_1640 (
        .y(_T_3093),
        .a(_T_3091),
        .b(32'h100F)
    );
    wire _T_3095;
    BITWISEOR #(.width(1)) bitwiseor_1641 (
        .y(_T_3095),
        .a(1'h0),
        .b(_T_3085)
    );
    wire _T_3096;
    BITWISEOR #(.width(1)) bitwiseor_1642 (
        .y(_T_3096),
        .a(_T_3095),
        .b(_T_2605)
    );
    wire _T_3097;
    BITWISEOR #(.width(1)) bitwiseor_1643 (
        .y(_T_3097),
        .a(_T_3096),
        .b(_T_3089)
    );
    wire _T_3098;
    BITWISEOR #(.width(1)) bitwiseor_1644 (
        .y(_T_3098),
        .a(_T_3097),
        .b(_T_3093)
    );
    wire _T_3099;
    BITWISEOR #(.width(1)) bitwiseor_1645 (
        .y(_T_3099),
        .a(_T_3098),
        .b(_T_2661)
    );
    wire _T_3100;
    BITWISEOR #(.width(1)) bitwiseor_1646 (
        .y(_T_3100),
        .a(_T_3099),
        .b(_T_2669)
    );
    wire _T_3101;
    BITWISEOR #(.width(1)) bitwiseor_1647 (
        .y(_T_3101),
        .a(_T_3100),
        .b(_T_2693)
    );
    wire _T_3102;
    BITWISEOR #(.width(1)) bitwiseor_1648 (
        .y(_T_3102),
        .a(_T_3101),
        .b(_T_2697)
    );
    wire [31:0] _T_3104;
    BITWISEAND #(.width(32)) bitwiseand_1649 (
        .y(_T_3104),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h2008)
    );
    wire _T_3106;
    EQ_UNSIGNED #(.width(32)) u_eq_1650 (
        .y(_T_3106),
        .a(_T_3104),
        .b(32'h8)
    );
    wire [31:0] _T_3108;
    BITWISEAND #(.width(32)) bitwiseand_1651 (
        .y(_T_3108),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h28)
    );
    wire _T_3110;
    EQ_UNSIGNED #(.width(32)) u_eq_1652 (
        .y(_T_3110),
        .a(_T_3108),
        .b(32'h20)
    );
    wire [31:0] _T_3112;
    BITWISEAND #(.width(32)) bitwiseand_1653 (
        .y(_T_3112),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h18000020)
    );
    wire _T_3114;
    EQ_UNSIGNED #(.width(32)) u_eq_1654 (
        .y(_T_3114),
        .a(_T_3112),
        .b(32'h18000020)
    );
    wire [31:0] _T_3116;
    BITWISEAND #(.width(32)) bitwiseand_1655 (
        .y(_T_3116),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h20000020)
    );
    wire _T_3118;
    EQ_UNSIGNED #(.width(32)) u_eq_1656 (
        .y(_T_3118),
        .a(_T_3116),
        .b(32'h20000020)
    );
    wire _T_3120;
    BITWISEOR #(.width(1)) bitwiseor_1657 (
        .y(_T_3120),
        .a(1'h0),
        .b(_T_3106)
    );
    wire _T_3121;
    BITWISEOR #(.width(1)) bitwiseor_1658 (
        .y(_T_3121),
        .a(_T_3120),
        .b(_T_3110)
    );
    wire _T_3122;
    BITWISEOR #(.width(1)) bitwiseor_1659 (
        .y(_T_3122),
        .a(_T_3121),
        .b(_T_3114)
    );
    wire _T_3123;
    BITWISEOR #(.width(1)) bitwiseor_1660 (
        .y(_T_3123),
        .a(_T_3122),
        .b(_T_3118)
    );
    wire [31:0] _T_3125;
    BITWISEAND #(.width(32)) bitwiseand_1661 (
        .y(_T_3125),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h10002008)
    );
    wire _T_3127;
    EQ_UNSIGNED #(.width(32)) u_eq_1662 (
        .y(_T_3127),
        .a(_T_3125),
        .b(32'h10002008)
    );
    wire [31:0] _T_3129;
    BITWISEAND #(.width(32)) bitwiseand_1663 (
        .y(_T_3129),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h40002008)
    );
    wire _T_3131;
    EQ_UNSIGNED #(.width(32)) u_eq_1664 (
        .y(_T_3131),
        .a(_T_3129),
        .b(32'h40002008)
    );
    wire _T_3133;
    BITWISEOR #(.width(1)) bitwiseor_1665 (
        .y(_T_3133),
        .a(1'h0),
        .b(_T_3127)
    );
    wire _T_3134;
    BITWISEOR #(.width(1)) bitwiseor_1666 (
        .y(_T_3134),
        .a(_T_3133),
        .b(_T_3131)
    );
    wire [31:0] _T_3136;
    BITWISEAND #(.width(32)) bitwiseand_1667 (
        .y(_T_3136),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h8000008)
    );
    wire _T_3138;
    EQ_UNSIGNED #(.width(32)) u_eq_1668 (
        .y(_T_3138),
        .a(_T_3136),
        .b(32'h8000008)
    );
    wire [31:0] _T_3140;
    BITWISEAND #(.width(32)) bitwiseand_1669 (
        .y(_T_3140),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h10000008)
    );
    wire _T_3142;
    EQ_UNSIGNED #(.width(32)) u_eq_1670 (
        .y(_T_3142),
        .a(_T_3140),
        .b(32'h10000008)
    );
    wire [31:0] _T_3144;
    BITWISEAND #(.width(32)) bitwiseand_1671 (
        .y(_T_3144),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h80000008)
    );
    wire _T_3146;
    EQ_UNSIGNED #(.width(32)) u_eq_1672 (
        .y(_T_3146),
        .a(_T_3144),
        .b(32'h80000008)
    );
    wire _T_3148;
    BITWISEOR #(.width(1)) bitwiseor_1673 (
        .y(_T_3148),
        .a(1'h0),
        .b(_T_3106)
    );
    wire _T_3149;
    BITWISEOR #(.width(1)) bitwiseor_1674 (
        .y(_T_3149),
        .a(_T_3148),
        .b(_T_3138)
    );
    wire _T_3150;
    BITWISEOR #(.width(1)) bitwiseor_1675 (
        .y(_T_3150),
        .a(_T_3149),
        .b(_T_3142)
    );
    wire _T_3151;
    BITWISEOR #(.width(1)) bitwiseor_1676 (
        .y(_T_3151),
        .a(_T_3150),
        .b(_T_3146)
    );
    wire [31:0] _T_3153;
    BITWISEAND #(.width(32)) bitwiseand_1677 (
        .y(_T_3153),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h18002008)
    );
    wire _T_3155;
    EQ_UNSIGNED #(.width(32)) u_eq_1678 (
        .y(_T_3155),
        .a(_T_3153),
        .b(32'h2008)
    );
    wire _T_3157;
    BITWISEOR #(.width(1)) bitwiseor_1679 (
        .y(_T_3157),
        .a(1'h0),
        .b(_T_3155)
    );
    wire [1:0] _T_3159;
    CAT #(.width_a(1), .width_b(1)) cat_1680 (
        .y(_T_3159),
        .a(_T_3134),
        .b(_T_3123)
    );
    wire [1:0] _T_3160;
    CAT #(.width_a(1), .width_b(1)) cat_1681 (
        .y(_T_3160),
        .a(1'h0),
        .b(_T_3157)
    );
    wire [2:0] _T_3161;
    CAT #(.width_a(2), .width_b(1)) cat_1682 (
        .y(_T_3161),
        .a(_T_3160),
        .b(_T_3151)
    );
    wire [4:0] _T_3162;
    CAT #(.width_a(3), .width_b(2)) cat_1683 (
        .y(_T_3162),
        .a(_T_3161),
        .b(_T_3159)
    );
    wire [31:0] _T_3164;
    BITWISEAND #(.width(32)) bitwiseand_1684 (
        .y(_T_3164),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h1000)
    );
    wire _T_3166;
    EQ_UNSIGNED #(.width(32)) u_eq_1685 (
        .y(_T_3166),
        .a(_T_3164),
        .b(32'h1000)
    );
    wire _T_3168;
    BITWISEOR #(.width(1)) bitwiseor_1686 (
        .y(_T_3168),
        .a(1'h0),
        .b(_T_3166)
    );
    wire [31:0] _T_3170;
    BITWISEAND #(.width(32)) bitwiseand_1687 (
        .y(_T_3170),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h2000)
    );
    wire _T_3172;
    EQ_UNSIGNED #(.width(32)) u_eq_1688 (
        .y(_T_3172),
        .a(_T_3170),
        .b(32'h2000)
    );
    wire _T_3174;
    BITWISEOR #(.width(1)) bitwiseor_1689 (
        .y(_T_3174),
        .a(1'h0),
        .b(_T_3172)
    );
    wire [31:0] _T_3176;
    BITWISEAND #(.width(32)) bitwiseand_1690 (
        .y(_T_3176),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h4000)
    );
    wire _T_3178;
    EQ_UNSIGNED #(.width(32)) u_eq_1691 (
        .y(_T_3178),
        .a(_T_3176),
        .b(32'h4000)
    );
    wire _T_3180;
    BITWISEOR #(.width(1)) bitwiseor_1692 (
        .y(_T_3180),
        .a(1'h0),
        .b(_T_3178)
    );
    wire [1:0] _T_3181;
    CAT #(.width_a(1), .width_b(1)) cat_1693 (
        .y(_T_3181),
        .a(_T_3180),
        .b(_T_3174)
    );
    wire [2:0] _T_3182;
    CAT #(.width_a(2), .width_b(1)) cat_1694 (
        .y(_T_3182),
        .a(_T_3181),
        .b(_T_3168)
    );
    wire [31:0] _T_3184;
    BITWISEAND #(.width(32)) bitwiseand_1695 (
        .y(_T_3184),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h80000060)
    );
    wire _T_3186;
    EQ_UNSIGNED #(.width(32)) u_eq_1696 (
        .y(_T_3186),
        .a(_T_3184),
        .b(32'h40)
    );
    wire [31:0] _T_3188;
    BITWISEAND #(.width(32)) bitwiseand_1697 (
        .y(_T_3188),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h10000060)
    );
    wire _T_3190;
    EQ_UNSIGNED #(.width(32)) u_eq_1698 (
        .y(_T_3190),
        .a(_T_3188),
        .b(32'h40)
    );
    wire [31:0] _T_3192;
    BITWISEAND #(.width(32)) bitwiseand_1699 (
        .y(_T_3192),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h70)
    );
    wire _T_3194;
    EQ_UNSIGNED #(.width(32)) u_eq_1700 (
        .y(_T_3194),
        .a(_T_3192),
        .b(32'h40)
    );
    wire _T_3196;
    BITWISEOR #(.width(1)) bitwiseor_1701 (
        .y(_T_3196),
        .a(1'h0),
        .b(_T_3186)
    );
    wire _T_3197;
    BITWISEOR #(.width(1)) bitwiseor_1702 (
        .y(_T_3197),
        .a(_T_3196),
        .b(_T_3190)
    );
    wire _T_3198;
    BITWISEOR #(.width(1)) bitwiseor_1703 (
        .y(_T_3198),
        .a(_T_3197),
        .b(_T_3194)
    );
    wire [31:0] _T_3200;
    BITWISEAND #(.width(32)) bitwiseand_1704 (
        .y(_T_3200),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h7C)
    );
    wire _T_3202;
    EQ_UNSIGNED #(.width(32)) u_eq_1705 (
        .y(_T_3202),
        .a(_T_3200),
        .b(32'h24)
    );
    wire [31:0] _T_3204;
    BITWISEAND #(.width(32)) bitwiseand_1706 (
        .y(_T_3204),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h40000060)
    );
    wire _T_3206;
    EQ_UNSIGNED #(.width(32)) u_eq_1707 (
        .y(_T_3206),
        .a(_T_3204),
        .b(32'h40)
    );
    wire [31:0] _T_3208;
    BITWISEAND #(.width(32)) bitwiseand_1708 (
        .y(_T_3208),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h90000060)
    );
    wire _T_3210;
    EQ_UNSIGNED #(.width(32)) u_eq_1709 (
        .y(_T_3210),
        .a(_T_3208),
        .b(32'h10000040)
    );
    wire _T_3212;
    BITWISEOR #(.width(1)) bitwiseor_1710 (
        .y(_T_3212),
        .a(1'h0),
        .b(_T_3202)
    );
    wire _T_3213;
    BITWISEOR #(.width(1)) bitwiseor_1711 (
        .y(_T_3213),
        .a(_T_3212),
        .b(_T_3206)
    );
    wire _T_3214;
    BITWISEOR #(.width(1)) bitwiseor_1712 (
        .y(_T_3214),
        .a(_T_3213),
        .b(_T_3194)
    );
    wire _T_3215;
    BITWISEOR #(.width(1)) bitwiseor_1713 (
        .y(_T_3215),
        .a(_T_3214),
        .b(_T_3210)
    );
    wire _T_3217;
    BITWISEOR #(.width(1)) bitwiseor_1714 (
        .y(_T_3217),
        .a(1'h0),
        .b(_T_3194)
    );
    wire [31:0] _T_3219;
    BITWISEAND #(.width(32)) bitwiseand_1715 (
        .y(_T_3219),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h3C)
    );
    wire _T_3221;
    EQ_UNSIGNED #(.width(32)) u_eq_1716 (
        .y(_T_3221),
        .a(_T_3219),
        .b(32'h4)
    );
    wire [31:0] _T_3223;
    BITWISEAND #(.width(32)) bitwiseand_1717 (
        .y(_T_3223),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h10000060)
    );
    wire _T_3225;
    EQ_UNSIGNED #(.width(32)) u_eq_1718 (
        .y(_T_3225),
        .a(_T_3223),
        .b(32'h10000040)
    );
    wire _T_3227;
    BITWISEOR #(.width(1)) bitwiseor_1719 (
        .y(_T_3227),
        .a(1'h0),
        .b(_T_3221)
    );
    wire _T_3228;
    BITWISEOR #(.width(1)) bitwiseor_1720 (
        .y(_T_3228),
        .a(_T_3227),
        .b(_T_3186)
    );
    wire _T_3229;
    BITWISEOR #(.width(1)) bitwiseor_1721 (
        .y(_T_3229),
        .a(_T_3228),
        .b(_T_3194)
    );
    wire _T_3230;
    BITWISEOR #(.width(1)) bitwiseor_1722 (
        .y(_T_3230),
        .a(_T_3229),
        .b(_T_3225)
    );
    wire [31:0] _T_3232;
    BITWISEAND #(.width(32)) bitwiseand_1723 (
        .y(_T_3232),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h2000074)
    );
    wire _T_3234;
    EQ_UNSIGNED #(.width(32)) u_eq_1724 (
        .y(_T_3234),
        .a(_T_3232),
        .b(32'h2000030)
    );
    wire _T_3236;
    BITWISEOR #(.width(1)) bitwiseor_1725 (
        .y(_T_3236),
        .a(1'h0),
        .b(_T_3234)
    );
    wire [31:0] _T_3238;
    BITWISEAND #(.width(32)) bitwiseand_1726 (
        .y(_T_3238),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h64)
    );
    wire _T_3240;
    EQ_UNSIGNED #(.width(32)) u_eq_1727 (
        .y(_T_3240),
        .a(_T_3238),
        .b(32'h0)
    );
    wire [31:0] _T_3242;
    BITWISEAND #(.width(32)) bitwiseand_1728 (
        .y(_T_3242),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h50)
    );
    wire _T_3244;
    EQ_UNSIGNED #(.width(32)) u_eq_1729 (
        .y(_T_3244),
        .a(_T_3242),
        .b(32'h10)
    );
    wire [31:0] _T_3246;
    BITWISEAND #(.width(32)) bitwiseand_1730 (
        .y(_T_3246),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h2024)
    );
    wire _T_3248;
    EQ_UNSIGNED #(.width(32)) u_eq_1731 (
        .y(_T_3248),
        .a(_T_3246),
        .b(32'h24)
    );
    wire [31:0] _T_3250;
    BITWISEAND #(.width(32)) bitwiseand_1732 (
        .y(_T_3250),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h28)
    );
    wire _T_3252;
    EQ_UNSIGNED #(.width(32)) u_eq_1733 (
        .y(_T_3252),
        .a(_T_3250),
        .b(32'h28)
    );
    wire [31:0] _T_3254;
    BITWISEAND #(.width(32)) bitwiseand_1734 (
        .y(_T_3254),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h1030)
    );
    wire _T_3256;
    EQ_UNSIGNED #(.width(32)) u_eq_1735 (
        .y(_T_3256),
        .a(_T_3254),
        .b(32'h1030)
    );
    wire [31:0] _T_3258;
    BITWISEAND #(.width(32)) bitwiseand_1736 (
        .y(_T_3258),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h2030)
    );
    wire _T_3260;
    EQ_UNSIGNED #(.width(32)) u_eq_1737 (
        .y(_T_3260),
        .a(_T_3258),
        .b(32'h2030)
    );
    wire [31:0] _T_3262;
    BITWISEAND #(.width(32)) bitwiseand_1738 (
        .y(_T_3262),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h90000010)
    );
    wire _T_3264;
    EQ_UNSIGNED #(.width(32)) u_eq_1739 (
        .y(_T_3264),
        .a(_T_3262),
        .b(32'h80000010)
    );
    wire _T_3266;
    BITWISEOR #(.width(1)) bitwiseor_1740 (
        .y(_T_3266),
        .a(1'h0),
        .b(_T_3240)
    );
    wire _T_3267;
    BITWISEOR #(.width(1)) bitwiseor_1741 (
        .y(_T_3267),
        .a(_T_3266),
        .b(_T_3244)
    );
    wire _T_3268;
    BITWISEOR #(.width(1)) bitwiseor_1742 (
        .y(_T_3268),
        .a(_T_3267),
        .b(_T_3248)
    );
    wire _T_3269;
    BITWISEOR #(.width(1)) bitwiseor_1743 (
        .y(_T_3269),
        .a(_T_3268),
        .b(_T_3252)
    );
    wire _T_3270;
    BITWISEOR #(.width(1)) bitwiseor_1744 (
        .y(_T_3270),
        .a(_T_3269),
        .b(_T_3256)
    );
    wire _T_3271;
    BITWISEOR #(.width(1)) bitwiseor_1745 (
        .y(_T_3271),
        .a(_T_3270),
        .b(_T_3260)
    );
    wire _T_3272;
    BITWISEOR #(.width(1)) bitwiseor_1746 (
        .y(_T_3272),
        .a(_T_3271),
        .b(_T_3264)
    );
    wire [31:0] _T_3274;
    BITWISEAND #(.width(32)) bitwiseand_1747 (
        .y(_T_3274),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h1070)
    );
    wire _T_3276;
    EQ_UNSIGNED #(.width(32)) u_eq_1748 (
        .y(_T_3276),
        .a(_T_3274),
        .b(32'h1070)
    );
    wire _T_3278;
    BITWISEOR #(.width(1)) bitwiseor_1749 (
        .y(_T_3278),
        .a(1'h0),
        .b(_T_3276)
    );
    wire [31:0] _T_3280;
    BITWISEAND #(.width(32)) bitwiseand_1750 (
        .y(_T_3280),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h2070)
    );
    wire _T_3282;
    EQ_UNSIGNED #(.width(32)) u_eq_1751 (
        .y(_T_3282),
        .a(_T_3280),
        .b(32'h2070)
    );
    wire _T_3284;
    BITWISEOR #(.width(1)) bitwiseor_1752 (
        .y(_T_3284),
        .a(1'h0),
        .b(_T_3282)
    );
    wire [31:0] _T_3286;
    BITWISEAND #(.width(32)) bitwiseand_1753 (
        .y(_T_3286),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h3070)
    );
    wire _T_3288;
    EQ_UNSIGNED #(.width(32)) u_eq_1754 (
        .y(_T_3288),
        .a(_T_3286),
        .b(32'h70)
    );
    wire _T_3290;
    BITWISEOR #(.width(1)) bitwiseor_1755 (
        .y(_T_3290),
        .a(1'h0),
        .b(_T_3288)
    );
    wire [1:0] _T_3291;
    CAT #(.width_a(1), .width_b(1)) cat_1756 (
        .y(_T_3291),
        .a(_T_3290),
        .b(_T_3284)
    );
    wire [2:0] _T_3292;
    CAT #(.width_a(2), .width_b(1)) cat_1757 (
        .y(_T_3292),
        .a(_T_3291),
        .b(_T_3278)
    );
    wire [31:0] _T_3294;
    BITWISEAND #(.width(32)) bitwiseand_1758 (
        .y(_T_3294),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h3058)
    );
    wire _T_3296;
    EQ_UNSIGNED #(.width(32)) u_eq_1759 (
        .y(_T_3296),
        .a(_T_3294),
        .b(32'h1008)
    );
    wire _T_3298;
    BITWISEOR #(.width(1)) bitwiseor_1760 (
        .y(_T_3298),
        .a(1'h0),
        .b(_T_3296)
    );
    wire [31:0] _T_3300;
    BITWISEAND #(.width(32)) bitwiseand_1761 (
        .y(_T_3300),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h3058)
    );
    wire _T_3302;
    EQ_UNSIGNED #(.width(32)) u_eq_1762 (
        .y(_T_3302),
        .a(_T_3300),
        .b(32'h8)
    );
    wire _T_3304;
    BITWISEOR #(.width(1)) bitwiseor_1763 (
        .y(_T_3304),
        .a(1'h0),
        .b(_T_3302)
    );
    wire [31:0] _T_3306;
    BITWISEAND #(.width(32)) bitwiseand_1764 (
        .y(_T_3306),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h6048)
    );
    wire _T_3308;
    EQ_UNSIGNED #(.width(32)) u_eq_1765 (
        .y(_T_3308),
        .a(_T_3306),
        .b(32'h2008)
    );
    wire _T_3310;
    BITWISEOR #(.width(1)) bitwiseor_1766 (
        .y(_T_3310),
        .a(1'h0),
        .b(_T_3308)
    );
    wire [31:0] _T_3312;
    BITWISEAND #(.width(32)) bitwiseand_1767 (
        .y(_T_3312),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h105C)
    );
    wire _T_3314;
    EQ_UNSIGNED #(.width(32)) u_eq_1768 (
        .y(_T_3314),
        .a(_T_3312),
        .b(32'h1004)
    );
    wire [31:0] _T_3316;
    BITWISEAND #(.width(32)) bitwiseand_1769 (
        .y(_T_3316),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'h2000060)
    );
    wire _T_3318;
    EQ_UNSIGNED #(.width(32)) u_eq_1770 (
        .y(_T_3318),
        .a(_T_3316),
        .b(32'h2000040)
    );
    wire [31:0] _T_3320;
    BITWISEAND #(.width(32)) bitwiseand_1771 (
        .y(_T_3320),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(32'hD0000070)
    );
    wire _T_3322;
    EQ_UNSIGNED #(.width(32)) u_eq_1772 (
        .y(_T_3322),
        .a(_T_3320),
        .b(32'h40000050)
    );
    wire _T_3324;
    BITWISEOR #(.width(1)) bitwiseor_1773 (
        .y(_T_3324),
        .a(1'h0),
        .b(_T_3314)
    );
    wire _T_3325;
    BITWISEOR #(.width(1)) bitwiseor_1774 (
        .y(_T_3325),
        .a(_T_3324),
        .b(_T_3318)
    );
    wire _T_3326;
    BITWISEOR #(.width(1)) bitwiseor_1775 (
        .y(_T_3326),
        .a(_T_3325),
        .b(_T_3322)
    );
    wire id_load_use;
    wire _id_reg_fence__q;
    wire _id_reg_fence__d;
    DFF_POSCLK #(.width(1)) id_reg_fence (
        .q(_id_reg_fence__q),
        .d(_id_reg_fence__d),
        .clk(clock)
    );
    wire _WTEMP_114;
    MUX_UNSIGNED #(.width(1)) u_mux_1776 (
        .y(_id_reg_fence__d),
        .sel(reset),
        .a(1'h0),
        .b(_WTEMP_114)
    );
    wire [63:0] _T_3331__T_3340_data;
    wire _T_3331__T_3340_clk;
    wire _T_3331__T_3340_en;
    wire [4:0] _T_3331__T_3340_addr;
    wire [63:0] _T_3331__T_3350_data;
    wire _T_3331__T_3350_clk;
    wire _T_3331__T_3350_en;
    wire [4:0] _T_3331__T_3350_addr;
    wire _T_3331__T_4200_clk;
    wire _T_3331__T_4200_en;
    wire _T_3331__T_4200_mask;
    wire [4:0] _T_3331__T_4200_addr;
    wire [63:0] _T_3331__T_4200_data;
    wire [127:0] _T_3331_read_datas;
    wire [1:0] _T_3331_read_clks;
    wire [1:0] _T_3331_read_ens;
    wire [9:0] _T_3331_read_addrs;
    wire _T_3331_write_clks;
    wire _T_3331_write_ens;
    wire _T_3331_write_masks;
    wire [4:0] _T_3331_write_addrs;
    wire [63:0] _T_3331_write_datas;
    BITS #(.width(128), .high(63), .low(0)) bits_1777 (
        .y(_T_3331__T_3340_data),
        .in(_T_3331_read_datas)
    );
    BITS #(.width(128), .high(127), .low(64)) bits_1778 (
        .y(_T_3331__T_3350_data),
        .in(_T_3331_read_datas)
    );
    CAT #(.width_a(1), .width_b(1)) cat_1779 (
        .y(_T_3331_read_clks),
        .a(_T_3331__T_3350_clk),
        .b(_T_3331__T_3340_clk)
    );
    CAT #(.width_a(1), .width_b(1)) cat_1780 (
        .y(_T_3331_read_ens),
        .a(_T_3331__T_3350_en),
        .b(_T_3331__T_3340_en)
    );
    CAT #(.width_a(5), .width_b(5)) cat_1781 (
        .y(_T_3331_read_addrs),
        .a(_T_3331__T_3350_addr),
        .b(_T_3331__T_3340_addr)
    );
    assign _T_3331_write_datas = _T_3331__T_4200_data;
    assign _T_3331_write_clks = _T_3331__T_4200_clk;
    assign _T_3331_write_ens = _T_3331__T_4200_en;
    assign _T_3331_write_addrs = _T_3331__T_4200_addr;
    assign _T_3331_write_masks = _T_3331__T_4200_mask;
    MRMWMEM #(.depth(31), .addrbits(5), .width(64), .readernum(2), .writernum(1), .isSyncRead(0)) _T_3331 (
        .read_datas(_T_3331_read_datas),
        .read_clks(_T_3331_read_clks),
        .read_ens(_T_3331_read_ens),
        .read_addrs(_T_3331_read_addrs),
        .write_clks(_T_3331_write_clks),
        .write_ens(_T_3331_write_ens),
        .write_masks(_T_3331_write_masks),
        .write_addrs(_T_3331_write_addrs),
        .write_datas(_T_3331_write_datas)
    );
    wire [63:0] id_rs_0;
    wire _T_3335;
    wire [4:0] _WTEMP_115;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_1782 (
        .y(_WTEMP_115),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(5)) u_eq_1783 (
        .y(_T_3335),
        .a(_ibuf__io_inst_0_bits_inst_rs1),
        .b(_WTEMP_115)
    );
    wire _T_3336;
    assign _T_3336 = 1'h0;
    wire [4:0] _T_3338;
    BITS #(.width(5), .high(4), .low(0)) bits_1784 (
        .y(_T_3338),
        .in(_ibuf__io_inst_0_bits_inst_rs1)
    );
    wire [4:0] _T_3339;
    BITWISENOT #(.width(5)) bitwisenot_1785 (
        .y(_T_3339),
        .in(_T_3338)
    );
    assign _T_3331__T_3340_addr = _T_3339;
    assign _T_3331__T_3340_en = 1'h1;
    assign _T_3331__T_3340_clk = clock;
    wire [63:0] _T_3341;
    assign _T_3341 = _T_3331__T_3340_data;
    wire [63:0] id_rs_1;
    wire _T_3345;
    wire [4:0] _WTEMP_116;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_1786 (
        .y(_WTEMP_116),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(5)) u_eq_1787 (
        .y(_T_3345),
        .a(_ibuf__io_inst_0_bits_inst_rs2),
        .b(_WTEMP_116)
    );
    wire _T_3346;
    assign _T_3346 = 1'h0;
    wire [4:0] _T_3348;
    BITS #(.width(5), .high(4), .low(0)) bits_1788 (
        .y(_T_3348),
        .in(_ibuf__io_inst_0_bits_inst_rs2)
    );
    wire [4:0] _T_3349;
    BITWISENOT #(.width(5)) bitwisenot_1789 (
        .y(_T_3349),
        .in(_T_3348)
    );
    assign _T_3331__T_3350_addr = _T_3349;
    assign _T_3331__T_3350_en = 1'h1;
    assign _T_3331__T_3350_clk = clock;
    wire [63:0] _T_3351;
    assign _T_3351 = _T_3331__T_3350_data;
    wire ctrl_killd;
    wire [39:0] _T_3353;
    ASSINT #(.width(40)) assint_1790 (
        .y(_T_3353),
        .in(_ibuf__io_pc)
    );
    wire _T_3356;
    assign _T_3356 = 1'h0;
    wire _T_3358;
    BITS #(.width(32), .high(31), .low(31)) bits_1791 (
        .y(_T_3358),
        .in(_ibuf__io_inst_0_bits_inst_bits)
    );
    wire _T_3359;
    ASSINT #(.width(1)) assint_1792 (
        .y(_T_3359),
        .in(_T_3358)
    );
    wire _T_3360;
    assign _T_3360 = _T_3359;
    wire _T_3362;
    assign _T_3362 = 1'h0;
    wire [10:0] _T_3363;
    BITS #(.width(32), .high(30), .low(20)) bits_1793 (
        .y(_T_3363),
        .in(_ibuf__io_inst_0_bits_inst_bits)
    );
    wire [10:0] _T_3364;
    ASSINT #(.width(11)) assint_1794 (
        .y(_T_3364),
        .in(_T_3363)
    );
    wire _T_3365;
    assign _T_3365 = _T_3360;
    wire _T_3367;
    assign _T_3367 = 1'h1;
    wire _T_3369;
    assign _T_3369 = 1'h0;
    wire _T_3370;
    assign _T_3370 = 1'h0;
    wire [7:0] _T_3371;
    BITS #(.width(32), .high(19), .low(12)) bits_1795 (
        .y(_T_3371),
        .in(_ibuf__io_inst_0_bits_inst_bits)
    );
    wire [7:0] _T_3372;
    ASSINT #(.width(8)) assint_1796 (
        .y(_T_3372),
        .in(_T_3371)
    );
    wire [7:0] _T_3373;
    assign _T_3373 = _T_3372;
    wire _T_3375;
    assign _T_3375 = 1'h0;
    wire _T_3377;
    assign _T_3377 = 1'h0;
    wire _T_3378;
    assign _T_3378 = 1'h0;
    wire _T_3381;
    assign _T_3381 = 1'h1;
    wire _T_3382;
    BITS #(.width(32), .high(20), .low(20)) bits_1797 (
        .y(_T_3382),
        .in(_ibuf__io_inst_0_bits_inst_bits)
    );
    wire _T_3383;
    ASSINT #(.width(1)) assint_1798 (
        .y(_T_3383),
        .in(_T_3382)
    );
    wire _T_3385;
    assign _T_3385 = 1'h0;
    wire _T_3386;
    BITS #(.width(32), .high(7), .low(7)) bits_1799 (
        .y(_T_3386),
        .in(_ibuf__io_inst_0_bits_inst_bits)
    );
    wire _T_3387;
    ASSINT #(.width(1)) assint_1800 (
        .y(_T_3387),
        .in(_T_3386)
    );
    wire _T_3388;
    assign _T_3388 = _T_3360;
    wire _T_3389;
    assign _T_3389 = _T_3383;
    wire _T_3390;
    assign _T_3390 = _T_3389;
    wire _T_3392;
    assign _T_3392 = 1'h0;
    wire _T_3394;
    assign _T_3394 = 1'h0;
    wire _T_3395;
    assign _T_3395 = 1'h0;
    wire [5:0] _T_3397;
    BITS #(.width(32), .high(30), .low(25)) bits_1801 (
        .y(_T_3397),
        .in(_ibuf__io_inst_0_bits_inst_bits)
    );
    wire [5:0] _T_3398;
    assign _T_3398 = _T_3397;
    wire _T_3400;
    assign _T_3400 = 1'h0;
    wire _T_3403;
    assign _T_3403 = 1'h0;
    wire _T_3405;
    assign _T_3405 = 1'h0;
    wire _T_3406;
    assign _T_3406 = 1'h0;
    wire [3:0] _T_3407;
    BITS #(.width(32), .high(11), .low(8)) bits_1802 (
        .y(_T_3407),
        .in(_ibuf__io_inst_0_bits_inst_bits)
    );
    wire _T_3409;
    assign _T_3409 = 1'h0;
    wire [3:0] _T_3410;
    BITS #(.width(32), .high(19), .low(16)) bits_1803 (
        .y(_T_3410),
        .in(_ibuf__io_inst_0_bits_inst_bits)
    );
    wire [3:0] _T_3411;
    BITS #(.width(32), .high(24), .low(21)) bits_1804 (
        .y(_T_3411),
        .in(_ibuf__io_inst_0_bits_inst_bits)
    );
    wire [3:0] _T_3412;
    assign _T_3412 = _T_3411;
    wire [3:0] _T_3413;
    assign _T_3413 = _T_3412;
    wire [3:0] _T_3414;
    assign _T_3414 = _T_3413;
    wire _T_3416;
    assign _T_3416 = 1'h0;
    wire _T_3417;
    BITS #(.width(32), .high(7), .low(7)) bits_1805 (
        .y(_T_3417),
        .in(_ibuf__io_inst_0_bits_inst_bits)
    );
    wire _T_3419;
    assign _T_3419 = 1'h0;
    wire _T_3420;
    BITS #(.width(32), .high(20), .low(20)) bits_1806 (
        .y(_T_3420),
        .in(_ibuf__io_inst_0_bits_inst_bits)
    );
    wire _T_3422;
    assign _T_3422 = 1'h0;
    wire _T_3423;
    BITS #(.width(32), .high(15), .low(15)) bits_1807 (
        .y(_T_3423),
        .in(_ibuf__io_inst_0_bits_inst_bits)
    );
    wire _T_3425;
    assign _T_3425 = 1'h0;
    wire _T_3426;
    assign _T_3426 = 1'h0;
    wire _T_3427;
    assign _T_3427 = 1'h0;
    wire [9:0] _T_3428;
    CAT #(.width_a(6), .width_b(4)) cat_1808 (
        .y(_T_3428),
        .a(_T_3398),
        .b(_T_3414)
    );
    wire [10:0] _T_3429;
    CAT #(.width_a(10), .width_b(1)) cat_1809 (
        .y(_T_3429),
        .a(_T_3428),
        .b(_T_3427)
    );
    wire _T_3430;
    ASUINT #(.width(1)) asuint_1810 (
        .y(_T_3430),
        .in(_T_3390)
    );
    wire [7:0] _T_3431;
    ASUINT #(.width(8)) asuint_1811 (
        .y(_T_3431),
        .in(_T_3373)
    );
    wire [8:0] _T_3432;
    CAT #(.width_a(8), .width_b(1)) cat_1812 (
        .y(_T_3432),
        .a(_T_3431),
        .b(_T_3430)
    );
    wire _T_3433;
    ASUINT #(.width(1)) asuint_1813 (
        .y(_T_3433),
        .in(_T_3365)
    );
    wire _T_3434;
    ASUINT #(.width(1)) asuint_1814 (
        .y(_T_3434),
        .in(_T_3360)
    );
    wire [1:0] _T_3435;
    CAT #(.width_a(1), .width_b(1)) cat_1815 (
        .y(_T_3435),
        .a(_T_3434),
        .b(_T_3433)
    );
    wire [10:0] _T_3436;
    CAT #(.width_a(2), .width_b(9)) cat_1816 (
        .y(_T_3436),
        .a(_T_3435),
        .b(_T_3432)
    );
    wire [21:0] _T_3437;
    CAT #(.width_a(11), .width_b(11)) cat_1817 (
        .y(_T_3437),
        .a(_T_3436),
        .b(_T_3429)
    );
    wire [21:0] _T_3438;
    ASSINT #(.width(22)) assint_1818 (
        .y(_T_3438),
        .in(_T_3437)
    );
    wire [40:0] _T_3439;
    wire [39:0] _WTEMP_117;
    PAD_SIGNED #(.width(22), .n(40)) s_pad_1819 (
        .y(_WTEMP_117),
        .in(_T_3438)
    );
    ADD_SIGNED #(.width(40)) s_add_1820 (
        .y(_T_3439),
        .a(_T_3353),
        .b(_WTEMP_117)
    );
    wire [39:0] _T_3440;
    TAIL #(.width(41), .n(1)) tail_1821 (
        .y(_T_3440),
        .in(_T_3439)
    );
    wire [39:0] _T_3441;
    ASSINT #(.width(40)) assint_1822 (
        .y(_T_3441),
        .in(_T_3440)
    );
    wire [39:0] id_npc;
    ASUINT #(.width(40)) asuint_1823 (
        .y(id_npc),
        .in(_T_3441)
    );
    wire _T_3444;
    EQ_UNSIGNED #(.width(1)) u_eq_1824 (
        .y(_T_3444),
        .a(ctrl_killd),
        .b(1'h0)
    );
    wire _T_3445;
    assign _T_3445 = 1'h0;
    wire _T_3446;
    assign _T_3446 = 1'h0;
    wire _csr__clock;
    wire _csr__reset;
    wire _csr__io_interrupts_debug;
    wire _csr__io_interrupts_mtip;
    wire _csr__io_interrupts_msip;
    wire _csr__io_interrupts_meip;
    wire _csr__io_interrupts_seip;
    wire [63:0] _csr__io_hartid;
    wire [11:0] _csr__io_rw_addr;
    wire [2:0] _csr__io_rw_cmd;
    wire [63:0] _csr__io_rw_rdata;
    wire [63:0] _csr__io_rw_wdata;
    wire [11:0] _csr__io_decode_csr;
    wire _csr__io_decode_fp_illegal;
    wire _csr__io_decode_rocc_illegal;
    wire _csr__io_decode_read_illegal;
    wire _csr__io_decode_write_illegal;
    wire _csr__io_decode_write_flush;
    wire _csr__io_decode_system_illegal;
    wire _csr__io_csr_stall;
    wire _csr__io_eret;
    wire _csr__io_singleStep;
    wire _csr__io_status_debug;
    wire [31:0] _csr__io_status_isa;
    wire [1:0] _csr__io_status_prv;
    wire _csr__io_status_sd;
    wire [26:0] _csr__io_status_zero2;
    wire [1:0] _csr__io_status_sxl;
    wire [1:0] _csr__io_status_uxl;
    wire _csr__io_status_sd_rv32;
    wire [7:0] _csr__io_status_zero1;
    wire _csr__io_status_tsr;
    wire _csr__io_status_tw;
    wire _csr__io_status_tvm;
    wire _csr__io_status_mxr;
    wire _csr__io_status_pum;
    wire _csr__io_status_mprv;
    wire [1:0] _csr__io_status_xs;
    wire [1:0] _csr__io_status_fs;
    wire [1:0] _csr__io_status_mpp;
    wire [1:0] _csr__io_status_hpp;
    wire _csr__io_status_spp;
    wire _csr__io_status_mpie;
    wire _csr__io_status_hpie;
    wire _csr__io_status_spie;
    wire _csr__io_status_upie;
    wire _csr__io_status_mie;
    wire _csr__io_status_hie;
    wire _csr__io_status_sie;
    wire _csr__io_status_uie;
    wire [3:0] _csr__io_ptbr_mode;
    wire [15:0] _csr__io_ptbr_asid;
    wire [43:0] _csr__io_ptbr_ppn;
    wire [39:0] _csr__io_evec;
    wire _csr__io_exception;
    wire _csr__io_retire;
    wire [63:0] _csr__io_cause;
    wire [39:0] _csr__io_pc;
    wire [39:0] _csr__io_badaddr;
    wire _csr__io_fatc;
    wire [63:0] _csr__io_time;
    wire [2:0] _csr__io_fcsr_rm;
    wire _csr__io_fcsr_flags_valid;
    wire [4:0] _csr__io_fcsr_flags_bits;
    wire _csr__io_rocc_interrupt;
    wire _csr__io_interrupt;
    wire [63:0] _csr__io_interrupt_cause;
    wire [3:0] _csr__io_bp_0_control_ttype;
    wire _csr__io_bp_0_control_dmode;
    wire [5:0] _csr__io_bp_0_control_maskmax;
    wire [39:0] _csr__io_bp_0_control_reserved;
    wire _csr__io_bp_0_control_action;
    wire _csr__io_bp_0_control_chain;
    wire [1:0] _csr__io_bp_0_control_zero;
    wire [1:0] _csr__io_bp_0_control_tmatch;
    wire _csr__io_bp_0_control_m;
    wire _csr__io_bp_0_control_h;
    wire _csr__io_bp_0_control_s;
    wire _csr__io_bp_0_control_u;
    wire _csr__io_bp_0_control_x;
    wire _csr__io_bp_0_control_w;
    wire _csr__io_bp_0_control_r;
    wire [38:0] _csr__io_bp_0_address;
    CSRFile csr (
        .clock(_csr__clock),
        .reset(_csr__reset),
        .io_interrupts_debug(_csr__io_interrupts_debug),
        .io_interrupts_mtip(_csr__io_interrupts_mtip),
        .io_interrupts_msip(_csr__io_interrupts_msip),
        .io_interrupts_meip(_csr__io_interrupts_meip),
        .io_interrupts_seip(_csr__io_interrupts_seip),
        .io_hartid(_csr__io_hartid),
        .io_rw_addr(_csr__io_rw_addr),
        .io_rw_cmd(_csr__io_rw_cmd),
        .io_rw_rdata(_csr__io_rw_rdata),
        .io_rw_wdata(_csr__io_rw_wdata),
        .io_decode_csr(_csr__io_decode_csr),
        .io_decode_fp_illegal(_csr__io_decode_fp_illegal),
        .io_decode_rocc_illegal(_csr__io_decode_rocc_illegal),
        .io_decode_read_illegal(_csr__io_decode_read_illegal),
        .io_decode_write_illegal(_csr__io_decode_write_illegal),
        .io_decode_write_flush(_csr__io_decode_write_flush),
        .io_decode_system_illegal(_csr__io_decode_system_illegal),
        .io_csr_stall(_csr__io_csr_stall),
        .io_eret(_csr__io_eret),
        .io_singleStep(_csr__io_singleStep),
        .io_status_debug(_csr__io_status_debug),
        .io_status_isa(_csr__io_status_isa),
        .io_status_prv(_csr__io_status_prv),
        .io_status_sd(_csr__io_status_sd),
        .io_status_zero2(_csr__io_status_zero2),
        .io_status_sxl(_csr__io_status_sxl),
        .io_status_uxl(_csr__io_status_uxl),
        .io_status_sd_rv32(_csr__io_status_sd_rv32),
        .io_status_zero1(_csr__io_status_zero1),
        .io_status_tsr(_csr__io_status_tsr),
        .io_status_tw(_csr__io_status_tw),
        .io_status_tvm(_csr__io_status_tvm),
        .io_status_mxr(_csr__io_status_mxr),
        .io_status_pum(_csr__io_status_pum),
        .io_status_mprv(_csr__io_status_mprv),
        .io_status_xs(_csr__io_status_xs),
        .io_status_fs(_csr__io_status_fs),
        .io_status_mpp(_csr__io_status_mpp),
        .io_status_hpp(_csr__io_status_hpp),
        .io_status_spp(_csr__io_status_spp),
        .io_status_mpie(_csr__io_status_mpie),
        .io_status_hpie(_csr__io_status_hpie),
        .io_status_spie(_csr__io_status_spie),
        .io_status_upie(_csr__io_status_upie),
        .io_status_mie(_csr__io_status_mie),
        .io_status_hie(_csr__io_status_hie),
        .io_status_sie(_csr__io_status_sie),
        .io_status_uie(_csr__io_status_uie),
        .io_ptbr_mode(_csr__io_ptbr_mode),
        .io_ptbr_asid(_csr__io_ptbr_asid),
        .io_ptbr_ppn(_csr__io_ptbr_ppn),
        .io_evec(_csr__io_evec),
        .io_exception(_csr__io_exception),
        .io_retire(_csr__io_retire),
        .io_cause(_csr__io_cause),
        .io_pc(_csr__io_pc),
        .io_badaddr(_csr__io_badaddr),
        .io_fatc(_csr__io_fatc),
        .io_time(_csr__io_time),
        .io_fcsr_rm(_csr__io_fcsr_rm),
        .io_fcsr_flags_valid(_csr__io_fcsr_flags_valid),
        .io_fcsr_flags_bits(_csr__io_fcsr_flags_bits),
        .io_rocc_interrupt(_csr__io_rocc_interrupt),
        .io_interrupt(_csr__io_interrupt),
        .io_interrupt_cause(_csr__io_interrupt_cause),
        .io_bp_0_control_ttype(_csr__io_bp_0_control_ttype),
        .io_bp_0_control_dmode(_csr__io_bp_0_control_dmode),
        .io_bp_0_control_maskmax(_csr__io_bp_0_control_maskmax),
        .io_bp_0_control_reserved(_csr__io_bp_0_control_reserved),
        .io_bp_0_control_action(_csr__io_bp_0_control_action),
        .io_bp_0_control_chain(_csr__io_bp_0_control_chain),
        .io_bp_0_control_zero(_csr__io_bp_0_control_zero),
        .io_bp_0_control_tmatch(_csr__io_bp_0_control_tmatch),
        .io_bp_0_control_m(_csr__io_bp_0_control_m),
        .io_bp_0_control_h(_csr__io_bp_0_control_h),
        .io_bp_0_control_s(_csr__io_bp_0_control_s),
        .io_bp_0_control_u(_csr__io_bp_0_control_u),
        .io_bp_0_control_x(_csr__io_bp_0_control_x),
        .io_bp_0_control_w(_csr__io_bp_0_control_w),
        .io_bp_0_control_r(_csr__io_bp_0_control_r),
        .io_bp_0_address(_csr__io_bp_0_address)
    );
    wire _T_3450;
    EQ_UNSIGNED #(.width(3)) u_eq_3884 (
        .y(_T_3450),
        .a(id_ctrl_csr),
        .b(3'h2)
    );
    wire _T_3451;
    EQ_UNSIGNED #(.width(3)) u_eq_3885 (
        .y(_T_3451),
        .a(id_ctrl_csr),
        .b(3'h3)
    );
    wire _T_3452;
    EQ_UNSIGNED #(.width(3)) u_eq_3886 (
        .y(_T_3452),
        .a(id_ctrl_csr),
        .b(3'h1)
    );
    wire _T_3453;
    BITWISEOR #(.width(1)) bitwiseor_3887 (
        .y(_T_3453),
        .a(_T_3450),
        .b(_T_3451)
    );
    wire id_csr_en;
    BITWISEOR #(.width(1)) bitwiseor_3888 (
        .y(id_csr_en),
        .a(_T_3453),
        .b(_T_3452)
    );
    wire id_system_insn;
    GEQ_UNSIGNED #(.width(3)) u_geq_3889 (
        .y(id_system_insn),
        .a(id_ctrl_csr),
        .b(3'h4)
    );
    wire _T_3457;
    EQ_UNSIGNED #(.width(3)) u_eq_3890 (
        .y(_T_3457),
        .a(id_ctrl_csr),
        .b(3'h2)
    );
    wire _T_3458;
    EQ_UNSIGNED #(.width(3)) u_eq_3891 (
        .y(_T_3458),
        .a(id_ctrl_csr),
        .b(3'h3)
    );
    wire _T_3459;
    BITWISEOR #(.width(1)) bitwiseor_3892 (
        .y(_T_3459),
        .a(_T_3457),
        .b(_T_3458)
    );
    wire _T_3461;
    wire [4:0] _WTEMP_563;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_3893 (
        .y(_WTEMP_563),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(5)) u_eq_3894 (
        .y(_T_3461),
        .a(_ibuf__io_inst_0_bits_inst_rs1),
        .b(_WTEMP_563)
    );
    wire id_csr_ren;
    BITWISEAND #(.width(1)) bitwiseand_3895 (
        .y(id_csr_ren),
        .a(_T_3459),
        .b(_T_3461)
    );
    wire [2:0] id_csr;
    MUX_UNSIGNED #(.width(3)) u_mux_3896 (
        .y(id_csr),
        .sel(id_csr_ren),
        .a(3'h5),
        .b(id_ctrl_csr)
    );
    wire _T_3464;
    EQ_UNSIGNED #(.width(1)) u_eq_3897 (
        .y(_T_3464),
        .a(id_csr_ren),
        .b(1'h0)
    );
    wire _T_3465;
    BITWISEAND #(.width(1)) bitwiseand_3898 (
        .y(_T_3465),
        .a(id_csr_en),
        .b(_T_3464)
    );
    wire _T_3466;
    BITWISEAND #(.width(1)) bitwiseand_3899 (
        .y(_T_3466),
        .a(_T_3465),
        .b(_csr__io_decode_write_flush)
    );
    wire id_csr_flush;
    BITWISEOR #(.width(1)) bitwiseor_3900 (
        .y(id_csr_flush),
        .a(id_system_insn),
        .b(_T_3466)
    );
    wire _T_3468;
    EQ_UNSIGNED #(.width(1)) u_eq_3901 (
        .y(_T_3468),
        .a(id_ctrl_legal),
        .b(1'h0)
    );
    wire _T_3469;
    BITS #(.width(32), .high(12), .low(12)) bits_3902 (
        .y(_T_3469),
        .in(_csr__io_status_isa)
    );
    wire _T_3471;
    EQ_UNSIGNED #(.width(1)) u_eq_3903 (
        .y(_T_3471),
        .a(_T_3469),
        .b(1'h0)
    );
    wire _T_3472;
    BITWISEAND #(.width(1)) bitwiseand_3904 (
        .y(_T_3472),
        .a(id_ctrl_div),
        .b(_T_3471)
    );
    wire _T_3473;
    BITWISEOR #(.width(1)) bitwiseor_3905 (
        .y(_T_3473),
        .a(_T_3468),
        .b(_T_3472)
    );
    wire _T_3474;
    BITS #(.width(32), .high(0), .low(0)) bits_3906 (
        .y(_T_3474),
        .in(_csr__io_status_isa)
    );
    wire _T_3476;
    EQ_UNSIGNED #(.width(1)) u_eq_3907 (
        .y(_T_3476),
        .a(_T_3474),
        .b(1'h0)
    );
    wire _T_3477;
    BITWISEAND #(.width(1)) bitwiseand_3908 (
        .y(_T_3477),
        .a(id_ctrl_amo),
        .b(_T_3476)
    );
    wire _T_3478;
    BITWISEOR #(.width(1)) bitwiseor_3909 (
        .y(_T_3478),
        .a(_T_3473),
        .b(_T_3477)
    );
    wire _T_3479;
    BITWISEOR #(.width(1)) bitwiseor_3910 (
        .y(_T_3479),
        .a(_csr__io_decode_fp_illegal),
        .b(io_fpu_illegal_rm)
    );
    wire _T_3480;
    BITWISEAND #(.width(1)) bitwiseand_3911 (
        .y(_T_3480),
        .a(id_ctrl_fp),
        .b(_T_3479)
    );
    wire _T_3481;
    BITWISEOR #(.width(1)) bitwiseor_3912 (
        .y(_T_3481),
        .a(_T_3478),
        .b(_T_3480)
    );
    wire _T_3482;
    BITS #(.width(32), .high(3), .low(3)) bits_3913 (
        .y(_T_3482),
        .in(_csr__io_status_isa)
    );
    wire _T_3484;
    EQ_UNSIGNED #(.width(1)) u_eq_3914 (
        .y(_T_3484),
        .a(_T_3482),
        .b(1'h0)
    );
    wire _T_3485;
    BITWISEAND #(.width(1)) bitwiseand_3915 (
        .y(_T_3485),
        .a(id_ctrl_dp),
        .b(_T_3484)
    );
    wire _T_3486;
    BITWISEOR #(.width(1)) bitwiseor_3916 (
        .y(_T_3486),
        .a(_T_3481),
        .b(_T_3485)
    );
    wire _T_3487;
    BITS #(.width(32), .high(2), .low(2)) bits_3917 (
        .y(_T_3487),
        .in(_csr__io_status_isa)
    );
    wire _T_3489;
    EQ_UNSIGNED #(.width(1)) u_eq_3918 (
        .y(_T_3489),
        .a(_T_3487),
        .b(1'h0)
    );
    wire _T_3490;
    BITWISEAND #(.width(1)) bitwiseand_3919 (
        .y(_T_3490),
        .a(_ibuf__io_inst_0_bits_rvc),
        .b(_T_3489)
    );
    wire _T_3491;
    BITWISEOR #(.width(1)) bitwiseor_3920 (
        .y(_T_3491),
        .a(_T_3486),
        .b(_T_3490)
    );
    wire _T_3492;
    BITWISEAND #(.width(1)) bitwiseand_3921 (
        .y(_T_3492),
        .a(id_ctrl_rocc),
        .b(_csr__io_decode_rocc_illegal)
    );
    wire _T_3493;
    BITWISEOR #(.width(1)) bitwiseor_3922 (
        .y(_T_3493),
        .a(_T_3491),
        .b(_T_3492)
    );
    wire _T_3495;
    EQ_UNSIGNED #(.width(1)) u_eq_3923 (
        .y(_T_3495),
        .a(id_csr_ren),
        .b(1'h0)
    );
    wire _T_3496;
    BITWISEAND #(.width(1)) bitwiseand_3924 (
        .y(_T_3496),
        .a(_T_3495),
        .b(_csr__io_decode_write_illegal)
    );
    wire _T_3497;
    BITWISEOR #(.width(1)) bitwiseor_3925 (
        .y(_T_3497),
        .a(_csr__io_decode_read_illegal),
        .b(_T_3496)
    );
    wire _T_3498;
    BITWISEAND #(.width(1)) bitwiseand_3926 (
        .y(_T_3498),
        .a(id_csr_en),
        .b(_T_3497)
    );
    wire _T_3499;
    BITWISEOR #(.width(1)) bitwiseor_3927 (
        .y(_T_3499),
        .a(_T_3493),
        .b(_T_3498)
    );
    wire _T_3500;
    BITWISEAND #(.width(1)) bitwiseand_3928 (
        .y(_T_3500),
        .a(id_system_insn),
        .b(_csr__io_decode_system_illegal)
    );
    wire id_illegal_insn;
    BITWISEOR #(.width(1)) bitwiseor_3929 (
        .y(id_illegal_insn),
        .a(_T_3499),
        .b(_T_3500)
    );
    wire id_amo_aq;
    BITS #(.width(32), .high(26), .low(26)) bits_3930 (
        .y(id_amo_aq),
        .in(_ibuf__io_inst_0_bits_inst_bits)
    );
    wire id_amo_rl;
    BITS #(.width(32), .high(25), .low(25)) bits_3931 (
        .y(id_amo_rl),
        .in(_ibuf__io_inst_0_bits_inst_bits)
    );
    wire _T_3501;
    BITWISEAND #(.width(1)) bitwiseand_3932 (
        .y(_T_3501),
        .a(id_ctrl_amo),
        .b(id_amo_rl)
    );
    wire id_fence_next;
    BITWISEOR #(.width(1)) bitwiseor_3933 (
        .y(id_fence_next),
        .a(id_ctrl_fence),
        .b(_T_3501)
    );
    wire _T_3503;
    EQ_UNSIGNED #(.width(1)) u_eq_3934 (
        .y(_T_3503),
        .a(io_dmem_ordered),
        .b(1'h0)
    );
    wire id_mem_busy;
    BITWISEOR #(.width(1)) bitwiseor_3935 (
        .y(id_mem_busy),
        .a(_T_3503),
        .b(io_dmem_req_valid)
    );
    wire _T_3505;
    assign _T_3505 = 1'h0;
    wire _T_3506;
    BITWISEOR #(.width(1)) bitwiseor_3936 (
        .y(_T_3506),
        .a(io_rocc_busy),
        .b(_T_3505)
    );
    wire _T_3507;
    assign _T_3507 = 1'h0;
    wire _T_3508;
    BITWISEOR #(.width(1)) bitwiseor_3937 (
        .y(_T_3508),
        .a(_T_3506),
        .b(_T_3507)
    );
    wire _T_3509;
    assign _T_3509 = 1'h0;
    wire _T_3510;
    BITWISEOR #(.width(1)) bitwiseor_3938 (
        .y(_T_3510),
        .a(_T_3508),
        .b(_T_3509)
    );
    wire id_rocc_busy;
    assign id_rocc_busy = 1'h0;
    wire _T_3511;
    BITWISEAND #(.width(1)) bitwiseand_3939 (
        .y(_T_3511),
        .a(_id_reg_fence__q),
        .b(id_mem_busy)
    );
    wire _T_3512;
    BITWISEOR #(.width(1)) bitwiseor_3940 (
        .y(_T_3512),
        .a(id_fence_next),
        .b(_T_3511)
    );
    wire _T_3513;
    assign _T_3513 = 1'h0;
    wire _T_3514;
    BITWISEAND #(.width(1)) bitwiseand_3941 (
        .y(_T_3514),
        .a(id_ctrl_amo),
        .b(id_amo_aq)
    );
    wire _T_3515;
    BITWISEOR #(.width(1)) bitwiseor_3942 (
        .y(_T_3515),
        .a(_T_3514),
        .b(id_ctrl_fence_i)
    );
    wire _T_3516;
    BITWISEOR #(.width(1)) bitwiseor_3943 (
        .y(_T_3516),
        .a(id_ctrl_mem),
        .b(id_ctrl_rocc)
    );
    wire _T_3517;
    BITWISEAND #(.width(1)) bitwiseand_3944 (
        .y(_T_3517),
        .a(_id_reg_fence__q),
        .b(_T_3516)
    );
    wire _T_3518;
    BITWISEOR #(.width(1)) bitwiseor_3945 (
        .y(_T_3518),
        .a(_T_3515),
        .b(_T_3517)
    );
    wire _T_3519;
    BITWISEAND #(.width(1)) bitwiseand_3946 (
        .y(_T_3519),
        .a(id_mem_busy),
        .b(_T_3518)
    );
    wire id_do_fence;
    BITWISEOR #(.width(1)) bitwiseor_3947 (
        .y(id_do_fence),
        .a(_T_3513),
        .b(_T_3519)
    );
    wire _bpu__clock;
    wire _bpu__reset;
    wire _bpu__io_status_debug;
    wire [31:0] _bpu__io_status_isa;
    wire [1:0] _bpu__io_status_prv;
    wire _bpu__io_status_sd;
    wire [26:0] _bpu__io_status_zero2;
    wire [1:0] _bpu__io_status_sxl;
    wire [1:0] _bpu__io_status_uxl;
    wire _bpu__io_status_sd_rv32;
    wire [7:0] _bpu__io_status_zero1;
    wire _bpu__io_status_tsr;
    wire _bpu__io_status_tw;
    wire _bpu__io_status_tvm;
    wire _bpu__io_status_mxr;
    wire _bpu__io_status_pum;
    wire _bpu__io_status_mprv;
    wire [1:0] _bpu__io_status_xs;
    wire [1:0] _bpu__io_status_fs;
    wire [1:0] _bpu__io_status_mpp;
    wire [1:0] _bpu__io_status_hpp;
    wire _bpu__io_status_spp;
    wire _bpu__io_status_mpie;
    wire _bpu__io_status_hpie;
    wire _bpu__io_status_spie;
    wire _bpu__io_status_upie;
    wire _bpu__io_status_mie;
    wire _bpu__io_status_hie;
    wire _bpu__io_status_sie;
    wire _bpu__io_status_uie;
    wire [3:0] _bpu__io_bp_0_control_ttype;
    wire _bpu__io_bp_0_control_dmode;
    wire [5:0] _bpu__io_bp_0_control_maskmax;
    wire [39:0] _bpu__io_bp_0_control_reserved;
    wire _bpu__io_bp_0_control_action;
    wire _bpu__io_bp_0_control_chain;
    wire [1:0] _bpu__io_bp_0_control_zero;
    wire [1:0] _bpu__io_bp_0_control_tmatch;
    wire _bpu__io_bp_0_control_m;
    wire _bpu__io_bp_0_control_h;
    wire _bpu__io_bp_0_control_s;
    wire _bpu__io_bp_0_control_u;
    wire _bpu__io_bp_0_control_x;
    wire _bpu__io_bp_0_control_w;
    wire _bpu__io_bp_0_control_r;
    wire [38:0] _bpu__io_bp_0_address;
    wire [38:0] _bpu__io_pc;
    wire [38:0] _bpu__io_ea;
    wire _bpu__io_xcpt_if;
    wire _bpu__io_xcpt_ld;
    wire _bpu__io_xcpt_st;
    wire _bpu__io_debug_if;
    wire _bpu__io_debug_ld;
    wire _bpu__io_debug_st;
    BreakpointUnit bpu (
        .clock(_bpu__clock),
        .reset(_bpu__reset),
        .io_status_debug(_bpu__io_status_debug),
        .io_status_isa(_bpu__io_status_isa),
        .io_status_prv(_bpu__io_status_prv),
        .io_status_sd(_bpu__io_status_sd),
        .io_status_zero2(_bpu__io_status_zero2),
        .io_status_sxl(_bpu__io_status_sxl),
        .io_status_uxl(_bpu__io_status_uxl),
        .io_status_sd_rv32(_bpu__io_status_sd_rv32),
        .io_status_zero1(_bpu__io_status_zero1),
        .io_status_tsr(_bpu__io_status_tsr),
        .io_status_tw(_bpu__io_status_tw),
        .io_status_tvm(_bpu__io_status_tvm),
        .io_status_mxr(_bpu__io_status_mxr),
        .io_status_pum(_bpu__io_status_pum),
        .io_status_mprv(_bpu__io_status_mprv),
        .io_status_xs(_bpu__io_status_xs),
        .io_status_fs(_bpu__io_status_fs),
        .io_status_mpp(_bpu__io_status_mpp),
        .io_status_hpp(_bpu__io_status_hpp),
        .io_status_spp(_bpu__io_status_spp),
        .io_status_mpie(_bpu__io_status_mpie),
        .io_status_hpie(_bpu__io_status_hpie),
        .io_status_spie(_bpu__io_status_spie),
        .io_status_upie(_bpu__io_status_upie),
        .io_status_mie(_bpu__io_status_mie),
        .io_status_hie(_bpu__io_status_hie),
        .io_status_sie(_bpu__io_status_sie),
        .io_status_uie(_bpu__io_status_uie),
        .io_bp_0_control_ttype(_bpu__io_bp_0_control_ttype),
        .io_bp_0_control_dmode(_bpu__io_bp_0_control_dmode),
        .io_bp_0_control_maskmax(_bpu__io_bp_0_control_maskmax),
        .io_bp_0_control_reserved(_bpu__io_bp_0_control_reserved),
        .io_bp_0_control_action(_bpu__io_bp_0_control_action),
        .io_bp_0_control_chain(_bpu__io_bp_0_control_chain),
        .io_bp_0_control_zero(_bpu__io_bp_0_control_zero),
        .io_bp_0_control_tmatch(_bpu__io_bp_0_control_tmatch),
        .io_bp_0_control_m(_bpu__io_bp_0_control_m),
        .io_bp_0_control_h(_bpu__io_bp_0_control_h),
        .io_bp_0_control_s(_bpu__io_bp_0_control_s),
        .io_bp_0_control_u(_bpu__io_bp_0_control_u),
        .io_bp_0_control_x(_bpu__io_bp_0_control_x),
        .io_bp_0_control_w(_bpu__io_bp_0_control_w),
        .io_bp_0_control_r(_bpu__io_bp_0_control_r),
        .io_bp_0_address(_bpu__io_bp_0_address),
        .io_pc(_bpu__io_pc),
        .io_ea(_bpu__io_ea),
        .io_xcpt_if(_bpu__io_xcpt_if),
        .io_xcpt_ld(_bpu__io_xcpt_ld),
        .io_xcpt_st(_bpu__io_xcpt_st),
        .io_debug_if(_bpu__io_debug_if),
        .io_debug_ld(_bpu__io_debug_ld),
        .io_debug_st(_bpu__io_debug_st)
    );
    wire id_xcpt_if;
    BITWISEOR #(.width(1)) bitwiseor_4076 (
        .y(id_xcpt_if),
        .a(_ibuf__io_inst_0_bits_pf0),
        .b(_ibuf__io_inst_0_bits_pf1)
    );
    wire _T_3552;
    BITWISEOR #(.width(1)) bitwiseor_4077 (
        .y(_T_3552),
        .a(_csr__io_interrupt),
        .b(_bpu__io_debug_if)
    );
    wire _T_3553;
    BITWISEOR #(.width(1)) bitwiseor_4078 (
        .y(_T_3553),
        .a(_T_3552),
        .b(_bpu__io_xcpt_if)
    );
    wire _T_3554;
    BITWISEOR #(.width(1)) bitwiseor_4079 (
        .y(_T_3554),
        .a(_T_3553),
        .b(id_xcpt_if)
    );
    wire id_xcpt;
    BITWISEOR #(.width(1)) bitwiseor_4080 (
        .y(id_xcpt),
        .a(_T_3554),
        .b(id_illegal_insn)
    );
    wire [1:0] _T_3555;
    wire [1:0] _WTEMP_570;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_4081 (
        .y(_WTEMP_570),
        .in(1'h1)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_4082 (
        .y(_T_3555),
        .sel(id_xcpt_if),
        .a(_WTEMP_570),
        .b(2'h2)
    );
    wire [1:0] _T_3556;
    MUX_UNSIGNED #(.width(2)) u_mux_4083 (
        .y(_T_3556),
        .sel(_bpu__io_xcpt_if),
        .a(2'h3),
        .b(_T_3555)
    );
    wire [3:0] _T_3557;
    wire [3:0] _WTEMP_571;
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_4084 (
        .y(_WTEMP_571),
        .in(_T_3556)
    );
    MUX_UNSIGNED #(.width(4)) u_mux_4085 (
        .y(_T_3557),
        .sel(_bpu__io_debug_if),
        .a(4'hD),
        .b(_WTEMP_571)
    );
    wire [63:0] id_cause;
    wire [63:0] _WTEMP_572;
    PAD_UNSIGNED #(.width(4), .n(64)) u_pad_4086 (
        .y(_WTEMP_572),
        .in(_T_3557)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_4087 (
        .y(id_cause),
        .sel(_csr__io_interrupt),
        .a(_csr__io_interrupt_cause),
        .b(_WTEMP_572)
    );
    wire [4:0] ex_waddr;
    BITS #(.width(32), .high(11), .low(7)) bits_4088 (
        .y(ex_waddr),
        .in(_ex_reg_inst__q)
    );
    wire [4:0] mem_waddr;
    BITS #(.width(32), .high(11), .low(7)) bits_4089 (
        .y(mem_waddr),
        .in(_mem_reg_inst__q)
    );
    wire [4:0] wb_waddr;
    BITS #(.width(32), .high(11), .low(7)) bits_4090 (
        .y(wb_waddr),
        .in(_wb_reg_inst__q)
    );
    wire _T_3561;
    BITWISEAND #(.width(1)) bitwiseand_4091 (
        .y(_T_3561),
        .a(_ex_reg_valid__q),
        .b(_ex_ctrl_wxd__q)
    );
    wire _T_3562;
    BITWISEAND #(.width(1)) bitwiseand_4092 (
        .y(_T_3562),
        .a(_mem_reg_valid__q),
        .b(_mem_ctrl_wxd__q)
    );
    wire _T_3564;
    EQ_UNSIGNED #(.width(1)) u_eq_4093 (
        .y(_T_3564),
        .a(_mem_ctrl_mem__q),
        .b(1'h0)
    );
    wire _T_3565;
    BITWISEAND #(.width(1)) bitwiseand_4094 (
        .y(_T_3565),
        .a(_T_3562),
        .b(_T_3564)
    );
    wire _T_3566;
    BITWISEAND #(.width(1)) bitwiseand_4095 (
        .y(_T_3566),
        .a(_mem_reg_valid__q),
        .b(_mem_ctrl_wxd__q)
    );
    wire _T_3567;
    wire [4:0] _WTEMP_573;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_4096 (
        .y(_WTEMP_573),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(5)) u_eq_4097 (
        .y(_T_3567),
        .a(_WTEMP_573),
        .b(_ibuf__io_inst_0_bits_inst_rs1)
    );
    wire id_bypass_src_0_0;
    BITWISEAND #(.width(1)) bitwiseand_4098 (
        .y(id_bypass_src_0_0),
        .a(1'h1),
        .b(_T_3567)
    );
    wire _T_3568;
    EQ_UNSIGNED #(.width(5)) u_eq_4099 (
        .y(_T_3568),
        .a(ex_waddr),
        .b(_ibuf__io_inst_0_bits_inst_rs1)
    );
    wire id_bypass_src_0_1;
    BITWISEAND #(.width(1)) bitwiseand_4100 (
        .y(id_bypass_src_0_1),
        .a(_T_3561),
        .b(_T_3568)
    );
    wire _T_3569;
    EQ_UNSIGNED #(.width(5)) u_eq_4101 (
        .y(_T_3569),
        .a(mem_waddr),
        .b(_ibuf__io_inst_0_bits_inst_rs1)
    );
    wire id_bypass_src_0_2;
    BITWISEAND #(.width(1)) bitwiseand_4102 (
        .y(id_bypass_src_0_2),
        .a(_T_3565),
        .b(_T_3569)
    );
    wire _T_3570;
    EQ_UNSIGNED #(.width(5)) u_eq_4103 (
        .y(_T_3570),
        .a(mem_waddr),
        .b(_ibuf__io_inst_0_bits_inst_rs1)
    );
    wire id_bypass_src_0_3;
    BITWISEAND #(.width(1)) bitwiseand_4104 (
        .y(id_bypass_src_0_3),
        .a(_T_3566),
        .b(_T_3570)
    );
    wire _T_3571;
    wire [4:0] _WTEMP_574;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_4105 (
        .y(_WTEMP_574),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(5)) u_eq_4106 (
        .y(_T_3571),
        .a(_WTEMP_574),
        .b(_ibuf__io_inst_0_bits_inst_rs2)
    );
    wire id_bypass_src_1_0;
    BITWISEAND #(.width(1)) bitwiseand_4107 (
        .y(id_bypass_src_1_0),
        .a(1'h1),
        .b(_T_3571)
    );
    wire _T_3572;
    EQ_UNSIGNED #(.width(5)) u_eq_4108 (
        .y(_T_3572),
        .a(ex_waddr),
        .b(_ibuf__io_inst_0_bits_inst_rs2)
    );
    wire id_bypass_src_1_1;
    BITWISEAND #(.width(1)) bitwiseand_4109 (
        .y(id_bypass_src_1_1),
        .a(_T_3561),
        .b(_T_3572)
    );
    wire _T_3573;
    EQ_UNSIGNED #(.width(5)) u_eq_4110 (
        .y(_T_3573),
        .a(mem_waddr),
        .b(_ibuf__io_inst_0_bits_inst_rs2)
    );
    wire id_bypass_src_1_2;
    BITWISEAND #(.width(1)) bitwiseand_4111 (
        .y(id_bypass_src_1_2),
        .a(_T_3565),
        .b(_T_3573)
    );
    wire _T_3574;
    EQ_UNSIGNED #(.width(5)) u_eq_4112 (
        .y(_T_3574),
        .a(mem_waddr),
        .b(_ibuf__io_inst_0_bits_inst_rs2)
    );
    wire id_bypass_src_1_3;
    BITWISEAND #(.width(1)) bitwiseand_4113 (
        .y(id_bypass_src_1_3),
        .a(_T_3566),
        .b(_T_3574)
    );
    wire [63:0] bypass_mux_0;
    wire [63:0] bypass_mux_1;
    wire [63:0] bypass_mux_2;
    wire [63:0] bypass_mux_3;
    wire _ex_reg_rs_bypass_0__q;
    wire _ex_reg_rs_bypass_0__d;
    DFF_POSCLK #(.width(1)) ex_reg_rs_bypass_0 (
        .q(_ex_reg_rs_bypass_0__q),
        .d(_ex_reg_rs_bypass_0__d),
        .clk(clock)
    );
    wire _ex_reg_rs_bypass_1__q;
    wire _ex_reg_rs_bypass_1__d;
    DFF_POSCLK #(.width(1)) ex_reg_rs_bypass_1 (
        .q(_ex_reg_rs_bypass_1__q),
        .d(_ex_reg_rs_bypass_1__d),
        .clk(clock)
    );
    wire [1:0] _ex_reg_rs_lsb_0__q;
    wire [1:0] _ex_reg_rs_lsb_0__d;
    DFF_POSCLK #(.width(2)) ex_reg_rs_lsb_0 (
        .q(_ex_reg_rs_lsb_0__q),
        .d(_ex_reg_rs_lsb_0__d),
        .clk(clock)
    );
    wire [1:0] _ex_reg_rs_lsb_1__q;
    wire [1:0] _ex_reg_rs_lsb_1__d;
    DFF_POSCLK #(.width(2)) ex_reg_rs_lsb_1 (
        .q(_ex_reg_rs_lsb_1__q),
        .d(_ex_reg_rs_lsb_1__d),
        .clk(clock)
    );
    wire [61:0] _ex_reg_rs_msb_0__q;
    wire [61:0] _ex_reg_rs_msb_0__d;
    DFF_POSCLK #(.width(62)) ex_reg_rs_msb_0 (
        .q(_ex_reg_rs_msb_0__q),
        .d(_ex_reg_rs_msb_0__d),
        .clk(clock)
    );
    wire [61:0] _ex_reg_rs_msb_1__q;
    wire [61:0] _ex_reg_rs_msb_1__d;
    DFF_POSCLK #(.width(62)) ex_reg_rs_msb_1 (
        .q(_ex_reg_rs_msb_1__q),
        .d(_ex_reg_rs_msb_1__d),
        .clk(clock)
    );
    wire [63:0] _T_3605;
    CAT #(.width_a(62), .width_b(2)) cat_4114 (
        .y(_T_3605),
        .a(_ex_reg_rs_msb_0__q),
        .b(_ex_reg_rs_lsb_0__q)
    );
    wire _node_324;
    EQ_UNSIGNED #(.width(2)) u_eq_4115 (
        .y(_node_324),
        .a(2'd0),
        .b(_ex_reg_rs_lsb_0__q)
    );
    wire [63:0] _node_325;
    assign _node_325 = bypass_mux_0;
    wire _node_326;
    EQ_UNSIGNED #(.width(2)) u_eq_4116 (
        .y(_node_326),
        .a(2'd1),
        .b(_ex_reg_rs_lsb_0__q)
    );
    wire [63:0] _node_327;
    MUX_UNSIGNED #(.width(64)) u_mux_4117 (
        .y(_node_327),
        .sel(_node_326),
        .a(bypass_mux_1),
        .b(_node_325)
    );
    wire _node_328;
    EQ_UNSIGNED #(.width(2)) u_eq_4118 (
        .y(_node_328),
        .a(2'd2),
        .b(_ex_reg_rs_lsb_0__q)
    );
    wire [63:0] _node_329;
    MUX_UNSIGNED #(.width(64)) u_mux_4119 (
        .y(_node_329),
        .sel(_node_328),
        .a(bypass_mux_2),
        .b(_node_327)
    );
    wire _node_330;
    EQ_UNSIGNED #(.width(2)) u_eq_4120 (
        .y(_node_330),
        .a(2'd3),
        .b(_ex_reg_rs_lsb_0__q)
    );
    wire [63:0] _node_331;
    MUX_UNSIGNED #(.width(64)) u_mux_4121 (
        .y(_node_331),
        .sel(_node_330),
        .a(bypass_mux_3),
        .b(_node_329)
    );
    wire [63:0] ex_rs_0;
    MUX_UNSIGNED #(.width(64)) u_mux_4122 (
        .y(ex_rs_0),
        .sel(_ex_reg_rs_bypass_0__q),
        .a(_node_331),
        .b(_T_3605)
    );
    wire [63:0] _T_3607;
    CAT #(.width_a(62), .width_b(2)) cat_4123 (
        .y(_T_3607),
        .a(_ex_reg_rs_msb_1__q),
        .b(_ex_reg_rs_lsb_1__q)
    );
    wire _node_332;
    EQ_UNSIGNED #(.width(2)) u_eq_4124 (
        .y(_node_332),
        .a(2'd0),
        .b(_ex_reg_rs_lsb_1__q)
    );
    wire [63:0] _node_333;
    assign _node_333 = bypass_mux_0;
    wire _node_334;
    EQ_UNSIGNED #(.width(2)) u_eq_4125 (
        .y(_node_334),
        .a(2'd1),
        .b(_ex_reg_rs_lsb_1__q)
    );
    wire [63:0] _node_335;
    MUX_UNSIGNED #(.width(64)) u_mux_4126 (
        .y(_node_335),
        .sel(_node_334),
        .a(bypass_mux_1),
        .b(_node_333)
    );
    wire _node_336;
    EQ_UNSIGNED #(.width(2)) u_eq_4127 (
        .y(_node_336),
        .a(2'd2),
        .b(_ex_reg_rs_lsb_1__q)
    );
    wire [63:0] _node_337;
    MUX_UNSIGNED #(.width(64)) u_mux_4128 (
        .y(_node_337),
        .sel(_node_336),
        .a(bypass_mux_2),
        .b(_node_335)
    );
    wire _node_338;
    EQ_UNSIGNED #(.width(2)) u_eq_4129 (
        .y(_node_338),
        .a(2'd3),
        .b(_ex_reg_rs_lsb_1__q)
    );
    wire [63:0] _node_339;
    MUX_UNSIGNED #(.width(64)) u_mux_4130 (
        .y(_node_339),
        .sel(_node_338),
        .a(bypass_mux_3),
        .b(_node_337)
    );
    wire [63:0] ex_rs_1;
    MUX_UNSIGNED #(.width(64)) u_mux_4131 (
        .y(ex_rs_1),
        .sel(_ex_reg_rs_bypass_1__q),
        .a(_node_339),
        .b(_T_3607)
    );
    wire _T_3609;
    EQ_UNSIGNED #(.width(3)) u_eq_4132 (
        .y(_T_3609),
        .a(_ex_ctrl_sel_imm__q),
        .b(3'h5)
    );
    wire _T_3611;
    BITS #(.width(32), .high(31), .low(31)) bits_4133 (
        .y(_T_3611),
        .in(_ex_reg_inst__q)
    );
    wire _T_3612;
    ASSINT #(.width(1)) assint_4134 (
        .y(_T_3612),
        .in(_T_3611)
    );
    wire _T_3613;
    MUX_SIGNED #(.width(1)) s_mux_4135 (
        .y(_T_3613),
        .sel(_T_3609),
        .a(1'sh0),
        .b(_T_3612)
    );
    wire _T_3615;
    EQ_UNSIGNED #(.width(3)) u_eq_4136 (
        .y(_T_3615),
        .a(_ex_ctrl_sel_imm__q),
        .b(3'h2)
    );
    wire [10:0] _T_3616;
    BITS #(.width(32), .high(30), .low(20)) bits_4137 (
        .y(_T_3616),
        .in(_ex_reg_inst__q)
    );
    wire [10:0] _T_3617;
    ASSINT #(.width(11)) assint_4138 (
        .y(_T_3617),
        .in(_T_3616)
    );
    wire [10:0] _T_3618;
    wire [10:0] _WTEMP_575;
    PAD_SIGNED #(.width(1), .n(11)) s_pad_4139 (
        .y(_WTEMP_575),
        .in(_T_3613)
    );
    MUX_SIGNED #(.width(11)) s_mux_4140 (
        .y(_T_3618),
        .sel(_T_3615),
        .a(_T_3617),
        .b(_WTEMP_575)
    );
    wire _T_3620;
    NEQ_UNSIGNED #(.width(3)) u_neq_4141 (
        .y(_T_3620),
        .a(_ex_ctrl_sel_imm__q),
        .b(3'h2)
    );
    wire _T_3622;
    NEQ_UNSIGNED #(.width(3)) u_neq_4142 (
        .y(_T_3622),
        .a(_ex_ctrl_sel_imm__q),
        .b(3'h3)
    );
    wire _T_3623;
    BITWISEAND #(.width(1)) bitwiseand_4143 (
        .y(_T_3623),
        .a(_T_3620),
        .b(_T_3622)
    );
    wire [7:0] _T_3624;
    BITS #(.width(32), .high(19), .low(12)) bits_4144 (
        .y(_T_3624),
        .in(_ex_reg_inst__q)
    );
    wire [7:0] _T_3625;
    ASSINT #(.width(8)) assint_4145 (
        .y(_T_3625),
        .in(_T_3624)
    );
    wire [7:0] _T_3626;
    wire [7:0] _WTEMP_576;
    PAD_SIGNED #(.width(1), .n(8)) s_pad_4146 (
        .y(_WTEMP_576),
        .in(_T_3613)
    );
    MUX_SIGNED #(.width(8)) s_mux_4147 (
        .y(_T_3626),
        .sel(_T_3623),
        .a(_WTEMP_576),
        .b(_T_3625)
    );
    wire _T_3628;
    EQ_UNSIGNED #(.width(3)) u_eq_4148 (
        .y(_T_3628),
        .a(_ex_ctrl_sel_imm__q),
        .b(3'h2)
    );
    wire _T_3630;
    EQ_UNSIGNED #(.width(3)) u_eq_4149 (
        .y(_T_3630),
        .a(_ex_ctrl_sel_imm__q),
        .b(3'h5)
    );
    wire _T_3631;
    BITWISEOR #(.width(1)) bitwiseor_4150 (
        .y(_T_3631),
        .a(_T_3628),
        .b(_T_3630)
    );
    wire _T_3634;
    EQ_UNSIGNED #(.width(3)) u_eq_4151 (
        .y(_T_3634),
        .a(_ex_ctrl_sel_imm__q),
        .b(3'h3)
    );
    wire _T_3635;
    BITS #(.width(32), .high(20), .low(20)) bits_4152 (
        .y(_T_3635),
        .in(_ex_reg_inst__q)
    );
    wire _T_3636;
    ASSINT #(.width(1)) assint_4153 (
        .y(_T_3636),
        .in(_T_3635)
    );
    wire _T_3638;
    EQ_UNSIGNED #(.width(3)) u_eq_4154 (
        .y(_T_3638),
        .a(_ex_ctrl_sel_imm__q),
        .b(3'h1)
    );
    wire _T_3639;
    BITS #(.width(32), .high(7), .low(7)) bits_4155 (
        .y(_T_3639),
        .in(_ex_reg_inst__q)
    );
    wire _T_3640;
    ASSINT #(.width(1)) assint_4156 (
        .y(_T_3640),
        .in(_T_3639)
    );
    wire _T_3641;
    MUX_SIGNED #(.width(1)) s_mux_4157 (
        .y(_T_3641),
        .sel(_T_3638),
        .a(_T_3640),
        .b(_T_3613)
    );
    wire _T_3642;
    MUX_SIGNED #(.width(1)) s_mux_4158 (
        .y(_T_3642),
        .sel(_T_3634),
        .a(_T_3636),
        .b(_T_3641)
    );
    wire _T_3643;
    MUX_SIGNED #(.width(1)) s_mux_4159 (
        .y(_T_3643),
        .sel(_T_3631),
        .a(1'sh0),
        .b(_T_3642)
    );
    wire _T_3645;
    EQ_UNSIGNED #(.width(3)) u_eq_4160 (
        .y(_T_3645),
        .a(_ex_ctrl_sel_imm__q),
        .b(3'h2)
    );
    wire _T_3647;
    EQ_UNSIGNED #(.width(3)) u_eq_4161 (
        .y(_T_3647),
        .a(_ex_ctrl_sel_imm__q),
        .b(3'h5)
    );
    wire _T_3648;
    BITWISEOR #(.width(1)) bitwiseor_4162 (
        .y(_T_3648),
        .a(_T_3645),
        .b(_T_3647)
    );
    wire [5:0] _T_3650;
    BITS #(.width(32), .high(30), .low(25)) bits_4163 (
        .y(_T_3650),
        .in(_ex_reg_inst__q)
    );
    wire [5:0] _T_3651;
    wire [5:0] _WTEMP_577;
    PAD_UNSIGNED #(.width(1), .n(6)) u_pad_4164 (
        .y(_WTEMP_577),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(6)) u_mux_4165 (
        .y(_T_3651),
        .sel(_T_3648),
        .a(_WTEMP_577),
        .b(_T_3650)
    );
    wire _T_3653;
    EQ_UNSIGNED #(.width(3)) u_eq_4166 (
        .y(_T_3653),
        .a(_ex_ctrl_sel_imm__q),
        .b(3'h2)
    );
    wire _T_3656;
    EQ_UNSIGNED #(.width(3)) u_eq_4167 (
        .y(_T_3656),
        .a(_ex_ctrl_sel_imm__q),
        .b(3'h0)
    );
    wire _T_3658;
    EQ_UNSIGNED #(.width(3)) u_eq_4168 (
        .y(_T_3658),
        .a(_ex_ctrl_sel_imm__q),
        .b(3'h1)
    );
    wire _T_3659;
    BITWISEOR #(.width(1)) bitwiseor_4169 (
        .y(_T_3659),
        .a(_T_3656),
        .b(_T_3658)
    );
    wire [3:0] _T_3660;
    BITS #(.width(32), .high(11), .low(8)) bits_4170 (
        .y(_T_3660),
        .in(_ex_reg_inst__q)
    );
    wire _T_3662;
    EQ_UNSIGNED #(.width(3)) u_eq_4171 (
        .y(_T_3662),
        .a(_ex_ctrl_sel_imm__q),
        .b(3'h5)
    );
    wire [3:0] _T_3663;
    BITS #(.width(32), .high(19), .low(16)) bits_4172 (
        .y(_T_3663),
        .in(_ex_reg_inst__q)
    );
    wire [3:0] _T_3664;
    BITS #(.width(32), .high(24), .low(21)) bits_4173 (
        .y(_T_3664),
        .in(_ex_reg_inst__q)
    );
    wire [3:0] _T_3665;
    MUX_UNSIGNED #(.width(4)) u_mux_4174 (
        .y(_T_3665),
        .sel(_T_3662),
        .a(_T_3663),
        .b(_T_3664)
    );
    wire [3:0] _T_3666;
    MUX_UNSIGNED #(.width(4)) u_mux_4175 (
        .y(_T_3666),
        .sel(_T_3659),
        .a(_T_3660),
        .b(_T_3665)
    );
    wire [3:0] _T_3667;
    wire [3:0] _WTEMP_578;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_4176 (
        .y(_WTEMP_578),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(4)) u_mux_4177 (
        .y(_T_3667),
        .sel(_T_3653),
        .a(_WTEMP_578),
        .b(_T_3666)
    );
    wire _T_3669;
    EQ_UNSIGNED #(.width(3)) u_eq_4178 (
        .y(_T_3669),
        .a(_ex_ctrl_sel_imm__q),
        .b(3'h0)
    );
    wire _T_3670;
    BITS #(.width(32), .high(7), .low(7)) bits_4179 (
        .y(_T_3670),
        .in(_ex_reg_inst__q)
    );
    wire _T_3672;
    EQ_UNSIGNED #(.width(3)) u_eq_4180 (
        .y(_T_3672),
        .a(_ex_ctrl_sel_imm__q),
        .b(3'h4)
    );
    wire _T_3673;
    BITS #(.width(32), .high(20), .low(20)) bits_4181 (
        .y(_T_3673),
        .in(_ex_reg_inst__q)
    );
    wire _T_3675;
    EQ_UNSIGNED #(.width(3)) u_eq_4182 (
        .y(_T_3675),
        .a(_ex_ctrl_sel_imm__q),
        .b(3'h5)
    );
    wire _T_3676;
    BITS #(.width(32), .high(15), .low(15)) bits_4183 (
        .y(_T_3676),
        .in(_ex_reg_inst__q)
    );
    wire _T_3678;
    MUX_UNSIGNED #(.width(1)) u_mux_4184 (
        .y(_T_3678),
        .sel(_T_3675),
        .a(_T_3676),
        .b(1'h0)
    );
    wire _T_3679;
    MUX_UNSIGNED #(.width(1)) u_mux_4185 (
        .y(_T_3679),
        .sel(_T_3672),
        .a(_T_3673),
        .b(_T_3678)
    );
    wire _T_3680;
    MUX_UNSIGNED #(.width(1)) u_mux_4186 (
        .y(_T_3680),
        .sel(_T_3669),
        .a(_T_3670),
        .b(_T_3679)
    );
    wire [9:0] _T_3681;
    CAT #(.width_a(6), .width_b(4)) cat_4187 (
        .y(_T_3681),
        .a(_T_3651),
        .b(_T_3667)
    );
    wire [10:0] _T_3682;
    CAT #(.width_a(10), .width_b(1)) cat_4188 (
        .y(_T_3682),
        .a(_T_3681),
        .b(_T_3680)
    );
    wire _T_3683;
    ASUINT #(.width(1)) asuint_4189 (
        .y(_T_3683),
        .in(_T_3643)
    );
    wire [7:0] _T_3684;
    ASUINT #(.width(8)) asuint_4190 (
        .y(_T_3684),
        .in(_T_3626)
    );
    wire [8:0] _T_3685;
    CAT #(.width_a(8), .width_b(1)) cat_4191 (
        .y(_T_3685),
        .a(_T_3684),
        .b(_T_3683)
    );
    wire [10:0] _T_3686;
    ASUINT #(.width(11)) asuint_4192 (
        .y(_T_3686),
        .in(_T_3618)
    );
    wire _T_3687;
    ASUINT #(.width(1)) asuint_4193 (
        .y(_T_3687),
        .in(_T_3613)
    );
    wire [11:0] _T_3688;
    CAT #(.width_a(1), .width_b(11)) cat_4194 (
        .y(_T_3688),
        .a(_T_3687),
        .b(_T_3686)
    );
    wire [20:0] _T_3689;
    CAT #(.width_a(12), .width_b(9)) cat_4195 (
        .y(_T_3689),
        .a(_T_3688),
        .b(_T_3685)
    );
    wire [31:0] _T_3690;
    CAT #(.width_a(21), .width_b(11)) cat_4196 (
        .y(_T_3690),
        .a(_T_3689),
        .b(_T_3682)
    );
    wire [31:0] ex_imm;
    ASSINT #(.width(32)) assint_4197 (
        .y(ex_imm),
        .in(_T_3690)
    );
    wire [63:0] _T_3693;
    ASSINT #(.width(64)) assint_4198 (
        .y(_T_3693),
        .in(ex_rs_0)
    );
    wire [39:0] _T_3695;
    ASSINT #(.width(40)) assint_4199 (
        .y(_T_3695),
        .in(_ex_reg_pc__q)
    );
    wire _T_3696;
    EQ_UNSIGNED #(.width(2)) u_eq_4200 (
        .y(_T_3696),
        .a(2'h2),
        .b(_ex_ctrl_sel_alu1__q)
    );
    wire [39:0] _T_3697;
    wire [39:0] _WTEMP_579;
    PAD_SIGNED #(.width(1), .n(40)) s_pad_4201 (
        .y(_WTEMP_579),
        .in(1'sh0)
    );
    MUX_SIGNED #(.width(40)) s_mux_4202 (
        .y(_T_3697),
        .sel(_T_3696),
        .a(_T_3695),
        .b(_WTEMP_579)
    );
    wire _T_3698;
    EQ_UNSIGNED #(.width(2)) u_eq_4203 (
        .y(_T_3698),
        .a(2'h1),
        .b(_ex_ctrl_sel_alu1__q)
    );
    wire [63:0] ex_op1;
    wire [63:0] _WTEMP_580;
    PAD_SIGNED #(.width(40), .n(64)) s_pad_4204 (
        .y(_WTEMP_580),
        .in(_T_3697)
    );
    MUX_SIGNED #(.width(64)) s_mux_4205 (
        .y(ex_op1),
        .sel(_T_3698),
        .a(_T_3693),
        .b(_WTEMP_580)
    );
    wire [63:0] _T_3701;
    ASSINT #(.width(64)) assint_4206 (
        .y(_T_3701),
        .in(ex_rs_1)
    );
    wire [3:0] _T_3706;
    wire [3:0] _WTEMP_581;
    PAD_SIGNED #(.width(3), .n(4)) s_pad_4207 (
        .y(_WTEMP_581),
        .in(3'sh2)
    );
    MUX_SIGNED #(.width(4)) s_mux_4208 (
        .y(_T_3706),
        .sel(_ex_reg_rvc__q),
        .a(_WTEMP_581),
        .b(4'sh4)
    );
    wire _T_3707;
    EQ_UNSIGNED #(.width(2)) u_eq_4209 (
        .y(_T_3707),
        .a(2'h1),
        .b(_ex_ctrl_sel_alu2__q)
    );
    wire [3:0] _T_3708;
    wire [3:0] _WTEMP_582;
    PAD_SIGNED #(.width(1), .n(4)) s_pad_4210 (
        .y(_WTEMP_582),
        .in(1'sh0)
    );
    MUX_SIGNED #(.width(4)) s_mux_4211 (
        .y(_T_3708),
        .sel(_T_3707),
        .a(_T_3706),
        .b(_WTEMP_582)
    );
    wire _T_3709;
    EQ_UNSIGNED #(.width(2)) u_eq_4212 (
        .y(_T_3709),
        .a(2'h3),
        .b(_ex_ctrl_sel_alu2__q)
    );
    wire [31:0] _T_3710;
    wire [31:0] _WTEMP_583;
    PAD_SIGNED #(.width(4), .n(32)) s_pad_4213 (
        .y(_WTEMP_583),
        .in(_T_3708)
    );
    MUX_SIGNED #(.width(32)) s_mux_4214 (
        .y(_T_3710),
        .sel(_T_3709),
        .a(ex_imm),
        .b(_WTEMP_583)
    );
    wire _T_3711;
    EQ_UNSIGNED #(.width(2)) u_eq_4215 (
        .y(_T_3711),
        .a(2'h2),
        .b(_ex_ctrl_sel_alu2__q)
    );
    wire [63:0] ex_op2;
    wire [63:0] _WTEMP_584;
    PAD_SIGNED #(.width(32), .n(64)) s_pad_4216 (
        .y(_WTEMP_584),
        .in(_T_3710)
    );
    MUX_SIGNED #(.width(64)) s_mux_4217 (
        .y(ex_op2),
        .sel(_T_3711),
        .a(_T_3701),
        .b(_WTEMP_584)
    );
    wire _alu__clock;
    wire _alu__reset;
    wire _alu__io_dw;
    wire [3:0] _alu__io_fn;
    wire [63:0] _alu__io_in2;
    wire [63:0] _alu__io_in1;
    wire [63:0] _alu__io_out;
    wire [63:0] _alu__io_adder_out;
    wire _alu__io_cmp_out;
    ALU alu (
        .clock(_alu__clock),
        .reset(_alu__reset),
        .io_dw(_alu__io_dw),
        .io_fn(_alu__io_fn),
        .io_in2(_alu__io_in2),
        .io_in1(_alu__io_in1),
        .io_out(_alu__io_out),
        .io_adder_out(_alu__io_adder_out),
        .io_cmp_out(_alu__io_cmp_out)
    );
    wire [63:0] _T_3712;
    ASUINT #(.width(64)) asuint_4405 (
        .y(_T_3712),
        .in(ex_op2)
    );
    wire [63:0] _T_3713;
    ASUINT #(.width(64)) asuint_4406 (
        .y(_T_3713),
        .in(ex_op1)
    );
    wire _div__clock;
    wire _div__reset;
    wire _div__io_req_ready;
    wire _div__io_req_valid;
    wire [3:0] _div__io_req_bits_fn;
    wire _div__io_req_bits_dw;
    wire [63:0] _div__io_req_bits_in1;
    wire [63:0] _div__io_req_bits_in2;
    wire [4:0] _div__io_req_bits_tag;
    wire _div__io_kill;
    wire _div__io_resp_ready;
    wire _div__io_resp_valid;
    wire [63:0] _div__io_resp_bits_data;
    wire [4:0] _div__io_resp_bits_tag;
    MulDiv div (
        .clock(_div__clock),
        .reset(_div__reset),
        .io_req_ready(_div__io_req_ready),
        .io_req_valid(_div__io_req_valid),
        .io_req_bits_fn(_div__io_req_bits_fn),
        .io_req_bits_dw(_div__io_req_bits_dw),
        .io_req_bits_in1(_div__io_req_bits_in1),
        .io_req_bits_in2(_div__io_req_bits_in2),
        .io_req_bits_tag(_div__io_req_bits_tag),
        .io_kill(_div__io_kill),
        .io_resp_ready(_div__io_resp_ready),
        .io_resp_valid(_div__io_resp_valid),
        .io_resp_bits_data(_div__io_resp_bits_data),
        .io_resp_bits_tag(_div__io_resp_bits_tag)
    );
    wire _T_3714;
    BITWISEAND #(.width(1)) bitwiseand_5018 (
        .y(_T_3714),
        .a(_ex_reg_valid__q),
        .b(_ex_ctrl_div__q)
    );
    wire _T_3716;
    EQ_UNSIGNED #(.width(1)) u_eq_5019 (
        .y(_T_3716),
        .a(ctrl_killd),
        .b(1'h0)
    );
    wire _T_3718;
    EQ_UNSIGNED #(.width(1)) u_eq_5020 (
        .y(_T_3718),
        .a(take_pc),
        .b(1'h0)
    );
    wire _T_3719;
    BITWISEAND #(.width(1)) bitwiseand_5021 (
        .y(_T_3719),
        .a(_T_3718),
        .b(_ibuf__io_inst_0_valid)
    );
    wire _T_3720;
    BITWISEAND #(.width(1)) bitwiseand_5022 (
        .y(_T_3720),
        .a(_T_3719),
        .b(_ibuf__io_inst_0_bits_replay)
    );
    wire _T_3722;
    EQ_UNSIGNED #(.width(1)) u_eq_5023 (
        .y(_T_3722),
        .a(ctrl_killd),
        .b(1'h0)
    );
    wire _T_3723;
    BITWISEAND #(.width(1)) bitwiseand_5024 (
        .y(_T_3723),
        .a(_T_3722),
        .b(id_xcpt)
    );
    wire _T_3725;
    EQ_UNSIGNED #(.width(1)) u_eq_5025 (
        .y(_T_3725),
        .a(take_pc),
        .b(1'h0)
    );
    wire _T_3726;
    BITWISEAND #(.width(1)) bitwiseand_5026 (
        .y(_T_3726),
        .a(_T_3725),
        .b(_ibuf__io_inst_0_valid)
    );
    wire _T_3727;
    BITWISEAND #(.width(1)) bitwiseand_5027 (
        .y(_T_3727),
        .a(_T_3726),
        .b(_csr__io_interrupt)
    );
    wire _T_3729;
    EQ_UNSIGNED #(.width(1)) u_eq_5028 (
        .y(_T_3729),
        .a(ctrl_killd),
        .b(1'h0)
    );
    wire _T_3735;
    EQ_UNSIGNED #(.width(1)) u_eq_5029 (
        .y(_T_3735),
        .a(_bpu__io_xcpt_if),
        .b(1'h0)
    );
    wire _T_3737;
    EQ_UNSIGNED #(.width(1)) u_eq_5030 (
        .y(_T_3737),
        .a(_ibuf__io_inst_0_bits_pf0),
        .b(1'h0)
    );
    wire _T_3738;
    BITWISEAND #(.width(1)) bitwiseand_5031 (
        .y(_T_3738),
        .a(_T_3735),
        .b(_T_3737)
    );
    wire _T_3739;
    BITWISEAND #(.width(1)) bitwiseand_5032 (
        .y(_T_3739),
        .a(_T_3738),
        .b(_ibuf__io_inst_0_bits_pf1)
    );
    wire [1:0] _node_364;
    MUX_UNSIGNED #(.width(2)) u_mux_5033 (
        .y(_node_364),
        .sel(_T_3739),
        .a(2'h1),
        .b(2'h0)
    );
    wire _node_365;
    MUX_UNSIGNED #(.width(1)) u_mux_5034 (
        .y(_node_365),
        .sel(_T_3739),
        .a(1'h1),
        .b(_ibuf__io_inst_0_bits_rvc)
    );
    wire _T_3742;
    BITWISEOR #(.width(1)) bitwiseor_5035 (
        .y(_T_3742),
        .a(id_ctrl_fence_i),
        .b(id_csr_flush)
    );
    wire _T_3743;
    BITWISEOR #(.width(1)) bitwiseor_5036 (
        .y(_T_3743),
        .a(_T_3742),
        .b(_csr__io_singleStep)
    );
    wire _T_3744;
    BITWISEAND #(.width(1)) bitwiseand_5037 (
        .y(_T_3744),
        .a(id_ctrl_jalr),
        .b(_csr__io_status_debug)
    );
    wire _T_3747;
    BITWISEOR #(.width(1)) bitwiseor_5038 (
        .y(_T_3747),
        .a(id_bypass_src_0_0),
        .b(id_bypass_src_0_1)
    );
    wire _T_3748;
    BITWISEOR #(.width(1)) bitwiseor_5039 (
        .y(_T_3748),
        .a(_T_3747),
        .b(id_bypass_src_0_2)
    );
    wire _T_3749;
    BITWISEOR #(.width(1)) bitwiseor_5040 (
        .y(_T_3749),
        .a(_T_3748),
        .b(id_bypass_src_0_3)
    );
    wire [1:0] _T_3754;
    MUX_UNSIGNED #(.width(2)) u_mux_5041 (
        .y(_T_3754),
        .sel(id_bypass_src_0_2),
        .a(2'h2),
        .b(2'h3)
    );
    wire [1:0] _T_3755;
    wire [1:0] _WTEMP_697;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_5042 (
        .y(_WTEMP_697),
        .in(1'h1)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_5043 (
        .y(_T_3755),
        .sel(id_bypass_src_0_1),
        .a(_WTEMP_697),
        .b(_T_3754)
    );
    wire [1:0] _T_3756;
    wire [1:0] _WTEMP_698;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_5044 (
        .y(_WTEMP_698),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_5045 (
        .y(_T_3756),
        .sel(id_bypass_src_0_0),
        .a(_WTEMP_698),
        .b(_T_3755)
    );
    wire _T_3758;
    EQ_UNSIGNED #(.width(1)) u_eq_5046 (
        .y(_T_3758),
        .a(_T_3749),
        .b(1'h0)
    );
    wire _T_3759;
    BITWISEAND #(.width(1)) bitwiseand_5047 (
        .y(_T_3759),
        .a(id_ctrl_rxs1),
        .b(_T_3758)
    );
    wire [1:0] _T_3760;
    BITS #(.width(64), .high(1), .low(0)) bits_5048 (
        .y(_T_3760),
        .in(id_rs_0)
    );
    wire [61:0] _T_3761;
    SHR_UNSIGNED #(.width(64), .n(2)) u_shr_5049 (
        .y(_T_3761),
        .in(id_rs_0)
    );
    wire _T_3762;
    BITWISEOR #(.width(1)) bitwiseor_5050 (
        .y(_T_3762),
        .a(id_bypass_src_1_0),
        .b(id_bypass_src_1_1)
    );
    wire _T_3763;
    BITWISEOR #(.width(1)) bitwiseor_5051 (
        .y(_T_3763),
        .a(_T_3762),
        .b(id_bypass_src_1_2)
    );
    wire _T_3764;
    BITWISEOR #(.width(1)) bitwiseor_5052 (
        .y(_T_3764),
        .a(_T_3763),
        .b(id_bypass_src_1_3)
    );
    wire [1:0] _T_3769;
    MUX_UNSIGNED #(.width(2)) u_mux_5053 (
        .y(_T_3769),
        .sel(id_bypass_src_1_2),
        .a(2'h2),
        .b(2'h3)
    );
    wire [1:0] _T_3770;
    wire [1:0] _WTEMP_699;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_5054 (
        .y(_WTEMP_699),
        .in(1'h1)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_5055 (
        .y(_T_3770),
        .sel(id_bypass_src_1_1),
        .a(_WTEMP_699),
        .b(_T_3769)
    );
    wire [1:0] _T_3771;
    wire [1:0] _WTEMP_700;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_5056 (
        .y(_WTEMP_700),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_5057 (
        .y(_T_3771),
        .sel(id_bypass_src_1_0),
        .a(_WTEMP_700),
        .b(_T_3770)
    );
    wire _T_3773;
    EQ_UNSIGNED #(.width(1)) u_eq_5058 (
        .y(_T_3773),
        .a(_T_3764),
        .b(1'h0)
    );
    wire _T_3774;
    BITWISEAND #(.width(1)) bitwiseand_5059 (
        .y(_T_3774),
        .a(id_ctrl_rxs2),
        .b(_T_3773)
    );
    wire [1:0] _T_3775;
    BITS #(.width(64), .high(1), .low(0)) bits_5060 (
        .y(_T_3775),
        .in(id_rs_1)
    );
    wire [61:0] _T_3776;
    SHR_UNSIGNED #(.width(64), .n(2)) u_shr_5061 (
        .y(_T_3776),
        .in(id_rs_1)
    );
    wire _node_366;
    MUX_UNSIGNED #(.width(1)) u_mux_5062 (
        .y(_node_366),
        .sel(id_xcpt),
        .a(1'h1),
        .b(id_ctrl_alu_dw)
    );
    wire [3:0] _node_367;
    wire [3:0] _WTEMP_701;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_5063 (
        .y(_WTEMP_701),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(4)) u_mux_5064 (
        .y(_node_367),
        .sel(id_xcpt),
        .a(_WTEMP_701),
        .b(id_ctrl_alu_fn)
    );
    wire _node_368;
    MUX_UNSIGNED #(.width(1)) u_mux_5065 (
        .y(_node_368),
        .sel(_T_3744),
        .a(1'h1),
        .b(id_ctrl_fence_i)
    );
    wire [1:0] _node_369;
    MUX_UNSIGNED #(.width(2)) u_mux_5066 (
        .y(_node_369),
        .sel(id_xcpt),
        .a(2'h2),
        .b(id_ctrl_sel_alu1)
    );
    wire [1:0] _node_370;
    MUX_UNSIGNED #(.width(2)) u_mux_5067 (
        .y(_node_370),
        .sel(id_xcpt),
        .a(_node_364),
        .b(id_ctrl_sel_alu2)
    );
    wire _node_371;
    MUX_UNSIGNED #(.width(1)) u_mux_5068 (
        .y(_node_371),
        .sel(_T_3744),
        .a(1'h1),
        .b(_T_3743)
    );
    wire [1:0] _node_372;
    MUX_UNSIGNED #(.width(2)) u_mux_5069 (
        .y(_node_372),
        .sel(_T_3759),
        .a(_T_3760),
        .b(_T_3756)
    );
    wire [1:0] _node_373;
    MUX_UNSIGNED #(.width(2)) u_mux_5070 (
        .y(_node_373),
        .sel(_T_3774),
        .a(_T_3775),
        .b(_T_3771)
    );
    wire [61:0] _node_374;
    MUX_UNSIGNED #(.width(62)) u_mux_5071 (
        .y(_node_374),
        .sel(_T_3759),
        .a(_T_3761),
        .b(_ex_reg_rs_msb_0__q)
    );
    wire [61:0] _node_375;
    MUX_UNSIGNED #(.width(62)) u_mux_5072 (
        .y(_node_375),
        .sel(_T_3774),
        .a(_T_3776),
        .b(_ex_reg_rs_msb_1__q)
    );
    wire _node_376;
    MUX_UNSIGNED #(.width(1)) u_mux_5073 (
        .y(_node_376),
        .sel(id_xcpt),
        .a(_node_365),
        .b(_ibuf__io_inst_0_bits_rvc)
    );
    wire _T_3778;
    EQ_UNSIGNED #(.width(1)) u_eq_5074 (
        .y(_T_3778),
        .a(ctrl_killd),
        .b(1'h0)
    );
    wire _T_3779;
    BITWISEOR #(.width(1)) bitwiseor_5075 (
        .y(_T_3779),
        .a(_T_3778),
        .b(_csr__io_interrupt)
    );
    wire _T_3780;
    BITWISEOR #(.width(1)) bitwiseor_5076 (
        .y(_T_3780),
        .a(_T_3779),
        .b(_ibuf__io_inst_0_bits_replay)
    );
    wire _T_3781;
    BITWISEOR #(.width(1)) bitwiseor_5077 (
        .y(_T_3781),
        .a(_ex_reg_valid__q),
        .b(_ex_reg_replay__q)
    );
    wire ex_pc_valid;
    BITWISEOR #(.width(1)) bitwiseor_5078 (
        .y(ex_pc_valid),
        .a(_T_3781),
        .b(_ex_reg_xcpt_interrupt__q)
    );
    wire _T_3783;
    EQ_UNSIGNED #(.width(1)) u_eq_5079 (
        .y(_T_3783),
        .a(io_dmem_resp_valid),
        .b(1'h0)
    );
    wire wb_dcache_miss;
    BITWISEAND #(.width(1)) bitwiseand_5080 (
        .y(wb_dcache_miss),
        .a(_wb_ctrl_mem__q),
        .b(_T_3783)
    );
    wire _T_3785;
    EQ_UNSIGNED #(.width(1)) u_eq_5081 (
        .y(_T_3785),
        .a(io_dmem_req_ready),
        .b(1'h0)
    );
    wire _T_3786;
    BITWISEAND #(.width(1)) bitwiseand_5082 (
        .y(_T_3786),
        .a(_ex_ctrl_mem__q),
        .b(_T_3785)
    );
    wire _T_3788;
    EQ_UNSIGNED #(.width(1)) u_eq_5083 (
        .y(_T_3788),
        .a(_div__io_req_ready),
        .b(1'h0)
    );
    wire _T_3789;
    BITWISEAND #(.width(1)) bitwiseand_5084 (
        .y(_T_3789),
        .a(_ex_ctrl_div__q),
        .b(_T_3788)
    );
    wire replay_ex_structural;
    BITWISEOR #(.width(1)) bitwiseor_5085 (
        .y(replay_ex_structural),
        .a(_T_3786),
        .b(_T_3789)
    );
    wire replay_ex_load_use;
    BITWISEAND #(.width(1)) bitwiseand_5086 (
        .y(replay_ex_load_use),
        .a(wb_dcache_miss),
        .b(_ex_reg_load_use__q)
    );
    wire _T_3790;
    BITWISEOR #(.width(1)) bitwiseor_5087 (
        .y(_T_3790),
        .a(replay_ex_structural),
        .b(replay_ex_load_use)
    );
    wire _T_3791;
    BITWISEAND #(.width(1)) bitwiseand_5088 (
        .y(_T_3791),
        .a(_ex_reg_valid__q),
        .b(_T_3790)
    );
    wire replay_ex;
    BITWISEOR #(.width(1)) bitwiseor_5089 (
        .y(replay_ex),
        .a(_ex_reg_replay__q),
        .b(_T_3791)
    );
    wire _T_3792;
    BITWISEOR #(.width(1)) bitwiseor_5090 (
        .y(_T_3792),
        .a(take_pc_mem_wb),
        .b(replay_ex)
    );
    wire _T_3794;
    EQ_UNSIGNED #(.width(1)) u_eq_5091 (
        .y(_T_3794),
        .a(_ex_reg_valid__q),
        .b(1'h0)
    );
    wire ctrl_killx;
    BITWISEOR #(.width(1)) bitwiseor_5092 (
        .y(ctrl_killx),
        .a(_T_3792),
        .b(_T_3794)
    );
    wire _T_3796;
    wire [4:0] _WTEMP_702;
    PAD_UNSIGNED #(.width(3), .n(5)) u_pad_5093 (
        .y(_WTEMP_702),
        .in(3'h7)
    );
    EQ_UNSIGNED #(.width(5)) u_eq_5094 (
        .y(_T_3796),
        .a(_ex_ctrl_mem_cmd__q),
        .b(_WTEMP_702)
    );
    wire [2:0] _T_3803_0;
    wire [2:0] _T_3803_1;
    wire [2:0] _T_3803_2;
    wire [2:0] _T_3803_3;
    wire _T_3810;
    EQ_UNSIGNED #(.width(3)) u_eq_5095 (
        .y(_T_3810),
        .a(_T_3803_0),
        .b(_ex_ctrl_mem_type__q)
    );
    wire _T_3811;
    EQ_UNSIGNED #(.width(3)) u_eq_5096 (
        .y(_T_3811),
        .a(_T_3803_1),
        .b(_ex_ctrl_mem_type__q)
    );
    wire _T_3812;
    EQ_UNSIGNED #(.width(3)) u_eq_5097 (
        .y(_T_3812),
        .a(_T_3803_2),
        .b(_ex_ctrl_mem_type__q)
    );
    wire _T_3813;
    EQ_UNSIGNED #(.width(3)) u_eq_5098 (
        .y(_T_3813),
        .a(_T_3803_3),
        .b(_ex_ctrl_mem_type__q)
    );
    wire _T_3815;
    BITWISEOR #(.width(1)) bitwiseor_5099 (
        .y(_T_3815),
        .a(1'h0),
        .b(_T_3810)
    );
    wire _T_3816;
    BITWISEOR #(.width(1)) bitwiseor_5100 (
        .y(_T_3816),
        .a(_T_3815),
        .b(_T_3811)
    );
    wire _T_3817;
    BITWISEOR #(.width(1)) bitwiseor_5101 (
        .y(_T_3817),
        .a(_T_3816),
        .b(_T_3812)
    );
    wire _T_3818;
    BITWISEOR #(.width(1)) bitwiseor_5102 (
        .y(_T_3818),
        .a(_T_3817),
        .b(_T_3813)
    );
    wire ex_slow_bypass;
    BITWISEOR #(.width(1)) bitwiseor_5103 (
        .y(ex_slow_bypass),
        .a(_T_3796),
        .b(_T_3818)
    );
    wire ex_xcpt;
    BITWISEOR #(.width(1)) bitwiseor_5104 (
        .y(ex_xcpt),
        .a(_ex_reg_xcpt_interrupt__q),
        .b(_ex_reg_xcpt__q)
    );
    wire _T_3819;
    BITWISEOR #(.width(1)) bitwiseor_5105 (
        .y(_T_3819),
        .a(_mem_reg_valid__q),
        .b(_mem_reg_replay__q)
    );
    wire mem_pc_valid;
    BITWISEOR #(.width(1)) bitwiseor_5106 (
        .y(mem_pc_valid),
        .a(_T_3819),
        .b(_mem_reg_xcpt_interrupt__q)
    );
    wire mem_br_taken;
    BITS #(.width(64), .high(0), .low(0)) bits_5107 (
        .y(mem_br_taken),
        .in(_mem_reg_wdata__q)
    );
    wire [39:0] _T_3820;
    ASSINT #(.width(40)) assint_5108 (
        .y(_T_3820),
        .in(_mem_reg_pc__q)
    );
    wire _T_3821;
    BITWISEAND #(.width(1)) bitwiseand_5109 (
        .y(_T_3821),
        .a(_mem_ctrl_branch__q),
        .b(mem_br_taken)
    );
    wire _T_3824;
    assign _T_3824 = 1'h0;
    wire _T_3826;
    BITS #(.width(32), .high(31), .low(31)) bits_5110 (
        .y(_T_3826),
        .in(_mem_reg_inst__q)
    );
    wire _T_3827;
    ASSINT #(.width(1)) assint_5111 (
        .y(_T_3827),
        .in(_T_3826)
    );
    wire _T_3828;
    assign _T_3828 = _T_3827;
    wire _T_3830;
    assign _T_3830 = 1'h0;
    wire [10:0] _T_3831;
    BITS #(.width(32), .high(30), .low(20)) bits_5112 (
        .y(_T_3831),
        .in(_mem_reg_inst__q)
    );
    wire [10:0] _T_3832;
    ASSINT #(.width(11)) assint_5113 (
        .y(_T_3832),
        .in(_T_3831)
    );
    wire _T_3833;
    assign _T_3833 = _T_3828;
    wire _T_3835;
    assign _T_3835 = 1'h1;
    wire _T_3837;
    assign _T_3837 = 1'h1;
    wire _T_3838;
    assign _T_3838 = 1'h1;
    wire [7:0] _T_3839;
    BITS #(.width(32), .high(19), .low(12)) bits_5114 (
        .y(_T_3839),
        .in(_mem_reg_inst__q)
    );
    wire [7:0] _T_3840;
    ASSINT #(.width(8)) assint_5115 (
        .y(_T_3840),
        .in(_T_3839)
    );
    wire _T_3841;
    assign _T_3841 = _T_3828;
    wire _T_3843;
    assign _T_3843 = 1'h0;
    wire _T_3845;
    assign _T_3845 = 1'h0;
    wire _T_3846;
    assign _T_3846 = 1'h0;
    wire _T_3849;
    assign _T_3849 = 1'h0;
    wire _T_3850;
    BITS #(.width(32), .high(20), .low(20)) bits_5116 (
        .y(_T_3850),
        .in(_mem_reg_inst__q)
    );
    wire _T_3851;
    ASSINT #(.width(1)) assint_5117 (
        .y(_T_3851),
        .in(_T_3850)
    );
    wire _T_3853;
    assign _T_3853 = 1'h1;
    wire _T_3854;
    BITS #(.width(32), .high(7), .low(7)) bits_5118 (
        .y(_T_3854),
        .in(_mem_reg_inst__q)
    );
    wire _T_3855;
    ASSINT #(.width(1)) assint_5119 (
        .y(_T_3855),
        .in(_T_3854)
    );
    wire _T_3856;
    assign _T_3856 = _T_3855;
    wire _T_3857;
    assign _T_3857 = _T_3856;
    wire _T_3858;
    assign _T_3858 = _T_3857;
    wire _T_3860;
    assign _T_3860 = 1'h0;
    wire _T_3862;
    assign _T_3862 = 1'h0;
    wire _T_3863;
    assign _T_3863 = 1'h0;
    wire [5:0] _T_3865;
    BITS #(.width(32), .high(30), .low(25)) bits_5120 (
        .y(_T_3865),
        .in(_mem_reg_inst__q)
    );
    wire [5:0] _T_3866;
    assign _T_3866 = _T_3865;
    wire _T_3868;
    assign _T_3868 = 1'h0;
    wire _T_3871;
    assign _T_3871 = 1'h0;
    wire _T_3873;
    assign _T_3873 = 1'h1;
    wire _T_3874;
    assign _T_3874 = 1'h1;
    wire [3:0] _T_3875;
    BITS #(.width(32), .high(11), .low(8)) bits_5121 (
        .y(_T_3875),
        .in(_mem_reg_inst__q)
    );
    wire _T_3877;
    assign _T_3877 = 1'h0;
    wire [3:0] _T_3878;
    BITS #(.width(32), .high(19), .low(16)) bits_5122 (
        .y(_T_3878),
        .in(_mem_reg_inst__q)
    );
    wire [3:0] _T_3879;
    BITS #(.width(32), .high(24), .low(21)) bits_5123 (
        .y(_T_3879),
        .in(_mem_reg_inst__q)
    );
    wire [3:0] _T_3880;
    assign _T_3880 = _T_3879;
    wire [3:0] _T_3881;
    assign _T_3881 = _T_3875;
    wire [3:0] _T_3882;
    assign _T_3882 = _T_3881;
    wire _T_3884;
    assign _T_3884 = 1'h0;
    wire _T_3885;
    BITS #(.width(32), .high(7), .low(7)) bits_5124 (
        .y(_T_3885),
        .in(_mem_reg_inst__q)
    );
    wire _T_3887;
    assign _T_3887 = 1'h0;
    wire _T_3888;
    BITS #(.width(32), .high(20), .low(20)) bits_5125 (
        .y(_T_3888),
        .in(_mem_reg_inst__q)
    );
    wire _T_3890;
    assign _T_3890 = 1'h0;
    wire _T_3891;
    BITS #(.width(32), .high(15), .low(15)) bits_5126 (
        .y(_T_3891),
        .in(_mem_reg_inst__q)
    );
    wire _T_3893;
    assign _T_3893 = 1'h0;
    wire _T_3894;
    assign _T_3894 = 1'h0;
    wire _T_3895;
    assign _T_3895 = 1'h0;
    wire [9:0] _T_3896;
    CAT #(.width_a(6), .width_b(4)) cat_5127 (
        .y(_T_3896),
        .a(_T_3866),
        .b(_T_3882)
    );
    wire [10:0] _T_3897;
    CAT #(.width_a(10), .width_b(1)) cat_5128 (
        .y(_T_3897),
        .a(_T_3896),
        .b(_T_3895)
    );
    wire _T_3898;
    ASUINT #(.width(1)) asuint_5129 (
        .y(_T_3898),
        .in(_T_3858)
    );
    wire _T_3899;
    ASUINT #(.width(1)) asuint_5130 (
        .y(_T_3899),
        .in(_T_3841)
    );
    wire [1:0] _T_3900;
    CAT #(.width_a(1), .width_b(1)) cat_5131 (
        .y(_T_3900),
        .a(_T_3899),
        .b(_T_3898)
    );
    wire _T_3901;
    ASUINT #(.width(1)) asuint_5132 (
        .y(_T_3901),
        .in(_T_3833)
    );
    wire _T_3902;
    ASUINT #(.width(1)) asuint_5133 (
        .y(_T_3902),
        .in(_T_3828)
    );
    wire [1:0] _T_3903;
    CAT #(.width_a(1), .width_b(1)) cat_5134 (
        .y(_T_3903),
        .a(_T_3902),
        .b(_T_3901)
    );
    wire [3:0] _T_3904;
    CAT #(.width_a(2), .width_b(2)) cat_5135 (
        .y(_T_3904),
        .a(_T_3903),
        .b(_T_3900)
    );
    wire [14:0] _T_3905;
    CAT #(.width_a(4), .width_b(11)) cat_5136 (
        .y(_T_3905),
        .a(_T_3904),
        .b(_T_3897)
    );
    wire [14:0] _T_3906;
    ASSINT #(.width(15)) assint_5137 (
        .y(_T_3906),
        .in(_T_3905)
    );
    wire _T_3908;
    BITWISEAND #(.width(1)) bitwiseand_5138 (
        .y(_T_3908),
        .a(1'h1),
        .b(_mem_ctrl_jal__q)
    );
    wire _T_3911;
    assign _T_3911 = 1'h0;
    wire _T_3913;
    BITS #(.width(32), .high(31), .low(31)) bits_5139 (
        .y(_T_3913),
        .in(_mem_reg_inst__q)
    );
    wire _T_3914;
    ASSINT #(.width(1)) assint_5140 (
        .y(_T_3914),
        .in(_T_3913)
    );
    wire _T_3915;
    assign _T_3915 = _T_3914;
    wire _T_3917;
    assign _T_3917 = 1'h0;
    wire [10:0] _T_3918;
    BITS #(.width(32), .high(30), .low(20)) bits_5141 (
        .y(_T_3918),
        .in(_mem_reg_inst__q)
    );
    wire [10:0] _T_3919;
    ASSINT #(.width(11)) assint_5142 (
        .y(_T_3919),
        .in(_T_3918)
    );
    wire _T_3920;
    assign _T_3920 = _T_3915;
    wire _T_3922;
    assign _T_3922 = 1'h1;
    wire _T_3924;
    assign _T_3924 = 1'h0;
    wire _T_3925;
    assign _T_3925 = 1'h0;
    wire [7:0] _T_3926;
    BITS #(.width(32), .high(19), .low(12)) bits_5143 (
        .y(_T_3926),
        .in(_mem_reg_inst__q)
    );
    wire [7:0] _T_3927;
    ASSINT #(.width(8)) assint_5144 (
        .y(_T_3927),
        .in(_T_3926)
    );
    wire [7:0] _T_3928;
    assign _T_3928 = _T_3927;
    wire _T_3930;
    assign _T_3930 = 1'h0;
    wire _T_3932;
    assign _T_3932 = 1'h0;
    wire _T_3933;
    assign _T_3933 = 1'h0;
    wire _T_3936;
    assign _T_3936 = 1'h1;
    wire _T_3937;
    BITS #(.width(32), .high(20), .low(20)) bits_5145 (
        .y(_T_3937),
        .in(_mem_reg_inst__q)
    );
    wire _T_3938;
    ASSINT #(.width(1)) assint_5146 (
        .y(_T_3938),
        .in(_T_3937)
    );
    wire _T_3940;
    assign _T_3940 = 1'h0;
    wire _T_3941;
    BITS #(.width(32), .high(7), .low(7)) bits_5147 (
        .y(_T_3941),
        .in(_mem_reg_inst__q)
    );
    wire _T_3942;
    ASSINT #(.width(1)) assint_5148 (
        .y(_T_3942),
        .in(_T_3941)
    );
    wire _T_3943;
    assign _T_3943 = _T_3915;
    wire _T_3944;
    assign _T_3944 = _T_3938;
    wire _T_3945;
    assign _T_3945 = _T_3944;
    wire _T_3947;
    assign _T_3947 = 1'h0;
    wire _T_3949;
    assign _T_3949 = 1'h0;
    wire _T_3950;
    assign _T_3950 = 1'h0;
    wire [5:0] _T_3952;
    BITS #(.width(32), .high(30), .low(25)) bits_5149 (
        .y(_T_3952),
        .in(_mem_reg_inst__q)
    );
    wire [5:0] _T_3953;
    assign _T_3953 = _T_3952;
    wire _T_3955;
    assign _T_3955 = 1'h0;
    wire _T_3958;
    assign _T_3958 = 1'h0;
    wire _T_3960;
    assign _T_3960 = 1'h0;
    wire _T_3961;
    assign _T_3961 = 1'h0;
    wire [3:0] _T_3962;
    BITS #(.width(32), .high(11), .low(8)) bits_5150 (
        .y(_T_3962),
        .in(_mem_reg_inst__q)
    );
    wire _T_3964;
    assign _T_3964 = 1'h0;
    wire [3:0] _T_3965;
    BITS #(.width(32), .high(19), .low(16)) bits_5151 (
        .y(_T_3965),
        .in(_mem_reg_inst__q)
    );
    wire [3:0] _T_3966;
    BITS #(.width(32), .high(24), .low(21)) bits_5152 (
        .y(_T_3966),
        .in(_mem_reg_inst__q)
    );
    wire [3:0] _T_3967;
    assign _T_3967 = _T_3966;
    wire [3:0] _T_3968;
    assign _T_3968 = _T_3967;
    wire [3:0] _T_3969;
    assign _T_3969 = _T_3968;
    wire _T_3971;
    assign _T_3971 = 1'h0;
    wire _T_3972;
    BITS #(.width(32), .high(7), .low(7)) bits_5153 (
        .y(_T_3972),
        .in(_mem_reg_inst__q)
    );
    wire _T_3974;
    assign _T_3974 = 1'h0;
    wire _T_3975;
    BITS #(.width(32), .high(20), .low(20)) bits_5154 (
        .y(_T_3975),
        .in(_mem_reg_inst__q)
    );
    wire _T_3977;
    assign _T_3977 = 1'h0;
    wire _T_3978;
    BITS #(.width(32), .high(15), .low(15)) bits_5155 (
        .y(_T_3978),
        .in(_mem_reg_inst__q)
    );
    wire _T_3980;
    assign _T_3980 = 1'h0;
    wire _T_3981;
    assign _T_3981 = 1'h0;
    wire _T_3982;
    assign _T_3982 = 1'h0;
    wire [9:0] _T_3983;
    CAT #(.width_a(6), .width_b(4)) cat_5156 (
        .y(_T_3983),
        .a(_T_3953),
        .b(_T_3969)
    );
    wire [10:0] _T_3984;
    CAT #(.width_a(10), .width_b(1)) cat_5157 (
        .y(_T_3984),
        .a(_T_3983),
        .b(_T_3982)
    );
    wire _T_3985;
    ASUINT #(.width(1)) asuint_5158 (
        .y(_T_3985),
        .in(_T_3945)
    );
    wire [7:0] _T_3986;
    ASUINT #(.width(8)) asuint_5159 (
        .y(_T_3986),
        .in(_T_3928)
    );
    wire [8:0] _T_3987;
    CAT #(.width_a(8), .width_b(1)) cat_5160 (
        .y(_T_3987),
        .a(_T_3986),
        .b(_T_3985)
    );
    wire _T_3988;
    ASUINT #(.width(1)) asuint_5161 (
        .y(_T_3988),
        .in(_T_3920)
    );
    wire _T_3989;
    ASUINT #(.width(1)) asuint_5162 (
        .y(_T_3989),
        .in(_T_3915)
    );
    wire [1:0] _T_3990;
    CAT #(.width_a(1), .width_b(1)) cat_5163 (
        .y(_T_3990),
        .a(_T_3989),
        .b(_T_3988)
    );
    wire [10:0] _T_3991;
    CAT #(.width_a(2), .width_b(9)) cat_5164 (
        .y(_T_3991),
        .a(_T_3990),
        .b(_T_3987)
    );
    wire [21:0] _T_3992;
    CAT #(.width_a(11), .width_b(11)) cat_5165 (
        .y(_T_3992),
        .a(_T_3991),
        .b(_T_3984)
    );
    wire [21:0] _T_3993;
    ASSINT #(.width(22)) assint_5166 (
        .y(_T_3993),
        .in(_T_3992)
    );
    wire [3:0] _T_3996;
    wire [3:0] _WTEMP_703;
    PAD_SIGNED #(.width(3), .n(4)) s_pad_5167 (
        .y(_WTEMP_703),
        .in(3'sh2)
    );
    MUX_SIGNED #(.width(4)) s_mux_5168 (
        .y(_T_3996),
        .sel(_mem_reg_rvc__q),
        .a(_WTEMP_703),
        .b(4'sh4)
    );
    wire [21:0] _T_3997;
    wire [21:0] _WTEMP_704;
    PAD_SIGNED #(.width(4), .n(22)) s_pad_5169 (
        .y(_WTEMP_704),
        .in(_T_3996)
    );
    MUX_SIGNED #(.width(22)) s_mux_5170 (
        .y(_T_3997),
        .sel(_T_3908),
        .a(_T_3993),
        .b(_WTEMP_704)
    );
    wire [21:0] _T_3998;
    wire [21:0] _WTEMP_705;
    PAD_SIGNED #(.width(15), .n(22)) s_pad_5171 (
        .y(_WTEMP_705),
        .in(_T_3906)
    );
    MUX_SIGNED #(.width(22)) s_mux_5172 (
        .y(_T_3998),
        .sel(_T_3821),
        .a(_WTEMP_705),
        .b(_T_3997)
    );
    wire [40:0] _T_3999;
    wire [39:0] _WTEMP_706;
    PAD_SIGNED #(.width(22), .n(40)) s_pad_5173 (
        .y(_WTEMP_706),
        .in(_T_3998)
    );
    ADD_SIGNED #(.width(40)) s_add_5174 (
        .y(_T_3999),
        .a(_T_3820),
        .b(_WTEMP_706)
    );
    wire [39:0] _T_4000;
    TAIL #(.width(41), .n(1)) tail_5175 (
        .y(_T_4000),
        .in(_T_3999)
    );
    wire [39:0] mem_br_target;
    ASSINT #(.width(40)) assint_5176 (
        .y(mem_br_target),
        .in(_T_4000)
    );
    wire [25:0] _T_4001;
    SHR_UNSIGNED #(.width(64), .n(38)) u_shr_5177 (
        .y(_T_4001),
        .in(_mem_reg_wdata__q)
    );
    wire [1:0] _T_4002;
    BITS #(.width(64), .high(39), .low(38)) bits_5178 (
        .y(_T_4002),
        .in(_mem_reg_wdata__q)
    );
    wire [1:0] _T_4003;
    ASSINT #(.width(2)) assint_5179 (
        .y(_T_4003),
        .in(_T_4002)
    );
    wire _T_4005;
    wire [25:0] _WTEMP_707;
    PAD_UNSIGNED #(.width(1), .n(26)) u_pad_5180 (
        .y(_WTEMP_707),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(26)) u_eq_5181 (
        .y(_T_4005),
        .a(_T_4001),
        .b(_WTEMP_707)
    );
    wire _T_4007;
    wire [25:0] _WTEMP_708;
    PAD_UNSIGNED #(.width(1), .n(26)) u_pad_5182 (
        .y(_WTEMP_708),
        .in(1'h1)
    );
    EQ_UNSIGNED #(.width(26)) u_eq_5183 (
        .y(_T_4007),
        .a(_T_4001),
        .b(_WTEMP_708)
    );
    wire _T_4008;
    BITWISEOR #(.width(1)) bitwiseor_5184 (
        .y(_T_4008),
        .a(_T_4005),
        .b(_T_4007)
    );
    wire _T_4010;
    wire [1:0] _WTEMP_709;
    PAD_SIGNED #(.width(1), .n(2)) s_pad_5185 (
        .y(_WTEMP_709),
        .in(1'sh0)
    );
    NEQ_SIGNED #(.width(2)) s_neq_5186 (
        .y(_T_4010),
        .a(_T_4003),
        .b(_WTEMP_709)
    );
    wire [25:0] _T_4011;
    ASSINT #(.width(26)) assint_5187 (
        .y(_T_4011),
        .in(_T_4001)
    );
    wire _T_4013;
    wire [25:0] _WTEMP_710;
    PAD_SIGNED #(.width(1), .n(26)) s_pad_5188 (
        .y(_WTEMP_710),
        .in(-1'sh1)
    );
    EQ_SIGNED #(.width(26)) s_eq_5189 (
        .y(_T_4013),
        .a(_T_4011),
        .b(_WTEMP_710)
    );
    wire [25:0] _T_4014;
    ASSINT #(.width(26)) assint_5190 (
        .y(_T_4014),
        .in(_T_4001)
    );
    wire _T_4016;
    wire [25:0] _WTEMP_711;
    PAD_SIGNED #(.width(2), .n(26)) s_pad_5191 (
        .y(_WTEMP_711),
        .in(-2'sh2)
    );
    EQ_SIGNED #(.width(26)) s_eq_5192 (
        .y(_T_4016),
        .a(_T_4014),
        .b(_WTEMP_711)
    );
    wire _T_4017;
    BITWISEOR #(.width(1)) bitwiseor_5193 (
        .y(_T_4017),
        .a(_T_4013),
        .b(_T_4016)
    );
    wire _T_4019;
    wire [1:0] _WTEMP_712;
    PAD_SIGNED #(.width(1), .n(2)) s_pad_5194 (
        .y(_WTEMP_712),
        .in(-1'sh1)
    );
    EQ_SIGNED #(.width(2)) s_eq_5195 (
        .y(_T_4019),
        .a(_T_4003),
        .b(_WTEMP_712)
    );
    wire _T_4020;
    BITS #(.width(2), .high(0), .low(0)) bits_5196 (
        .y(_T_4020),
        .in(_T_4003)
    );
    wire _T_4021;
    MUX_UNSIGNED #(.width(1)) u_mux_5197 (
        .y(_T_4021),
        .sel(_T_4017),
        .a(_T_4019),
        .b(_T_4020)
    );
    wire _T_4022;
    MUX_UNSIGNED #(.width(1)) u_mux_5198 (
        .y(_T_4022),
        .sel(_T_4008),
        .a(_T_4010),
        .b(_T_4021)
    );
    wire [38:0] _T_4023;
    BITS #(.width(64), .high(38), .low(0)) bits_5199 (
        .y(_T_4023),
        .in(_mem_reg_wdata__q)
    );
    wire [39:0] _T_4024;
    CAT #(.width_a(1), .width_b(39)) cat_5200 (
        .y(_T_4024),
        .a(_T_4022),
        .b(_T_4023)
    );
    wire [39:0] _T_4025;
    ASSINT #(.width(40)) assint_5201 (
        .y(_T_4025),
        .in(_T_4024)
    );
    wire [39:0] _T_4026;
    MUX_SIGNED #(.width(40)) s_mux_5202 (
        .y(_T_4026),
        .sel(_mem_ctrl_jalr__q),
        .a(_T_4025),
        .b(mem_br_target)
    );
    wire [39:0] _T_4028;
    wire [39:0] _WTEMP_713;
    PAD_SIGNED #(.width(2), .n(40)) s_pad_5203 (
        .y(_WTEMP_713),
        .in(-2'sh2)
    );
    BITWISEAND #(.width(40)) bitwiseand_5204 (
        .y(_T_4028),
        .a(_T_4026),
        .b(_WTEMP_713)
    );
    wire [39:0] _T_4029;
    ASSINT #(.width(40)) assint_5205 (
        .y(_T_4029),
        .in(_T_4028)
    );
    wire [39:0] mem_npc;
    ASUINT #(.width(40)) asuint_5206 (
        .y(mem_npc),
        .in(_T_4029)
    );
    wire _T_4030;
    NEQ_UNSIGNED #(.width(40)) u_neq_5207 (
        .y(_T_4030),
        .a(mem_npc),
        .b(_ex_reg_pc__q)
    );
    wire _T_4031;
    NEQ_UNSIGNED #(.width(40)) u_neq_5208 (
        .y(_T_4031),
        .a(mem_npc),
        .b(_ibuf__io_pc)
    );
    wire _T_4033;
    MUX_UNSIGNED #(.width(1)) u_mux_5209 (
        .y(_T_4033),
        .sel(_ibuf__io_inst_0_valid),
        .a(_T_4031),
        .b(1'h1)
    );
    wire mem_misprediction;
    MUX_UNSIGNED #(.width(1)) u_mux_5210 (
        .y(mem_misprediction),
        .sel(ex_pc_valid),
        .a(_T_4030),
        .b(_T_4033)
    );
    wire _T_4034;
    BITS #(.width(32), .high(2), .low(2)) bits_5211 (
        .y(_T_4034),
        .in(_csr__io_status_isa)
    );
    wire _T_4036;
    EQ_UNSIGNED #(.width(1)) u_eq_5212 (
        .y(_T_4036),
        .a(_T_4034),
        .b(1'h0)
    );
    wire _T_4037;
    BITS #(.width(40), .high(1), .low(1)) bits_5213 (
        .y(_T_4037),
        .in(mem_npc)
    );
    wire mem_npc_misaligned;
    BITWISEAND #(.width(1)) bitwiseand_5214 (
        .y(mem_npc_misaligned),
        .a(_T_4036),
        .b(_T_4037)
    );
    wire _T_4039;
    EQ_UNSIGNED #(.width(1)) u_eq_5215 (
        .y(_T_4039),
        .a(_mem_reg_xcpt__q),
        .b(1'h0)
    );
    wire _T_4040;
    BITWISEXOR #(.width(1)) bitwisexor_5216 (
        .y(_T_4040),
        .a(_mem_ctrl_jalr__q),
        .b(mem_npc_misaligned)
    );
    wire _T_4041;
    BITWISEAND #(.width(1)) bitwiseand_5217 (
        .y(_T_4041),
        .a(_T_4039),
        .b(_T_4040)
    );
    wire [63:0] _T_4042;
    ASSINT #(.width(64)) assint_5218 (
        .y(_T_4042),
        .in(_mem_reg_wdata__q)
    );
    wire [63:0] _T_4043;
    wire [63:0] _WTEMP_714;
    PAD_SIGNED #(.width(40), .n(64)) s_pad_5219 (
        .y(_WTEMP_714),
        .in(mem_br_target)
    );
    MUX_SIGNED #(.width(64)) s_mux_5220 (
        .y(_T_4043),
        .sel(_T_4041),
        .a(_WTEMP_714),
        .b(_T_4042)
    );
    wire [63:0] mem_int_wdata;
    ASUINT #(.width(64)) asuint_5221 (
        .y(mem_int_wdata),
        .in(_T_4043)
    );
    wire _T_4044;
    BITWISEOR #(.width(1)) bitwiseor_5222 (
        .y(_T_4044),
        .a(_mem_ctrl_branch__q),
        .b(_mem_ctrl_jalr__q)
    );
    wire mem_cfi;
    BITWISEOR #(.width(1)) bitwiseor_5223 (
        .y(mem_cfi),
        .a(_T_4044),
        .b(_mem_ctrl_jal__q)
    );
    wire _T_4045;
    BITWISEAND #(.width(1)) bitwiseand_5224 (
        .y(_T_4045),
        .a(_mem_ctrl_branch__q),
        .b(mem_br_taken)
    );
    wire _T_4046;
    BITWISEOR #(.width(1)) bitwiseor_5225 (
        .y(_T_4046),
        .a(_T_4045),
        .b(_mem_ctrl_jalr__q)
    );
    wire _T_4048;
    BITWISEAND #(.width(1)) bitwiseand_5226 (
        .y(_T_4048),
        .a(1'h1),
        .b(_mem_ctrl_jal__q)
    );
    wire mem_cfi_taken;
    BITWISEOR #(.width(1)) bitwiseor_5227 (
        .y(mem_cfi_taken),
        .a(_T_4046),
        .b(_T_4048)
    );
    wire _T_4049;
    BITWISEAND #(.width(1)) bitwiseand_5228 (
        .y(_T_4049),
        .a(_mem_reg_btb_hit__q),
        .b(_mem_ctrl_branch__q)
    );
    wire _T_4050;
    NEQ_UNSIGNED #(.width(1)) u_neq_5229 (
        .y(_T_4050),
        .a(mem_br_taken),
        .b(_mem_reg_btb_resp_taken__q)
    );
    wire mem_direction_misprediction;
    BITWISEAND #(.width(1)) bitwiseand_5230 (
        .y(mem_direction_misprediction),
        .a(_T_4049),
        .b(_T_4050)
    );
    wire _T_4051;
    BITWISEOR #(.width(1)) bitwiseor_5231 (
        .y(_T_4051),
        .a(mem_misprediction),
        .b(_mem_reg_flush_pipe__q)
    );
    wire _T_4052;
    BITWISEAND #(.width(1)) bitwiseand_5232 (
        .y(_T_4052),
        .a(_mem_reg_valid__q),
        .b(_T_4051)
    );
    wire _T_4054;
    EQ_UNSIGNED #(.width(1)) u_eq_5233 (
        .y(_T_4054),
        .a(ctrl_killx),
        .b(1'h0)
    );
    wire _T_4056;
    EQ_UNSIGNED #(.width(1)) u_eq_5234 (
        .y(_T_4056),
        .a(take_pc_mem_wb),
        .b(1'h0)
    );
    wire _T_4057;
    BITWISEAND #(.width(1)) bitwiseand_5235 (
        .y(_T_4057),
        .a(_T_4056),
        .b(replay_ex)
    );
    wire _T_4059;
    EQ_UNSIGNED #(.width(1)) u_eq_5236 (
        .y(_T_4059),
        .a(ctrl_killx),
        .b(1'h0)
    );
    wire _T_4060;
    BITWISEAND #(.width(1)) bitwiseand_5237 (
        .y(_T_4060),
        .a(_T_4059),
        .b(ex_xcpt)
    );
    wire _T_4062;
    EQ_UNSIGNED #(.width(1)) u_eq_5238 (
        .y(_T_4062),
        .a(take_pc_mem_wb),
        .b(1'h0)
    );
    wire _T_4063;
    BITWISEAND #(.width(1)) bitwiseand_5239 (
        .y(_T_4063),
        .a(_T_4062),
        .b(_ex_reg_xcpt_interrupt__q)
    );
    wire _T_4065;
    wire [4:0] _WTEMP_715;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_5240 (
        .y(_WTEMP_715),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(5)) u_eq_5241 (
        .y(_T_4065),
        .a(_ex_ctrl_mem_cmd__q),
        .b(_WTEMP_715)
    );
    wire _T_4067;
    wire [4:0] _WTEMP_716;
    PAD_UNSIGNED #(.width(3), .n(5)) u_pad_5242 (
        .y(_WTEMP_716),
        .in(3'h6)
    );
    EQ_UNSIGNED #(.width(5)) u_eq_5243 (
        .y(_T_4067),
        .a(_ex_ctrl_mem_cmd__q),
        .b(_WTEMP_716)
    );
    wire _T_4068;
    BITWISEOR #(.width(1)) bitwiseor_5244 (
        .y(_T_4068),
        .a(_T_4065),
        .b(_T_4067)
    );
    wire _T_4070;
    wire [4:0] _WTEMP_717;
    PAD_UNSIGNED #(.width(3), .n(5)) u_pad_5245 (
        .y(_WTEMP_717),
        .in(3'h7)
    );
    EQ_UNSIGNED #(.width(5)) u_eq_5246 (
        .y(_T_4070),
        .a(_ex_ctrl_mem_cmd__q),
        .b(_WTEMP_717)
    );
    wire _T_4071;
    BITWISEOR #(.width(1)) bitwiseor_5247 (
        .y(_T_4071),
        .a(_T_4068),
        .b(_T_4070)
    );
    wire _T_4072;
    BITS #(.width(5), .high(3), .low(3)) bits_5248 (
        .y(_T_4072),
        .in(_ex_ctrl_mem_cmd__q)
    );
    wire _T_4074;
    wire [4:0] _WTEMP_718;
    PAD_UNSIGNED #(.width(3), .n(5)) u_pad_5249 (
        .y(_WTEMP_718),
        .in(3'h4)
    );
    EQ_UNSIGNED #(.width(5)) u_eq_5250 (
        .y(_T_4074),
        .a(_ex_ctrl_mem_cmd__q),
        .b(_WTEMP_718)
    );
    wire _T_4075;
    BITWISEOR #(.width(1)) bitwiseor_5251 (
        .y(_T_4075),
        .a(_T_4072),
        .b(_T_4074)
    );
    wire _T_4076;
    BITWISEOR #(.width(1)) bitwiseor_5252 (
        .y(_T_4076),
        .a(_T_4071),
        .b(_T_4075)
    );
    wire _T_4077;
    BITWISEAND #(.width(1)) bitwiseand_5253 (
        .y(_T_4077),
        .a(_ex_ctrl_mem__q),
        .b(_T_4076)
    );
    wire _T_4079;
    wire [4:0] _WTEMP_719;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_5254 (
        .y(_WTEMP_719),
        .in(1'h1)
    );
    EQ_UNSIGNED #(.width(5)) u_eq_5255 (
        .y(_T_4079),
        .a(_ex_ctrl_mem_cmd__q),
        .b(_WTEMP_719)
    );
    wire _T_4081;
    wire [4:0] _WTEMP_720;
    PAD_UNSIGNED #(.width(3), .n(5)) u_pad_5256 (
        .y(_WTEMP_720),
        .in(3'h7)
    );
    EQ_UNSIGNED #(.width(5)) u_eq_5257 (
        .y(_T_4081),
        .a(_ex_ctrl_mem_cmd__q),
        .b(_WTEMP_720)
    );
    wire _T_4082;
    BITWISEOR #(.width(1)) bitwiseor_5258 (
        .y(_T_4082),
        .a(_T_4079),
        .b(_T_4081)
    );
    wire _T_4083;
    BITS #(.width(5), .high(3), .low(3)) bits_5259 (
        .y(_T_4083),
        .in(_ex_ctrl_mem_cmd__q)
    );
    wire _T_4085;
    wire [4:0] _WTEMP_721;
    PAD_UNSIGNED #(.width(3), .n(5)) u_pad_5260 (
        .y(_WTEMP_721),
        .in(3'h4)
    );
    EQ_UNSIGNED #(.width(5)) u_eq_5261 (
        .y(_T_4085),
        .a(_ex_ctrl_mem_cmd__q),
        .b(_WTEMP_721)
    );
    wire _T_4086;
    BITWISEOR #(.width(1)) bitwiseor_5262 (
        .y(_T_4086),
        .a(_T_4083),
        .b(_T_4085)
    );
    wire _T_4087;
    BITWISEOR #(.width(1)) bitwiseor_5263 (
        .y(_T_4087),
        .a(_T_4082),
        .b(_T_4086)
    );
    wire _T_4088;
    BITWISEAND #(.width(1)) bitwiseand_5264 (
        .y(_T_4088),
        .a(_ex_ctrl_mem__q),
        .b(_T_4087)
    );
    wire _T_4089;
    BITWISEOR #(.width(1)) bitwiseor_5265 (
        .y(_T_4089),
        .a(_ex_ctrl_mem__q),
        .b(1'h0)
    );
    wire _T_4090;
    BITWISEAND #(.width(1)) bitwiseand_5266 (
        .y(_T_4090),
        .a(_ex_ctrl_rxs2__q),
        .b(_T_4089)
    );
    wire [6:0] _node_377;
    MUX_UNSIGNED #(.width(7)) u_mux_5267 (
        .y(_node_377),
        .sel(_ex_reg_btb_hit__q),
        .a(_ex_reg_btb_resp_bht_history__q),
        .b(_mem_reg_btb_resp_bht_history__q)
    );
    wire [1:0] _node_378;
    MUX_UNSIGNED #(.width(2)) u_mux_5268 (
        .y(_node_378),
        .sel(_ex_reg_btb_hit__q),
        .a(_ex_reg_btb_resp_bht_value__q),
        .b(_mem_reg_btb_resp_bht_value__q)
    );
    wire _node_379;
    MUX_UNSIGNED #(.width(1)) u_mux_5269 (
        .y(_node_379),
        .sel(_ex_reg_btb_hit__q),
        .a(_ex_reg_btb_resp_bridx__q),
        .b(_mem_reg_btb_resp_bridx__q)
    );
    wire [5:0] _node_380;
    MUX_UNSIGNED #(.width(6)) u_mux_5270 (
        .y(_node_380),
        .sel(_ex_reg_btb_hit__q),
        .a(_ex_reg_btb_resp_entry__q),
        .b(_mem_reg_btb_resp_entry__q)
    );
    wire [1:0] _node_381;
    MUX_UNSIGNED #(.width(2)) u_mux_5271 (
        .y(_node_381),
        .sel(_ex_reg_btb_hit__q),
        .a(_ex_reg_btb_resp_mask__q),
        .b(_mem_reg_btb_resp_mask__q)
    );
    wire _node_382;
    MUX_UNSIGNED #(.width(1)) u_mux_5272 (
        .y(_node_382),
        .sel(_ex_reg_btb_hit__q),
        .a(_ex_reg_btb_resp_taken__q),
        .b(_mem_reg_btb_resp_taken__q)
    );
    wire [38:0] _node_383;
    MUX_UNSIGNED #(.width(39)) u_mux_5273 (
        .y(_node_383),
        .sel(_ex_reg_btb_hit__q),
        .a(_ex_reg_btb_resp_target__q),
        .b(_mem_reg_btb_resp_target__q)
    );
    wire [63:0] _node_384;
    MUX_UNSIGNED #(.width(64)) u_mux_5274 (
        .y(_node_384),
        .sel(_T_4090),
        .a(ex_rs_1),
        .b(_mem_reg_rs2__q)
    );
    wire _T_4091;
    BITWISEAND #(.width(1)) bitwiseand_5275 (
        .y(_T_4091),
        .a(_mem_reg_load__q),
        .b(_bpu__io_xcpt_ld)
    );
    wire _T_4092;
    BITWISEAND #(.width(1)) bitwiseand_5276 (
        .y(_T_4092),
        .a(_mem_reg_store__q),
        .b(_bpu__io_xcpt_st)
    );
    wire mem_breakpoint;
    BITWISEOR #(.width(1)) bitwiseor_5277 (
        .y(mem_breakpoint),
        .a(_T_4091),
        .b(_T_4092)
    );
    wire _T_4093;
    BITWISEAND #(.width(1)) bitwiseand_5278 (
        .y(_T_4093),
        .a(_mem_reg_load__q),
        .b(_bpu__io_debug_ld)
    );
    wire _T_4094;
    BITWISEAND #(.width(1)) bitwiseand_5279 (
        .y(_T_4094),
        .a(_mem_reg_store__q),
        .b(_bpu__io_debug_st)
    );
    wire mem_debug_breakpoint;
    BITWISEOR #(.width(1)) bitwiseor_5280 (
        .y(mem_debug_breakpoint),
        .a(_T_4093),
        .b(_T_4094)
    );
    wire _T_4126;
    BITWISEAND #(.width(1)) bitwiseand_5281 (
        .y(_T_4126),
        .a(_mem_ctrl_mem__q),
        .b(io_dmem_xcpt_ma_st)
    );
    wire _T_4128;
    BITWISEAND #(.width(1)) bitwiseand_5282 (
        .y(_T_4128),
        .a(_mem_ctrl_mem__q),
        .b(io_dmem_xcpt_ma_ld)
    );
    wire _T_4130;
    BITWISEAND #(.width(1)) bitwiseand_5283 (
        .y(_T_4130),
        .a(_mem_ctrl_mem__q),
        .b(io_dmem_xcpt_pf_st)
    );
    wire _T_4132;
    BITWISEAND #(.width(1)) bitwiseand_5284 (
        .y(_T_4132),
        .a(_mem_ctrl_mem__q),
        .b(io_dmem_xcpt_pf_ld)
    );
    wire _T_4134;
    BITWISEOR #(.width(1)) bitwiseor_5285 (
        .y(_T_4134),
        .a(mem_debug_breakpoint),
        .b(mem_breakpoint)
    );
    wire _T_4135;
    BITWISEOR #(.width(1)) bitwiseor_5286 (
        .y(_T_4135),
        .a(_T_4134),
        .b(mem_npc_misaligned)
    );
    wire _T_4136;
    BITWISEOR #(.width(1)) bitwiseor_5287 (
        .y(_T_4136),
        .a(_T_4135),
        .b(_T_4126)
    );
    wire _T_4137;
    BITWISEOR #(.width(1)) bitwiseor_5288 (
        .y(_T_4137),
        .a(_T_4136),
        .b(_T_4128)
    );
    wire _T_4138;
    BITWISEOR #(.width(1)) bitwiseor_5289 (
        .y(_T_4138),
        .a(_T_4137),
        .b(_T_4130)
    );
    wire mem_new_xcpt;
    BITWISEOR #(.width(1)) bitwiseor_5290 (
        .y(mem_new_xcpt),
        .a(_T_4138),
        .b(_T_4132)
    );
    wire [2:0] _T_4139;
    MUX_UNSIGNED #(.width(3)) u_mux_5291 (
        .y(_T_4139),
        .sel(_T_4130),
        .a(3'h7),
        .b(3'h5)
    );
    wire [2:0] _T_4140;
    MUX_UNSIGNED #(.width(3)) u_mux_5292 (
        .y(_T_4140),
        .sel(_T_4128),
        .a(3'h4),
        .b(_T_4139)
    );
    wire [2:0] _T_4141;
    MUX_UNSIGNED #(.width(3)) u_mux_5293 (
        .y(_T_4141),
        .sel(_T_4126),
        .a(3'h6),
        .b(_T_4140)
    );
    wire [2:0] _T_4142;
    wire [2:0] _WTEMP_722;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_5294 (
        .y(_WTEMP_722),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(3)) u_mux_5295 (
        .y(_T_4142),
        .sel(mem_npc_misaligned),
        .a(_WTEMP_722),
        .b(_T_4141)
    );
    wire [2:0] _T_4143;
    wire [2:0] _WTEMP_723;
    PAD_UNSIGNED #(.width(2), .n(3)) u_pad_5296 (
        .y(_WTEMP_723),
        .in(2'h3)
    );
    MUX_UNSIGNED #(.width(3)) u_mux_5297 (
        .y(_T_4143),
        .sel(mem_breakpoint),
        .a(_WTEMP_723),
        .b(_T_4142)
    );
    wire [3:0] mem_new_cause;
    wire [3:0] _WTEMP_724;
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_5298 (
        .y(_WTEMP_724),
        .in(_T_4143)
    );
    MUX_UNSIGNED #(.width(4)) u_mux_5299 (
        .y(mem_new_cause),
        .sel(mem_debug_breakpoint),
        .a(4'hD),
        .b(_WTEMP_724)
    );
    wire _T_4144;
    BITWISEOR #(.width(1)) bitwiseor_5300 (
        .y(_T_4144),
        .a(_mem_reg_xcpt_interrupt__q),
        .b(_mem_reg_xcpt__q)
    );
    wire _T_4145;
    BITWISEAND #(.width(1)) bitwiseand_5301 (
        .y(_T_4145),
        .a(_mem_reg_valid__q),
        .b(mem_new_xcpt)
    );
    wire mem_xcpt;
    BITWISEOR #(.width(1)) bitwiseor_5302 (
        .y(mem_xcpt),
        .a(_T_4144),
        .b(_T_4145)
    );
    wire [63:0] mem_cause;
    wire [63:0] _WTEMP_725;
    PAD_UNSIGNED #(.width(4), .n(64)) u_pad_5303 (
        .y(_WTEMP_725),
        .in(mem_new_cause)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_5304 (
        .y(mem_cause),
        .sel(_T_4144),
        .a(_mem_reg_cause__q),
        .b(_WTEMP_725)
    );
    wire _T_4146;
    BITWISEAND #(.width(1)) bitwiseand_5305 (
        .y(_T_4146),
        .a(_mem_reg_valid__q),
        .b(_mem_ctrl_wxd__q)
    );
    wire dcache_kill_mem;
    BITWISEAND #(.width(1)) bitwiseand_5306 (
        .y(dcache_kill_mem),
        .a(_T_4146),
        .b(io_dmem_replay_next)
    );
    wire _T_4147;
    BITWISEAND #(.width(1)) bitwiseand_5307 (
        .y(_T_4147),
        .a(_mem_reg_valid__q),
        .b(_mem_ctrl_fp__q)
    );
    wire fpu_kill_mem;
    BITWISEAND #(.width(1)) bitwiseand_5308 (
        .y(fpu_kill_mem),
        .a(_T_4147),
        .b(io_fpu_nack_mem)
    );
    wire _T_4148;
    BITWISEOR #(.width(1)) bitwiseor_5309 (
        .y(_T_4148),
        .a(dcache_kill_mem),
        .b(_mem_reg_replay__q)
    );
    wire replay_mem;
    BITWISEOR #(.width(1)) bitwiseor_5310 (
        .y(replay_mem),
        .a(_T_4148),
        .b(fpu_kill_mem)
    );
    wire _T_4149;
    BITWISEOR #(.width(1)) bitwiseor_5311 (
        .y(_T_4149),
        .a(dcache_kill_mem),
        .b(take_pc_wb)
    );
    wire _T_4150;
    BITWISEOR #(.width(1)) bitwiseor_5312 (
        .y(_T_4150),
        .a(_T_4149),
        .b(_mem_reg_xcpt__q)
    );
    wire _T_4152;
    EQ_UNSIGNED #(.width(1)) u_eq_5313 (
        .y(_T_4152),
        .a(_mem_reg_valid__q),
        .b(1'h0)
    );
    wire killm_common;
    BITWISEOR #(.width(1)) bitwiseor_5314 (
        .y(killm_common),
        .a(_T_4150),
        .b(_T_4152)
    );
    wire _T_4153;
    BITWISEAND #(.width(1)) bitwiseand_5315 (
        .y(_T_4153),
        .a(_div__io_req_ready),
        .b(_div__io_req_valid)
    );
    wire __T_4154__q;
    wire __T_4154__d;
    DFF_POSCLK #(.width(1)) _T_4154 (
        .q(__T_4154__q),
        .d(__T_4154__d),
        .clk(clock)
    );
    wire _T_4155;
    BITWISEAND #(.width(1)) bitwiseand_5316 (
        .y(_T_4155),
        .a(killm_common),
        .b(__T_4154__q)
    );
    wire _T_4156;
    BITWISEOR #(.width(1)) bitwiseor_5317 (
        .y(_T_4156),
        .a(killm_common),
        .b(mem_xcpt)
    );
    wire ctrl_killm;
    BITWISEOR #(.width(1)) bitwiseor_5318 (
        .y(ctrl_killm),
        .a(_T_4156),
        .b(fpu_kill_mem)
    );
    wire _T_4158;
    EQ_UNSIGNED #(.width(1)) u_eq_5319 (
        .y(_T_4158),
        .a(ctrl_killm),
        .b(1'h0)
    );
    wire _T_4160;
    EQ_UNSIGNED #(.width(1)) u_eq_5320 (
        .y(_T_4160),
        .a(take_pc_wb),
        .b(1'h0)
    );
    wire _T_4161;
    BITWISEAND #(.width(1)) bitwiseand_5321 (
        .y(_T_4161),
        .a(replay_mem),
        .b(_T_4160)
    );
    wire _T_4163;
    EQ_UNSIGNED #(.width(1)) u_eq_5322 (
        .y(_T_4163),
        .a(take_pc_wb),
        .b(1'h0)
    );
    wire _T_4164;
    BITWISEAND #(.width(1)) bitwiseand_5323 (
        .y(_T_4164),
        .a(mem_xcpt),
        .b(_T_4163)
    );
    wire _T_4166;
    EQ_UNSIGNED #(.width(1)) u_eq_5324 (
        .y(_T_4166),
        .a(_mem_reg_xcpt__q),
        .b(1'h0)
    );
    wire _T_4167;
    BITWISEAND #(.width(1)) bitwiseand_5325 (
        .y(_T_4167),
        .a(_T_4166),
        .b(_mem_ctrl_fp__q)
    );
    wire _T_4168;
    BITWISEAND #(.width(1)) bitwiseand_5326 (
        .y(_T_4168),
        .a(_T_4167),
        .b(_mem_ctrl_wxd__q)
    );
    wire [63:0] _T_4169;
    MUX_UNSIGNED #(.width(64)) u_mux_5327 (
        .y(_T_4169),
        .sel(_T_4168),
        .a(io_fpu_toint_data),
        .b(mem_int_wdata)
    );
    wire wb_wxd;
    BITWISEAND #(.width(1)) bitwiseand_5328 (
        .y(wb_wxd),
        .a(_wb_reg_valid__q),
        .b(_wb_ctrl_wxd__q)
    );
    wire _T_4170;
    BITWISEOR #(.width(1)) bitwiseor_5329 (
        .y(_T_4170),
        .a(_wb_ctrl_div__q),
        .b(wb_dcache_miss)
    );
    wire wb_set_sboard;
    BITWISEOR #(.width(1)) bitwiseor_5330 (
        .y(wb_set_sboard),
        .a(_T_4170),
        .b(1'h0)
    );
    wire replay_wb_common;
    BITWISEOR #(.width(1)) bitwiseor_5331 (
        .y(replay_wb_common),
        .a(io_dmem_s2_nack),
        .b(_wb_reg_replay__q)
    );
    wire _T_4171;
    assign _T_4171 = 1'h0;
    wire _T_4173;
    EQ_UNSIGNED #(.width(1)) u_eq_5332 (
        .y(_T_4173),
        .a(io_rocc_cmd_ready),
        .b(1'h0)
    );
    wire replay_wb_rocc;
    assign replay_wb_rocc = 1'h0;
    wire replay_wb;
    BITWISEOR #(.width(1)) bitwiseor_5333 (
        .y(replay_wb),
        .a(replay_wb_common),
        .b(replay_wb_rocc)
    );
    wire _T_4174;
    BITWISEOR #(.width(1)) bitwiseor_5334 (
        .y(_T_4174),
        .a(replay_wb),
        .b(_wb_reg_xcpt__q)
    );
    wire _T_4175;
    BITWISEOR #(.width(1)) bitwiseor_5335 (
        .y(_T_4175),
        .a(_T_4174),
        .b(_csr__io_eret)
    );
    wire _T_4176;
    BITS #(.width(7), .high(0), .low(0)) bits_5336 (
        .y(_T_4176),
        .in(io_dmem_resp_bits_tag)
    );
    wire _T_4177;
    BITS #(.width(1), .high(0), .low(0)) bits_5337 (
        .y(_T_4177),
        .in(_T_4176)
    );
    wire dmem_resp_xpu;
    EQ_UNSIGNED #(.width(1)) u_eq_5338 (
        .y(dmem_resp_xpu),
        .a(_T_4177),
        .b(1'h0)
    );
    wire _T_4179;
    BITS #(.width(7), .high(0), .low(0)) bits_5339 (
        .y(_T_4179),
        .in(io_dmem_resp_bits_tag)
    );
    wire dmem_resp_fpu;
    BITS #(.width(1), .high(0), .low(0)) bits_5340 (
        .y(dmem_resp_fpu),
        .in(_T_4179)
    );
    wire [4:0] dmem_resp_waddr;
    BITS #(.width(7), .high(5), .low(1)) bits_5341 (
        .y(dmem_resp_waddr),
        .in(io_dmem_resp_bits_tag)
    );
    wire dmem_resp_valid;
    BITWISEAND #(.width(1)) bitwiseand_5342 (
        .y(dmem_resp_valid),
        .a(io_dmem_resp_valid),
        .b(io_dmem_resp_bits_has_data)
    );
    wire dmem_resp_replay;
    BITWISEAND #(.width(1)) bitwiseand_5343 (
        .y(dmem_resp_replay),
        .a(dmem_resp_valid),
        .b(io_dmem_resp_bits_replay)
    );
    wire _T_4181;
    EQ_UNSIGNED #(.width(1)) u_eq_5344 (
        .y(_T_4181),
        .a(wb_wxd),
        .b(1'h0)
    );
    wire [63:0] ll_wdata;
    wire [4:0] ll_waddr;
    wire _T_4182;
    BITWISEAND #(.width(1)) bitwiseand_5345 (
        .y(_T_4182),
        .a(_div__io_resp_ready),
        .b(_div__io_resp_valid)
    );
    wire ll_wen;
    wire _T_4183;
    BITWISEAND #(.width(1)) bitwiseand_5346 (
        .y(_T_4183),
        .a(dmem_resp_replay),
        .b(dmem_resp_xpu)
    );
    wire _T_4187;
    EQ_UNSIGNED #(.width(1)) u_eq_5347 (
        .y(_T_4187),
        .a(replay_wb),
        .b(1'h0)
    );
    wire _T_4188;
    BITWISEAND #(.width(1)) bitwiseand_5348 (
        .y(_T_4188),
        .a(_wb_reg_valid__q),
        .b(_T_4187)
    );
    wire _T_4190;
    EQ_UNSIGNED #(.width(1)) u_eq_5349 (
        .y(_T_4190),
        .a(_wb_reg_xcpt__q),
        .b(1'h0)
    );
    wire wb_valid;
    BITWISEAND #(.width(1)) bitwiseand_5350 (
        .y(wb_valid),
        .a(_T_4188),
        .b(_T_4190)
    );
    wire wb_wen;
    BITWISEAND #(.width(1)) bitwiseand_5351 (
        .y(wb_wen),
        .a(wb_valid),
        .b(_wb_ctrl_wxd__q)
    );
    wire rf_wen;
    BITWISEOR #(.width(1)) bitwiseor_5352 (
        .y(rf_wen),
        .a(wb_wen),
        .b(ll_wen)
    );
    wire [4:0] rf_waddr;
    MUX_UNSIGNED #(.width(5)) u_mux_5353 (
        .y(rf_waddr),
        .sel(ll_wen),
        .a(ll_waddr),
        .b(wb_waddr)
    );
    wire _T_4191;
    BITWISEAND #(.width(1)) bitwiseand_5354 (
        .y(_T_4191),
        .a(dmem_resp_valid),
        .b(dmem_resp_xpu)
    );
    wire _T_4193;
    NEQ_UNSIGNED #(.width(3)) u_neq_5355 (
        .y(_T_4193),
        .a(_wb_ctrl_csr__q),
        .b(3'h0)
    );
    wire [63:0] _T_4194;
    MUX_UNSIGNED #(.width(64)) u_mux_5356 (
        .y(_T_4194),
        .sel(_T_4193),
        .a(_csr__io_rw_rdata),
        .b(_wb_reg_wdata__q)
    );
    wire [63:0] _T_4195;
    MUX_UNSIGNED #(.width(64)) u_mux_5357 (
        .y(_T_4195),
        .sel(ll_wen),
        .a(ll_wdata),
        .b(_T_4194)
    );
    wire [63:0] rf_wdata;
    MUX_UNSIGNED #(.width(64)) u_mux_5358 (
        .y(rf_wdata),
        .sel(_T_4191),
        .a(io_dmem_resp_bits_data),
        .b(_T_4195)
    );
    wire _T_4197;
    wire [4:0] _WTEMP_726;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_5359 (
        .y(_WTEMP_726),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(5)) u_neq_5360 (
        .y(_T_4197),
        .a(rf_waddr),
        .b(_WTEMP_726)
    );
    wire [4:0] _T_4198;
    BITS #(.width(5), .high(4), .low(0)) bits_5361 (
        .y(_T_4198),
        .in(rf_waddr)
    );
    wire [4:0] _T_4199;
    BITWISENOT #(.width(5)) bitwisenot_5362 (
        .y(_T_4199),
        .in(_T_4198)
    );
    wire _node_385;
    BITWISEAND #(.width(1)) bitwiseand_5363 (
        .y(_node_385),
        .a(_T_4197),
        .b(rf_wen)
    );
    wire _node_386;
    BITWISEAND #(.width(1)) bitwiseand_5364 (
        .y(_node_386),
        .a(_T_4197),
        .b(rf_wen)
    );
    assign _T_3331__T_4200_addr = _T_4199;
    assign _T_3331__T_4200_en = _node_386;
    assign _T_3331__T_4200_clk = clock;
    assign _T_3331__T_4200_mask = 1'h1;
    wire _T_4201;
    EQ_UNSIGNED #(.width(5)) u_eq_5365 (
        .y(_T_4201),
        .a(rf_waddr),
        .b(_ibuf__io_inst_0_bits_inst_rs1)
    );
    wire _T_4202;
    EQ_UNSIGNED #(.width(5)) u_eq_5366 (
        .y(_T_4202),
        .a(rf_waddr),
        .b(_ibuf__io_inst_0_bits_inst_rs2)
    );
    wire [63:0] _node_387;
    MUX_UNSIGNED #(.width(64)) u_mux_5367 (
        .y(_node_387),
        .sel(_T_4201),
        .a(rf_wdata),
        .b(_T_3341)
    );
    wire [63:0] _node_388;
    MUX_UNSIGNED #(.width(64)) u_mux_5368 (
        .y(_node_388),
        .sel(_T_4202),
        .a(rf_wdata),
        .b(_T_3351)
    );
    wire [63:0] _node_389;
    assign _node_389 = rf_wdata;
    wire [63:0] _node_390;
    MUX_UNSIGNED #(.width(64)) u_mux_5369 (
        .y(_node_390),
        .sel(_T_4197),
        .a(_node_387),
        .b(_T_3341)
    );
    wire [63:0] _node_391;
    MUX_UNSIGNED #(.width(64)) u_mux_5370 (
        .y(_node_391),
        .sel(_T_4197),
        .a(_node_388),
        .b(_T_3351)
    );
    wire [11:0] _T_4203;
    BITS #(.width(32), .high(31), .low(20)) bits_5371 (
        .y(_T_4203),
        .in(_ibuf__io_inst_0_bits_raw)
    );
    wire [25:0] _T_4204;
    SHR_UNSIGNED #(.width(64), .n(38)) u_shr_5372 (
        .y(_T_4204),
        .in(_wb_reg_wdata__q)
    );
    wire [1:0] _T_4205;
    BITS #(.width(64), .high(39), .low(38)) bits_5373 (
        .y(_T_4205),
        .in(_wb_reg_wdata__q)
    );
    wire [1:0] _T_4206;
    ASSINT #(.width(2)) assint_5374 (
        .y(_T_4206),
        .in(_T_4205)
    );
    wire _T_4208;
    wire [25:0] _WTEMP_727;
    PAD_UNSIGNED #(.width(1), .n(26)) u_pad_5375 (
        .y(_WTEMP_727),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(26)) u_eq_5376 (
        .y(_T_4208),
        .a(_T_4204),
        .b(_WTEMP_727)
    );
    wire _T_4210;
    wire [25:0] _WTEMP_728;
    PAD_UNSIGNED #(.width(1), .n(26)) u_pad_5377 (
        .y(_WTEMP_728),
        .in(1'h1)
    );
    EQ_UNSIGNED #(.width(26)) u_eq_5378 (
        .y(_T_4210),
        .a(_T_4204),
        .b(_WTEMP_728)
    );
    wire _T_4211;
    BITWISEOR #(.width(1)) bitwiseor_5379 (
        .y(_T_4211),
        .a(_T_4208),
        .b(_T_4210)
    );
    wire _T_4213;
    wire [1:0] _WTEMP_729;
    PAD_SIGNED #(.width(1), .n(2)) s_pad_5380 (
        .y(_WTEMP_729),
        .in(1'sh0)
    );
    NEQ_SIGNED #(.width(2)) s_neq_5381 (
        .y(_T_4213),
        .a(_T_4206),
        .b(_WTEMP_729)
    );
    wire [25:0] _T_4214;
    ASSINT #(.width(26)) assint_5382 (
        .y(_T_4214),
        .in(_T_4204)
    );
    wire _T_4216;
    wire [25:0] _WTEMP_730;
    PAD_SIGNED #(.width(1), .n(26)) s_pad_5383 (
        .y(_WTEMP_730),
        .in(-1'sh1)
    );
    EQ_SIGNED #(.width(26)) s_eq_5384 (
        .y(_T_4216),
        .a(_T_4214),
        .b(_WTEMP_730)
    );
    wire [25:0] _T_4217;
    ASSINT #(.width(26)) assint_5385 (
        .y(_T_4217),
        .in(_T_4204)
    );
    wire _T_4219;
    wire [25:0] _WTEMP_731;
    PAD_SIGNED #(.width(2), .n(26)) s_pad_5386 (
        .y(_WTEMP_731),
        .in(-2'sh2)
    );
    EQ_SIGNED #(.width(26)) s_eq_5387 (
        .y(_T_4219),
        .a(_T_4217),
        .b(_WTEMP_731)
    );
    wire _T_4220;
    BITWISEOR #(.width(1)) bitwiseor_5388 (
        .y(_T_4220),
        .a(_T_4216),
        .b(_T_4219)
    );
    wire _T_4222;
    wire [1:0] _WTEMP_732;
    PAD_SIGNED #(.width(1), .n(2)) s_pad_5389 (
        .y(_WTEMP_732),
        .in(-1'sh1)
    );
    EQ_SIGNED #(.width(2)) s_eq_5390 (
        .y(_T_4222),
        .a(_T_4206),
        .b(_WTEMP_732)
    );
    wire _T_4223;
    BITS #(.width(2), .high(0), .low(0)) bits_5391 (
        .y(_T_4223),
        .in(_T_4206)
    );
    wire _T_4224;
    MUX_UNSIGNED #(.width(1)) u_mux_5392 (
        .y(_T_4224),
        .sel(_T_4220),
        .a(_T_4222),
        .b(_T_4223)
    );
    wire _T_4225;
    MUX_UNSIGNED #(.width(1)) u_mux_5393 (
        .y(_T_4225),
        .sel(_T_4211),
        .a(_T_4213),
        .b(_T_4224)
    );
    wire [38:0] _T_4226;
    BITS #(.width(64), .high(38), .low(0)) bits_5394 (
        .y(_T_4226),
        .in(_wb_reg_wdata__q)
    );
    wire [39:0] _T_4227;
    CAT #(.width_a(1), .width_b(39)) cat_5395 (
        .y(_T_4227),
        .a(_T_4225),
        .b(_T_4226)
    );
    wire [11:0] _T_4228;
    BITS #(.width(32), .high(31), .low(20)) bits_5396 (
        .y(_T_4228),
        .in(_wb_reg_inst__q)
    );
    wire [2:0] _T_4230;
    MUX_UNSIGNED #(.width(3)) u_mux_5397 (
        .y(_T_4230),
        .sel(_wb_reg_valid__q),
        .a(_wb_ctrl_csr__q),
        .b(3'h0)
    );
    wire _T_4232;
    wire [4:0] _WTEMP_733;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_5398 (
        .y(_WTEMP_733),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(5)) u_neq_5399 (
        .y(_T_4232),
        .a(_ibuf__io_inst_0_bits_inst_rs1),
        .b(_WTEMP_733)
    );
    wire _T_4233;
    BITWISEAND #(.width(1)) bitwiseand_5400 (
        .y(_T_4233),
        .a(id_ctrl_rxs1),
        .b(_T_4232)
    );
    wire _T_4235;
    wire [4:0] _WTEMP_734;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_5401 (
        .y(_WTEMP_734),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(5)) u_neq_5402 (
        .y(_T_4235),
        .a(_ibuf__io_inst_0_bits_inst_rs2),
        .b(_WTEMP_734)
    );
    wire _T_4236;
    BITWISEAND #(.width(1)) bitwiseand_5403 (
        .y(_T_4236),
        .a(id_ctrl_rxs2),
        .b(_T_4235)
    );
    wire _T_4238;
    wire [4:0] _WTEMP_735;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_5404 (
        .y(_WTEMP_735),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(5)) u_neq_5405 (
        .y(_T_4238),
        .a(_ibuf__io_inst_0_bits_inst_rd),
        .b(_WTEMP_735)
    );
    wire _T_4239;
    BITWISEAND #(.width(1)) bitwiseand_5406 (
        .y(_T_4239),
        .a(id_ctrl_wxd),
        .b(_T_4238)
    );
    wire [31:0] __T_4241__q;
    wire [31:0] __T_4241__d;
    DFF_POSCLK #(.width(32)) _T_4241 (
        .q(__T_4241__q),
        .d(__T_4241__d),
        .clk(clock)
    );
    wire [31:0] _WTEMP_736;
    MUX_UNSIGNED #(.width(32)) u_mux_5407 (
        .y(__T_4241__d),
        .sel(reset),
        .a(32'h0),
        .b(_WTEMP_736)
    );
    wire [30:0] _T_4242;
    SHR_UNSIGNED #(.width(32), .n(1)) u_shr_5408 (
        .y(_T_4242),
        .in(__T_4241__q)
    );
    wire [31:0] _T_4243;
    SHL_UNSIGNED #(.width(31), .n(1)) u_shl_5409 (
        .y(_T_4243),
        .in(_T_4242)
    );
    wire [31:0] _T_4246;
    DSHL_UNSIGNED #(.width_in(1), .width_n(5)) u_dshl_5410 (
        .y(_T_4246),
        .in(1'h1),
        .n(ll_waddr)
    );
    wire [31:0] _T_4248;
    wire [31:0] _WTEMP_737;
    PAD_UNSIGNED #(.width(1), .n(32)) u_pad_5411 (
        .y(_WTEMP_737),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(32)) u_mux_5412 (
        .y(_T_4248),
        .sel(ll_wen),
        .a(_T_4246),
        .b(_WTEMP_737)
    );
    wire [31:0] _T_4249;
    BITWISENOT #(.width(32)) bitwisenot_5413 (
        .y(_T_4249),
        .in(_T_4248)
    );
    wire [31:0] _T_4250;
    BITWISEAND #(.width(32)) bitwiseand_5414 (
        .y(_T_4250),
        .a(_T_4243),
        .b(_T_4249)
    );
    wire _T_4251;
    BITWISEOR #(.width(1)) bitwiseor_5415 (
        .y(_T_4251),
        .a(1'h0),
        .b(ll_wen)
    );
    wire [31:0] _T_4252;
    DSHR_UNSIGNED #(.width_in(32), .width_n(5)) u_dshr_5416 (
        .y(_T_4252),
        .in(_T_4243),
        .n(_ibuf__io_inst_0_bits_inst_rs1)
    );
    wire _T_4253;
    BITS #(.width(32), .high(0), .low(0)) bits_5417 (
        .y(_T_4253),
        .in(_T_4252)
    );
    wire _T_4254;
    BITWISEAND #(.width(1)) bitwiseand_5418 (
        .y(_T_4254),
        .a(_T_4233),
        .b(_T_4253)
    );
    wire [31:0] _T_4255;
    DSHR_UNSIGNED #(.width_in(32), .width_n(5)) u_dshr_5419 (
        .y(_T_4255),
        .in(_T_4243),
        .n(_ibuf__io_inst_0_bits_inst_rs2)
    );
    wire _T_4256;
    BITS #(.width(32), .high(0), .low(0)) bits_5420 (
        .y(_T_4256),
        .in(_T_4255)
    );
    wire _T_4257;
    BITWISEAND #(.width(1)) bitwiseand_5421 (
        .y(_T_4257),
        .a(_T_4236),
        .b(_T_4256)
    );
    wire [31:0] _T_4258;
    DSHR_UNSIGNED #(.width_in(32), .width_n(5)) u_dshr_5422 (
        .y(_T_4258),
        .in(_T_4243),
        .n(_ibuf__io_inst_0_bits_inst_rd)
    );
    wire _T_4259;
    BITS #(.width(32), .high(0), .low(0)) bits_5423 (
        .y(_T_4259),
        .in(_T_4258)
    );
    wire _T_4260;
    BITWISEAND #(.width(1)) bitwiseand_5424 (
        .y(_T_4260),
        .a(_T_4239),
        .b(_T_4259)
    );
    wire _T_4261;
    BITWISEOR #(.width(1)) bitwiseor_5425 (
        .y(_T_4261),
        .a(_T_4254),
        .b(_T_4257)
    );
    wire id_sboard_hazard;
    BITWISEOR #(.width(1)) bitwiseor_5426 (
        .y(id_sboard_hazard),
        .a(_T_4261),
        .b(_T_4260)
    );
    wire _T_4262;
    BITWISEAND #(.width(1)) bitwiseand_5427 (
        .y(_T_4262),
        .a(wb_set_sboard),
        .b(wb_wen)
    );
    wire [31:0] _T_4264;
    DSHL_UNSIGNED #(.width_in(1), .width_n(5)) u_dshl_5428 (
        .y(_T_4264),
        .in(1'h1),
        .n(wb_waddr)
    );
    wire [31:0] _T_4266;
    wire [31:0] _WTEMP_738;
    PAD_UNSIGNED #(.width(1), .n(32)) u_pad_5429 (
        .y(_WTEMP_738),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(32)) u_mux_5430 (
        .y(_T_4266),
        .sel(_T_4262),
        .a(_T_4264),
        .b(_WTEMP_738)
    );
    wire [31:0] _T_4267;
    BITWISEOR #(.width(32)) bitwiseor_5431 (
        .y(_T_4267),
        .a(_T_4250),
        .b(_T_4266)
    );
    wire _T_4268;
    BITWISEOR #(.width(1)) bitwiseor_5432 (
        .y(_T_4268),
        .a(_T_4251),
        .b(_T_4262)
    );
    wire [31:0] _node_392;
    MUX_UNSIGNED #(.width(32)) u_mux_5433 (
        .y(_node_392),
        .sel(_T_4251),
        .a(_T_4250),
        .b(__T_4241__q)
    );
    wire _T_4270;
    NEQ_UNSIGNED #(.width(3)) u_neq_5434 (
        .y(_T_4270),
        .a(_ex_ctrl_csr__q),
        .b(3'h0)
    );
    wire _T_4271;
    BITWISEOR #(.width(1)) bitwiseor_5435 (
        .y(_T_4271),
        .a(_T_4270),
        .b(_ex_ctrl_jalr__q)
    );
    wire _T_4272;
    BITWISEOR #(.width(1)) bitwiseor_5436 (
        .y(_T_4272),
        .a(_T_4271),
        .b(_ex_ctrl_mem__q)
    );
    wire _T_4273;
    BITWISEOR #(.width(1)) bitwiseor_5437 (
        .y(_T_4273),
        .a(_T_4272),
        .b(_ex_ctrl_div__q)
    );
    wire _T_4274;
    BITWISEOR #(.width(1)) bitwiseor_5438 (
        .y(_T_4274),
        .a(_T_4273),
        .b(_ex_ctrl_fp__q)
    );
    wire ex_cannot_bypass;
    BITWISEOR #(.width(1)) bitwiseor_5439 (
        .y(ex_cannot_bypass),
        .a(_T_4274),
        .b(1'h0)
    );
    wire _T_4275;
    EQ_UNSIGNED #(.width(5)) u_eq_5440 (
        .y(_T_4275),
        .a(_ibuf__io_inst_0_bits_inst_rs1),
        .b(ex_waddr)
    );
    wire _T_4276;
    BITWISEAND #(.width(1)) bitwiseand_5441 (
        .y(_T_4276),
        .a(_T_4233),
        .b(_T_4275)
    );
    wire _T_4277;
    EQ_UNSIGNED #(.width(5)) u_eq_5442 (
        .y(_T_4277),
        .a(_ibuf__io_inst_0_bits_inst_rs2),
        .b(ex_waddr)
    );
    wire _T_4278;
    BITWISEAND #(.width(1)) bitwiseand_5443 (
        .y(_T_4278),
        .a(_T_4236),
        .b(_T_4277)
    );
    wire _T_4279;
    EQ_UNSIGNED #(.width(5)) u_eq_5444 (
        .y(_T_4279),
        .a(_ibuf__io_inst_0_bits_inst_rd),
        .b(ex_waddr)
    );
    wire _T_4280;
    BITWISEAND #(.width(1)) bitwiseand_5445 (
        .y(_T_4280),
        .a(_T_4239),
        .b(_T_4279)
    );
    wire _T_4281;
    BITWISEOR #(.width(1)) bitwiseor_5446 (
        .y(_T_4281),
        .a(_T_4276),
        .b(_T_4278)
    );
    wire _T_4282;
    BITWISEOR #(.width(1)) bitwiseor_5447 (
        .y(_T_4282),
        .a(_T_4281),
        .b(_T_4280)
    );
    wire data_hazard_ex;
    BITWISEAND #(.width(1)) bitwiseand_5448 (
        .y(data_hazard_ex),
        .a(_ex_ctrl_wxd__q),
        .b(_T_4282)
    );
    wire _T_4283;
    EQ_UNSIGNED #(.width(5)) u_eq_5449 (
        .y(_T_4283),
        .a(_ibuf__io_inst_0_bits_inst_rs1),
        .b(ex_waddr)
    );
    wire _T_4284;
    BITWISEAND #(.width(1)) bitwiseand_5450 (
        .y(_T_4284),
        .a(io_fpu_dec_ren1),
        .b(_T_4283)
    );
    wire _T_4285;
    EQ_UNSIGNED #(.width(5)) u_eq_5451 (
        .y(_T_4285),
        .a(_ibuf__io_inst_0_bits_inst_rs2),
        .b(ex_waddr)
    );
    wire _T_4286;
    BITWISEAND #(.width(1)) bitwiseand_5452 (
        .y(_T_4286),
        .a(io_fpu_dec_ren2),
        .b(_T_4285)
    );
    wire _T_4287;
    EQ_UNSIGNED #(.width(5)) u_eq_5453 (
        .y(_T_4287),
        .a(_ibuf__io_inst_0_bits_inst_rs3),
        .b(ex_waddr)
    );
    wire _T_4288;
    BITWISEAND #(.width(1)) bitwiseand_5454 (
        .y(_T_4288),
        .a(io_fpu_dec_ren3),
        .b(_T_4287)
    );
    wire _T_4289;
    EQ_UNSIGNED #(.width(5)) u_eq_5455 (
        .y(_T_4289),
        .a(_ibuf__io_inst_0_bits_inst_rd),
        .b(ex_waddr)
    );
    wire _T_4290;
    BITWISEAND #(.width(1)) bitwiseand_5456 (
        .y(_T_4290),
        .a(io_fpu_dec_wen),
        .b(_T_4289)
    );
    wire _T_4291;
    BITWISEOR #(.width(1)) bitwiseor_5457 (
        .y(_T_4291),
        .a(_T_4284),
        .b(_T_4286)
    );
    wire _T_4292;
    BITWISEOR #(.width(1)) bitwiseor_5458 (
        .y(_T_4292),
        .a(_T_4291),
        .b(_T_4288)
    );
    wire _T_4293;
    BITWISEOR #(.width(1)) bitwiseor_5459 (
        .y(_T_4293),
        .a(_T_4292),
        .b(_T_4290)
    );
    wire fp_data_hazard_ex;
    BITWISEAND #(.width(1)) bitwiseand_5460 (
        .y(fp_data_hazard_ex),
        .a(_ex_ctrl_wfd__q),
        .b(_T_4293)
    );
    wire _T_4294;
    BITWISEAND #(.width(1)) bitwiseand_5461 (
        .y(_T_4294),
        .a(data_hazard_ex),
        .b(ex_cannot_bypass)
    );
    wire _T_4295;
    BITWISEOR #(.width(1)) bitwiseor_5462 (
        .y(_T_4295),
        .a(_T_4294),
        .b(fp_data_hazard_ex)
    );
    wire id_ex_hazard;
    BITWISEAND #(.width(1)) bitwiseand_5463 (
        .y(id_ex_hazard),
        .a(_ex_reg_valid__q),
        .b(_T_4295)
    );
    wire mem_mem_cmd_bh;
    BITWISEAND #(.width(1)) bitwiseand_5464 (
        .y(mem_mem_cmd_bh),
        .a(1'h1),
        .b(_mem_reg_slow_bypass__q)
    );
    wire _T_4298;
    NEQ_UNSIGNED #(.width(3)) u_neq_5465 (
        .y(_T_4298),
        .a(_mem_ctrl_csr__q),
        .b(3'h0)
    );
    wire _T_4299;
    BITWISEAND #(.width(1)) bitwiseand_5466 (
        .y(_T_4299),
        .a(_mem_ctrl_mem__q),
        .b(mem_mem_cmd_bh)
    );
    wire _T_4300;
    BITWISEOR #(.width(1)) bitwiseor_5467 (
        .y(_T_4300),
        .a(_T_4298),
        .b(_T_4299)
    );
    wire _T_4301;
    BITWISEOR #(.width(1)) bitwiseor_5468 (
        .y(_T_4301),
        .a(_T_4300),
        .b(_mem_ctrl_div__q)
    );
    wire _T_4302;
    BITWISEOR #(.width(1)) bitwiseor_5469 (
        .y(_T_4302),
        .a(_T_4301),
        .b(_mem_ctrl_fp__q)
    );
    wire mem_cannot_bypass;
    BITWISEOR #(.width(1)) bitwiseor_5470 (
        .y(mem_cannot_bypass),
        .a(_T_4302),
        .b(1'h0)
    );
    wire _T_4303;
    EQ_UNSIGNED #(.width(5)) u_eq_5471 (
        .y(_T_4303),
        .a(_ibuf__io_inst_0_bits_inst_rs1),
        .b(mem_waddr)
    );
    wire _T_4304;
    BITWISEAND #(.width(1)) bitwiseand_5472 (
        .y(_T_4304),
        .a(_T_4233),
        .b(_T_4303)
    );
    wire _T_4305;
    EQ_UNSIGNED #(.width(5)) u_eq_5473 (
        .y(_T_4305),
        .a(_ibuf__io_inst_0_bits_inst_rs2),
        .b(mem_waddr)
    );
    wire _T_4306;
    BITWISEAND #(.width(1)) bitwiseand_5474 (
        .y(_T_4306),
        .a(_T_4236),
        .b(_T_4305)
    );
    wire _T_4307;
    EQ_UNSIGNED #(.width(5)) u_eq_5475 (
        .y(_T_4307),
        .a(_ibuf__io_inst_0_bits_inst_rd),
        .b(mem_waddr)
    );
    wire _T_4308;
    BITWISEAND #(.width(1)) bitwiseand_5476 (
        .y(_T_4308),
        .a(_T_4239),
        .b(_T_4307)
    );
    wire _T_4309;
    BITWISEOR #(.width(1)) bitwiseor_5477 (
        .y(_T_4309),
        .a(_T_4304),
        .b(_T_4306)
    );
    wire _T_4310;
    BITWISEOR #(.width(1)) bitwiseor_5478 (
        .y(_T_4310),
        .a(_T_4309),
        .b(_T_4308)
    );
    wire data_hazard_mem;
    BITWISEAND #(.width(1)) bitwiseand_5479 (
        .y(data_hazard_mem),
        .a(_mem_ctrl_wxd__q),
        .b(_T_4310)
    );
    wire _T_4311;
    EQ_UNSIGNED #(.width(5)) u_eq_5480 (
        .y(_T_4311),
        .a(_ibuf__io_inst_0_bits_inst_rs1),
        .b(mem_waddr)
    );
    wire _T_4312;
    BITWISEAND #(.width(1)) bitwiseand_5481 (
        .y(_T_4312),
        .a(io_fpu_dec_ren1),
        .b(_T_4311)
    );
    wire _T_4313;
    EQ_UNSIGNED #(.width(5)) u_eq_5482 (
        .y(_T_4313),
        .a(_ibuf__io_inst_0_bits_inst_rs2),
        .b(mem_waddr)
    );
    wire _T_4314;
    BITWISEAND #(.width(1)) bitwiseand_5483 (
        .y(_T_4314),
        .a(io_fpu_dec_ren2),
        .b(_T_4313)
    );
    wire _T_4315;
    EQ_UNSIGNED #(.width(5)) u_eq_5484 (
        .y(_T_4315),
        .a(_ibuf__io_inst_0_bits_inst_rs3),
        .b(mem_waddr)
    );
    wire _T_4316;
    BITWISEAND #(.width(1)) bitwiseand_5485 (
        .y(_T_4316),
        .a(io_fpu_dec_ren3),
        .b(_T_4315)
    );
    wire _T_4317;
    EQ_UNSIGNED #(.width(5)) u_eq_5486 (
        .y(_T_4317),
        .a(_ibuf__io_inst_0_bits_inst_rd),
        .b(mem_waddr)
    );
    wire _T_4318;
    BITWISEAND #(.width(1)) bitwiseand_5487 (
        .y(_T_4318),
        .a(io_fpu_dec_wen),
        .b(_T_4317)
    );
    wire _T_4319;
    BITWISEOR #(.width(1)) bitwiseor_5488 (
        .y(_T_4319),
        .a(_T_4312),
        .b(_T_4314)
    );
    wire _T_4320;
    BITWISEOR #(.width(1)) bitwiseor_5489 (
        .y(_T_4320),
        .a(_T_4319),
        .b(_T_4316)
    );
    wire _T_4321;
    BITWISEOR #(.width(1)) bitwiseor_5490 (
        .y(_T_4321),
        .a(_T_4320),
        .b(_T_4318)
    );
    wire fp_data_hazard_mem;
    BITWISEAND #(.width(1)) bitwiseand_5491 (
        .y(fp_data_hazard_mem),
        .a(_mem_ctrl_wfd__q),
        .b(_T_4321)
    );
    wire _T_4322;
    BITWISEAND #(.width(1)) bitwiseand_5492 (
        .y(_T_4322),
        .a(data_hazard_mem),
        .b(mem_cannot_bypass)
    );
    wire _T_4323;
    BITWISEOR #(.width(1)) bitwiseor_5493 (
        .y(_T_4323),
        .a(_T_4322),
        .b(fp_data_hazard_mem)
    );
    wire id_mem_hazard;
    BITWISEAND #(.width(1)) bitwiseand_5494 (
        .y(id_mem_hazard),
        .a(_mem_reg_valid__q),
        .b(_T_4323)
    );
    wire _T_4324;
    BITWISEAND #(.width(1)) bitwiseand_5495 (
        .y(_T_4324),
        .a(_mem_reg_valid__q),
        .b(data_hazard_mem)
    );
    wire _T_4325;
    BITWISEAND #(.width(1)) bitwiseand_5496 (
        .y(_T_4325),
        .a(_T_4324),
        .b(_mem_ctrl_mem__q)
    );
    wire _T_4326;
    EQ_UNSIGNED #(.width(5)) u_eq_5497 (
        .y(_T_4326),
        .a(_ibuf__io_inst_0_bits_inst_rs1),
        .b(wb_waddr)
    );
    wire _T_4327;
    BITWISEAND #(.width(1)) bitwiseand_5498 (
        .y(_T_4327),
        .a(_T_4233),
        .b(_T_4326)
    );
    wire _T_4328;
    EQ_UNSIGNED #(.width(5)) u_eq_5499 (
        .y(_T_4328),
        .a(_ibuf__io_inst_0_bits_inst_rs2),
        .b(wb_waddr)
    );
    wire _T_4329;
    BITWISEAND #(.width(1)) bitwiseand_5500 (
        .y(_T_4329),
        .a(_T_4236),
        .b(_T_4328)
    );
    wire _T_4330;
    EQ_UNSIGNED #(.width(5)) u_eq_5501 (
        .y(_T_4330),
        .a(_ibuf__io_inst_0_bits_inst_rd),
        .b(wb_waddr)
    );
    wire _T_4331;
    BITWISEAND #(.width(1)) bitwiseand_5502 (
        .y(_T_4331),
        .a(_T_4239),
        .b(_T_4330)
    );
    wire _T_4332;
    BITWISEOR #(.width(1)) bitwiseor_5503 (
        .y(_T_4332),
        .a(_T_4327),
        .b(_T_4329)
    );
    wire _T_4333;
    BITWISEOR #(.width(1)) bitwiseor_5504 (
        .y(_T_4333),
        .a(_T_4332),
        .b(_T_4331)
    );
    wire data_hazard_wb;
    BITWISEAND #(.width(1)) bitwiseand_5505 (
        .y(data_hazard_wb),
        .a(_wb_ctrl_wxd__q),
        .b(_T_4333)
    );
    wire _T_4334;
    EQ_UNSIGNED #(.width(5)) u_eq_5506 (
        .y(_T_4334),
        .a(_ibuf__io_inst_0_bits_inst_rs1),
        .b(wb_waddr)
    );
    wire _T_4335;
    BITWISEAND #(.width(1)) bitwiseand_5507 (
        .y(_T_4335),
        .a(io_fpu_dec_ren1),
        .b(_T_4334)
    );
    wire _T_4336;
    EQ_UNSIGNED #(.width(5)) u_eq_5508 (
        .y(_T_4336),
        .a(_ibuf__io_inst_0_bits_inst_rs2),
        .b(wb_waddr)
    );
    wire _T_4337;
    BITWISEAND #(.width(1)) bitwiseand_5509 (
        .y(_T_4337),
        .a(io_fpu_dec_ren2),
        .b(_T_4336)
    );
    wire _T_4338;
    EQ_UNSIGNED #(.width(5)) u_eq_5510 (
        .y(_T_4338),
        .a(_ibuf__io_inst_0_bits_inst_rs3),
        .b(wb_waddr)
    );
    wire _T_4339;
    BITWISEAND #(.width(1)) bitwiseand_5511 (
        .y(_T_4339),
        .a(io_fpu_dec_ren3),
        .b(_T_4338)
    );
    wire _T_4340;
    EQ_UNSIGNED #(.width(5)) u_eq_5512 (
        .y(_T_4340),
        .a(_ibuf__io_inst_0_bits_inst_rd),
        .b(wb_waddr)
    );
    wire _T_4341;
    BITWISEAND #(.width(1)) bitwiseand_5513 (
        .y(_T_4341),
        .a(io_fpu_dec_wen),
        .b(_T_4340)
    );
    wire _T_4342;
    BITWISEOR #(.width(1)) bitwiseor_5514 (
        .y(_T_4342),
        .a(_T_4335),
        .b(_T_4337)
    );
    wire _T_4343;
    BITWISEOR #(.width(1)) bitwiseor_5515 (
        .y(_T_4343),
        .a(_T_4342),
        .b(_T_4339)
    );
    wire _T_4344;
    BITWISEOR #(.width(1)) bitwiseor_5516 (
        .y(_T_4344),
        .a(_T_4343),
        .b(_T_4341)
    );
    wire fp_data_hazard_wb;
    BITWISEAND #(.width(1)) bitwiseand_5517 (
        .y(fp_data_hazard_wb),
        .a(_wb_ctrl_wfd__q),
        .b(_T_4344)
    );
    wire _T_4345;
    BITWISEAND #(.width(1)) bitwiseand_5518 (
        .y(_T_4345),
        .a(data_hazard_wb),
        .b(wb_set_sboard)
    );
    wire _T_4346;
    BITWISEOR #(.width(1)) bitwiseor_5519 (
        .y(_T_4346),
        .a(_T_4345),
        .b(fp_data_hazard_wb)
    );
    wire id_wb_hazard;
    BITWISEAND #(.width(1)) bitwiseand_5520 (
        .y(id_wb_hazard),
        .a(_wb_reg_valid__q),
        .b(_T_4346)
    );
    wire [31:0] __T_4348__q;
    wire [31:0] __T_4348__d;
    DFF_POSCLK #(.width(32)) _T_4348 (
        .q(__T_4348__q),
        .d(__T_4348__d),
        .clk(clock)
    );
    wire [31:0] _WTEMP_739;
    MUX_UNSIGNED #(.width(32)) u_mux_5521 (
        .y(__T_4348__d),
        .sel(reset),
        .a(32'h0),
        .b(_WTEMP_739)
    );
    wire _T_4350;
    BITWISEAND #(.width(1)) bitwiseand_5522 (
        .y(_T_4350),
        .a(wb_dcache_miss),
        .b(_wb_ctrl_wfd__q)
    );
    wire _T_4351;
    BITWISEOR #(.width(1)) bitwiseor_5523 (
        .y(_T_4351),
        .a(_T_4350),
        .b(io_fpu_sboard_set)
    );
    wire _T_4352;
    BITWISEAND #(.width(1)) bitwiseand_5524 (
        .y(_T_4352),
        .a(_T_4351),
        .b(wb_valid)
    );
    wire [31:0] _T_4354;
    DSHL_UNSIGNED #(.width_in(1), .width_n(5)) u_dshl_5525 (
        .y(_T_4354),
        .in(1'h1),
        .n(wb_waddr)
    );
    wire [31:0] _T_4356;
    wire [31:0] _WTEMP_740;
    PAD_UNSIGNED #(.width(1), .n(32)) u_pad_5526 (
        .y(_WTEMP_740),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(32)) u_mux_5527 (
        .y(_T_4356),
        .sel(_T_4352),
        .a(_T_4354),
        .b(_WTEMP_740)
    );
    wire [31:0] _T_4357;
    BITWISEOR #(.width(32)) bitwiseor_5528 (
        .y(_T_4357),
        .a(__T_4348__q),
        .b(_T_4356)
    );
    wire _T_4358;
    BITWISEOR #(.width(1)) bitwiseor_5529 (
        .y(_T_4358),
        .a(1'h0),
        .b(_T_4352)
    );
    wire _T_4359;
    BITWISEAND #(.width(1)) bitwiseand_5530 (
        .y(_T_4359),
        .a(dmem_resp_replay),
        .b(dmem_resp_fpu)
    );
    wire [31:0] _T_4361;
    DSHL_UNSIGNED #(.width_in(1), .width_n(5)) u_dshl_5531 (
        .y(_T_4361),
        .in(1'h1),
        .n(dmem_resp_waddr)
    );
    wire [31:0] _T_4363;
    wire [31:0] _WTEMP_741;
    PAD_UNSIGNED #(.width(1), .n(32)) u_pad_5532 (
        .y(_WTEMP_741),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(32)) u_mux_5533 (
        .y(_T_4363),
        .sel(_T_4359),
        .a(_T_4361),
        .b(_WTEMP_741)
    );
    wire [31:0] _T_4364;
    BITWISENOT #(.width(32)) bitwisenot_5534 (
        .y(_T_4364),
        .in(_T_4363)
    );
    wire [31:0] _T_4365;
    BITWISEAND #(.width(32)) bitwiseand_5535 (
        .y(_T_4365),
        .a(_T_4357),
        .b(_T_4364)
    );
    wire _T_4366;
    BITWISEOR #(.width(1)) bitwiseor_5536 (
        .y(_T_4366),
        .a(_T_4358),
        .b(_T_4359)
    );
    wire [31:0] _node_393;
    MUX_UNSIGNED #(.width(32)) u_mux_5537 (
        .y(_node_393),
        .sel(_T_4358),
        .a(_T_4357),
        .b(__T_4348__q)
    );
    wire [31:0] _T_4368;
    DSHL_UNSIGNED #(.width_in(1), .width_n(5)) u_dshl_5538 (
        .y(_T_4368),
        .in(1'h1),
        .n(io_fpu_sboard_clra)
    );
    wire [31:0] _T_4370;
    wire [31:0] _WTEMP_742;
    PAD_UNSIGNED #(.width(1), .n(32)) u_pad_5539 (
        .y(_WTEMP_742),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(32)) u_mux_5540 (
        .y(_T_4370),
        .sel(io_fpu_sboard_clr),
        .a(_T_4368),
        .b(_WTEMP_742)
    );
    wire [31:0] _T_4371;
    BITWISENOT #(.width(32)) bitwisenot_5541 (
        .y(_T_4371),
        .in(_T_4370)
    );
    wire [31:0] _T_4372;
    BITWISEAND #(.width(32)) bitwiseand_5542 (
        .y(_T_4372),
        .a(_T_4365),
        .b(_T_4371)
    );
    wire _T_4373;
    BITWISEOR #(.width(1)) bitwiseor_5543 (
        .y(_T_4373),
        .a(_T_4366),
        .b(io_fpu_sboard_clr)
    );
    wire [31:0] _node_394;
    MUX_UNSIGNED #(.width(32)) u_mux_5544 (
        .y(_node_394),
        .sel(_T_4366),
        .a(_T_4365),
        .b(_node_393)
    );
    wire _T_4375;
    EQ_UNSIGNED #(.width(1)) u_eq_5545 (
        .y(_T_4375),
        .a(io_fpu_fcsr_rdy),
        .b(1'h0)
    );
    wire _T_4376;
    BITWISEAND #(.width(1)) bitwiseand_5546 (
        .y(_T_4376),
        .a(id_csr_en),
        .b(_T_4375)
    );
    wire [31:0] _T_4377;
    DSHR_UNSIGNED #(.width_in(32), .width_n(5)) u_dshr_5547 (
        .y(_T_4377),
        .in(__T_4348__q),
        .n(_ibuf__io_inst_0_bits_inst_rs1)
    );
    wire _T_4378;
    BITS #(.width(32), .high(0), .low(0)) bits_5548 (
        .y(_T_4378),
        .in(_T_4377)
    );
    wire _T_4379;
    BITWISEAND #(.width(1)) bitwiseand_5549 (
        .y(_T_4379),
        .a(io_fpu_dec_ren1),
        .b(_T_4378)
    );
    wire [31:0] _T_4380;
    DSHR_UNSIGNED #(.width_in(32), .width_n(5)) u_dshr_5550 (
        .y(_T_4380),
        .in(__T_4348__q),
        .n(_ibuf__io_inst_0_bits_inst_rs2)
    );
    wire _T_4381;
    BITS #(.width(32), .high(0), .low(0)) bits_5551 (
        .y(_T_4381),
        .in(_T_4380)
    );
    wire _T_4382;
    BITWISEAND #(.width(1)) bitwiseand_5552 (
        .y(_T_4382),
        .a(io_fpu_dec_ren2),
        .b(_T_4381)
    );
    wire [31:0] _T_4383;
    DSHR_UNSIGNED #(.width_in(32), .width_n(5)) u_dshr_5553 (
        .y(_T_4383),
        .in(__T_4348__q),
        .n(_ibuf__io_inst_0_bits_inst_rs3)
    );
    wire _T_4384;
    BITS #(.width(32), .high(0), .low(0)) bits_5554 (
        .y(_T_4384),
        .in(_T_4383)
    );
    wire _T_4385;
    BITWISEAND #(.width(1)) bitwiseand_5555 (
        .y(_T_4385),
        .a(io_fpu_dec_ren3),
        .b(_T_4384)
    );
    wire [31:0] _T_4386;
    DSHR_UNSIGNED #(.width_in(32), .width_n(5)) u_dshr_5556 (
        .y(_T_4386),
        .in(__T_4348__q),
        .n(_ibuf__io_inst_0_bits_inst_rd)
    );
    wire _T_4387;
    BITS #(.width(32), .high(0), .low(0)) bits_5557 (
        .y(_T_4387),
        .in(_T_4386)
    );
    wire _T_4388;
    BITWISEAND #(.width(1)) bitwiseand_5558 (
        .y(_T_4388),
        .a(io_fpu_dec_wen),
        .b(_T_4387)
    );
    wire _T_4389;
    BITWISEOR #(.width(1)) bitwiseor_5559 (
        .y(_T_4389),
        .a(_T_4379),
        .b(_T_4382)
    );
    wire _T_4390;
    BITWISEOR #(.width(1)) bitwiseor_5560 (
        .y(_T_4390),
        .a(_T_4389),
        .b(_T_4385)
    );
    wire _T_4391;
    BITWISEOR #(.width(1)) bitwiseor_5561 (
        .y(_T_4391),
        .a(_T_4390),
        .b(_T_4388)
    );
    wire id_stall_fpu;
    BITWISEOR #(.width(1)) bitwiseor_5562 (
        .y(id_stall_fpu),
        .a(_T_4376),
        .b(_T_4391)
    );
    wire _dcache_blocked__q;
    wire _dcache_blocked__d;
    DFF_POSCLK #(.width(1)) dcache_blocked (
        .q(_dcache_blocked__q),
        .d(_dcache_blocked__d),
        .clk(clock)
    );
    wire _T_4394;
    EQ_UNSIGNED #(.width(1)) u_eq_5563 (
        .y(_T_4394),
        .a(io_dmem_req_ready),
        .b(1'h0)
    );
    wire _T_4395;
    BITWISEOR #(.width(1)) bitwiseor_5564 (
        .y(_T_4395),
        .a(io_dmem_req_valid),
        .b(_dcache_blocked__q)
    );
    wire _T_4396;
    BITWISEAND #(.width(1)) bitwiseand_5565 (
        .y(_T_4396),
        .a(_T_4394),
        .b(_T_4395)
    );
    wire _rocc_blocked__q;
    wire _rocc_blocked__d;
    DFF_POSCLK #(.width(1)) rocc_blocked (
        .q(_rocc_blocked__q),
        .d(_rocc_blocked__d),
        .clk(clock)
    );
    wire _T_4399;
    EQ_UNSIGNED #(.width(1)) u_eq_5566 (
        .y(_T_4399),
        .a(_wb_reg_xcpt__q),
        .b(1'h0)
    );
    wire _T_4401;
    EQ_UNSIGNED #(.width(1)) u_eq_5567 (
        .y(_T_4401),
        .a(io_rocc_cmd_ready),
        .b(1'h0)
    );
    wire _T_4402;
    BITWISEAND #(.width(1)) bitwiseand_5568 (
        .y(_T_4402),
        .a(_T_4399),
        .b(_T_4401)
    );
    wire _T_4403;
    BITWISEOR #(.width(1)) bitwiseor_5569 (
        .y(_T_4403),
        .a(io_rocc_cmd_valid),
        .b(_rocc_blocked__q)
    );
    wire _T_4404;
    BITWISEAND #(.width(1)) bitwiseand_5570 (
        .y(_T_4404),
        .a(_T_4402),
        .b(_T_4403)
    );
    wire _T_4405;
    BITWISEOR #(.width(1)) bitwiseor_5571 (
        .y(_T_4405),
        .a(id_ex_hazard),
        .b(id_mem_hazard)
    );
    wire _T_4406;
    BITWISEOR #(.width(1)) bitwiseor_5572 (
        .y(_T_4406),
        .a(_T_4405),
        .b(id_wb_hazard)
    );
    wire _T_4407;
    BITWISEOR #(.width(1)) bitwiseor_5573 (
        .y(_T_4407),
        .a(_T_4406),
        .b(id_sboard_hazard)
    );
    wire _T_4408;
    BITWISEAND #(.width(1)) bitwiseand_5574 (
        .y(_T_4408),
        .a(id_ctrl_fp),
        .b(id_stall_fpu)
    );
    wire _T_4409;
    BITWISEOR #(.width(1)) bitwiseor_5575 (
        .y(_T_4409),
        .a(_T_4407),
        .b(_T_4408)
    );
    wire _T_4410;
    BITWISEAND #(.width(1)) bitwiseand_5576 (
        .y(_T_4410),
        .a(id_ctrl_mem),
        .b(_dcache_blocked__q)
    );
    wire _T_4411;
    BITWISEOR #(.width(1)) bitwiseor_5577 (
        .y(_T_4411),
        .a(_T_4409),
        .b(_T_4410)
    );
    wire _T_4412;
    BITWISEAND #(.width(1)) bitwiseand_5578 (
        .y(_T_4412),
        .a(id_ctrl_rocc),
        .b(_rocc_blocked__q)
    );
    wire _T_4413;
    BITWISEOR #(.width(1)) bitwiseor_5579 (
        .y(_T_4413),
        .a(_T_4411),
        .b(_T_4412)
    );
    wire _T_4415;
    EQ_UNSIGNED #(.width(1)) u_eq_5580 (
        .y(_T_4415),
        .a(wb_wxd),
        .b(1'h0)
    );
    wire _T_4416;
    BITWISEAND #(.width(1)) bitwiseand_5581 (
        .y(_T_4416),
        .a(_div__io_resp_valid),
        .b(_T_4415)
    );
    wire _T_4417;
    BITWISEOR #(.width(1)) bitwiseor_5582 (
        .y(_T_4417),
        .a(_div__io_req_ready),
        .b(_T_4416)
    );
    wire _T_4419;
    EQ_UNSIGNED #(.width(1)) u_eq_5583 (
        .y(_T_4419),
        .a(_T_4417),
        .b(1'h0)
    );
    wire _T_4420;
    BITWISEOR #(.width(1)) bitwiseor_5584 (
        .y(_T_4420),
        .a(_T_4419),
        .b(_div__io_req_valid)
    );
    wire _T_4421;
    BITWISEAND #(.width(1)) bitwiseand_5585 (
        .y(_T_4421),
        .a(id_ctrl_div),
        .b(_T_4420)
    );
    wire _T_4422;
    BITWISEOR #(.width(1)) bitwiseor_5586 (
        .y(_T_4422),
        .a(_T_4413),
        .b(_T_4421)
    );
    wire _T_4423;
    BITWISEOR #(.width(1)) bitwiseor_5587 (
        .y(_T_4423),
        .a(_T_4422),
        .b(id_do_fence)
    );
    wire ctrl_stalld;
    BITWISEOR #(.width(1)) bitwiseor_5588 (
        .y(ctrl_stalld),
        .a(_T_4423),
        .b(_csr__io_csr_stall)
    );
    wire _T_4425;
    EQ_UNSIGNED #(.width(1)) u_eq_5589 (
        .y(_T_4425),
        .a(_ibuf__io_inst_0_valid),
        .b(1'h0)
    );
    wire _T_4426;
    BITWISEOR #(.width(1)) bitwiseor_5590 (
        .y(_T_4426),
        .a(_T_4425),
        .b(_ibuf__io_inst_0_bits_replay)
    );
    wire _T_4427;
    BITWISEOR #(.width(1)) bitwiseor_5591 (
        .y(_T_4427),
        .a(_T_4426),
        .b(take_pc_mem_wb)
    );
    wire _T_4428;
    BITWISEOR #(.width(1)) bitwiseor_5592 (
        .y(_T_4428),
        .a(_T_4427),
        .b(ctrl_stalld)
    );
    wire _T_4429;
    BITWISEOR #(.width(1)) bitwiseor_5593 (
        .y(_T_4429),
        .a(_T_4428),
        .b(_csr__io_interrupt)
    );
    wire _T_4431;
    EQ_UNSIGNED #(.width(1)) u_eq_5594 (
        .y(_T_4431),
        .a(take_pc_wb),
        .b(1'h0)
    );
    wire _T_4432;
    BITWISEOR #(.width(1)) bitwiseor_5595 (
        .y(_T_4432),
        .a(_wb_reg_xcpt__q),
        .b(_csr__io_eret)
    );
    wire _T_4434;
    assign _T_4434 = 1'h1;
    wire [39:0] _T_4435;
    assign _T_4435 = mem_npc;
    wire [39:0] _T_4436;
    MUX_UNSIGNED #(.width(40)) u_mux_5596 (
        .y(_T_4436),
        .sel(replay_wb),
        .a(_wb_reg_pc__q),
        .b(_T_4435)
    );
    wire [39:0] _T_4437;
    MUX_UNSIGNED #(.width(40)) u_mux_5597 (
        .y(_T_4437),
        .sel(_T_4432),
        .a(_csr__io_evec),
        .b(_T_4436)
    );
    wire _T_4438;
    BITWISEAND #(.width(1)) bitwiseand_5598 (
        .y(_T_4438),
        .a(_wb_reg_valid__q),
        .b(_wb_ctrl_fence_i__q)
    );
    wire _T_4440;
    EQ_UNSIGNED #(.width(1)) u_eq_5599 (
        .y(_T_4440),
        .a(io_dmem_s2_nack),
        .b(1'h0)
    );
    wire _T_4441;
    BITWISEAND #(.width(1)) bitwiseand_5600 (
        .y(_T_4441),
        .a(_T_4438),
        .b(_T_4440)
    );
    wire _T_4443;
    EQ_UNSIGNED #(.width(1)) u_eq_5601 (
        .y(_T_4443),
        .a(ctrl_stalld),
        .b(1'h0)
    );
    wire _T_4444;
    BITWISEOR #(.width(1)) bitwiseor_5602 (
        .y(_T_4444),
        .a(_T_4443),
        .b(_csr__io_interrupt)
    );
    wire _T_4445;
    BITWISEAND #(.width(1)) bitwiseand_5603 (
        .y(_T_4445),
        .a(_mem_reg_replay__q),
        .b(_mem_reg_btb_hit__q)
    );
    wire _T_4447;
    EQ_UNSIGNED #(.width(1)) u_eq_5604 (
        .y(_T_4447),
        .a(take_pc_wb),
        .b(1'h0)
    );
    wire _T_4448;
    BITWISEAND #(.width(1)) bitwiseand_5605 (
        .y(_T_4448),
        .a(_mem_reg_valid__q),
        .b(_T_4447)
    );
    wire _T_4450;
    EQ_UNSIGNED #(.width(1)) u_eq_5606 (
        .y(_T_4450),
        .a(mem_cfi),
        .b(1'h0)
    );
    wire _T_4451;
    BITWISEOR #(.width(1)) bitwiseor_5607 (
        .y(_T_4451),
        .a(mem_cfi_taken),
        .b(_T_4450)
    );
    wire _T_4452;
    BITWISEAND #(.width(1)) bitwiseand_5608 (
        .y(_T_4452),
        .a(_T_4451),
        .b(mem_misprediction)
    );
    wire _T_4454;
    assign _T_4454 = 1'h0;
    wire _T_4456;
    EQ_UNSIGNED #(.width(1)) u_eq_5609 (
        .y(_T_4456),
        .a(_mem_reg_btb_hit__q),
        .b(1'h0)
    );
    wire _T_4457;
    assign _T_4457 = 1'h0;
    wire _T_4458;
    BITWISEOR #(.width(1)) bitwiseor_5610 (
        .y(_T_4458),
        .a(_T_4452),
        .b(_T_4457)
    );
    wire _T_4459;
    BITWISEAND #(.width(1)) bitwiseand_5611 (
        .y(_T_4459),
        .a(_T_4448),
        .b(_T_4458)
    );
    wire _T_4460;
    BITWISEOR #(.width(1)) bitwiseor_5612 (
        .y(_T_4460),
        .a(_T_4445),
        .b(_T_4459)
    );
    wire _T_4462;
    EQ_UNSIGNED #(.width(1)) u_eq_5613 (
        .y(_T_4462),
        .a(_mem_reg_replay__q),
        .b(1'h0)
    );
    wire _T_4463;
    BITWISEAND #(.width(1)) bitwiseand_5614 (
        .y(_T_4463),
        .a(_T_4462),
        .b(mem_cfi)
    );
    wire _T_4464;
    BITWISEOR #(.width(1)) bitwiseor_5615 (
        .y(_T_4464),
        .a(_mem_ctrl_jal__q),
        .b(_mem_ctrl_jalr__q)
    );
    wire [4:0] _T_4465;
    BITS #(.width(32), .high(19), .low(15)) bits_5616 (
        .y(_T_4465),
        .in(_mem_reg_inst__q)
    );
    wire [4:0] _T_4468;
    BITWISEAND #(.width(5)) bitwiseand_5617 (
        .y(_T_4468),
        .a(_T_4465),
        .b(5'h1B)
    );
    wire _T_4469;
    wire [4:0] _WTEMP_743;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_5618 (
        .y(_WTEMP_743),
        .in(1'h1)
    );
    EQ_UNSIGNED #(.width(5)) u_eq_5619 (
        .y(_T_4469),
        .a(_WTEMP_743),
        .b(_T_4468)
    );
    wire _T_4470;
    BITWISEAND #(.width(1)) bitwiseand_5620 (
        .y(_T_4470),
        .a(_mem_ctrl_jalr__q),
        .b(_T_4469)
    );
    wire [1:0] _T_4473;
    wire [1:0] _WTEMP_744;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_5621 (
        .y(_WTEMP_744),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_5622 (
        .y(_T_4473),
        .sel(_mem_reg_rvc__q),
        .a(_WTEMP_744),
        .b(2'h2)
    );
    wire [40:0] _T_4474;
    wire [39:0] _WTEMP_745;
    PAD_UNSIGNED #(.width(2), .n(40)) u_pad_5623 (
        .y(_WTEMP_745),
        .in(_T_4473)
    );
    ADD_UNSIGNED #(.width(40)) u_add_5624 (
        .y(_T_4474),
        .a(_mem_reg_pc__q),
        .b(_WTEMP_745)
    );
    wire [39:0] _T_4475;
    TAIL #(.width(41), .n(1)) tail_5625 (
        .y(_T_4475),
        .in(_T_4474)
    );
    wire [38:0] _T_4476;
    BITWISENOT #(.width(39)) bitwisenot_5626 (
        .y(_T_4476),
        .in(io_imem_btb_update_bits_br_pc)
    );
    wire [38:0] _T_4478;
    wire [38:0] _WTEMP_746;
    PAD_UNSIGNED #(.width(2), .n(39)) u_pad_5627 (
        .y(_WTEMP_746),
        .in(2'h3)
    );
    BITWISEOR #(.width(39)) bitwiseor_5628 (
        .y(_T_4478),
        .a(_T_4476),
        .b(_WTEMP_746)
    );
    wire [38:0] _T_4479;
    BITWISENOT #(.width(39)) bitwisenot_5629 (
        .y(_T_4479),
        .in(_T_4478)
    );
    wire _T_4481;
    EQ_UNSIGNED #(.width(1)) u_eq_5630 (
        .y(_T_4481),
        .a(take_pc_wb),
        .b(1'h0)
    );
    wire _T_4482;
    BITWISEAND #(.width(1)) bitwiseand_5631 (
        .y(_T_4482),
        .a(_mem_reg_valid__q),
        .b(_T_4481)
    );
    wire _T_4483;
    BITWISEAND #(.width(1)) bitwiseand_5632 (
        .y(_T_4483),
        .a(_T_4482),
        .b(_mem_ctrl_branch__q)
    );
    wire _T_4485;
    EQ_UNSIGNED #(.width(1)) u_eq_5633 (
        .y(_T_4485),
        .a(take_pc_wb),
        .b(1'h0)
    );
    wire _T_4486;
    BITWISEAND #(.width(1)) bitwiseand_5634 (
        .y(_T_4486),
        .a(_mem_reg_valid__q),
        .b(_T_4485)
    );
    wire _T_4487;
    BITS #(.width(5), .high(0), .low(0)) bits_5635 (
        .y(_T_4487),
        .in(mem_waddr)
    );
    wire _T_4488;
    BITWISEAND #(.width(1)) bitwiseand_5636 (
        .y(_T_4488),
        .a(io_imem_btb_update_bits_isJump),
        .b(_T_4487)
    );
    wire _T_4490;
    EQ_UNSIGNED #(.width(1)) u_eq_5637 (
        .y(_T_4490),
        .a(ctrl_killd),
        .b(1'h0)
    );
    wire _T_4491;
    BITWISEAND #(.width(1)) bitwiseand_5638 (
        .y(_T_4491),
        .a(_T_4490),
        .b(id_ctrl_fp)
    );
    wire _T_4492;
    BITWISEAND #(.width(1)) bitwiseand_5639 (
        .y(_T_4492),
        .a(dmem_resp_valid),
        .b(dmem_resp_fpu)
    );
    wire _T_4493;
    BITWISEAND #(.width(1)) bitwiseand_5640 (
        .y(_T_4493),
        .a(_ex_reg_valid__q),
        .b(_ex_ctrl_mem__q)
    );
    wire [5:0] ex_dcache_tag;
    CAT #(.width_a(5), .width_b(1)) cat_5641 (
        .y(ex_dcache_tag),
        .a(ex_waddr),
        .b(_ex_ctrl_fp__q)
    );
    wire [25:0] _T_4495;
    SHR_UNSIGNED #(.width(64), .n(38)) u_shr_5642 (
        .y(_T_4495),
        .in(ex_rs_0)
    );
    wire [1:0] _T_4496;
    BITS #(.width(64), .high(39), .low(38)) bits_5643 (
        .y(_T_4496),
        .in(_alu__io_adder_out)
    );
    wire [1:0] _T_4497;
    ASSINT #(.width(2)) assint_5644 (
        .y(_T_4497),
        .in(_T_4496)
    );
    wire _T_4499;
    wire [25:0] _WTEMP_747;
    PAD_UNSIGNED #(.width(1), .n(26)) u_pad_5645 (
        .y(_WTEMP_747),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(26)) u_eq_5646 (
        .y(_T_4499),
        .a(_T_4495),
        .b(_WTEMP_747)
    );
    wire _T_4501;
    wire [25:0] _WTEMP_748;
    PAD_UNSIGNED #(.width(1), .n(26)) u_pad_5647 (
        .y(_WTEMP_748),
        .in(1'h1)
    );
    EQ_UNSIGNED #(.width(26)) u_eq_5648 (
        .y(_T_4501),
        .a(_T_4495),
        .b(_WTEMP_748)
    );
    wire _T_4502;
    BITWISEOR #(.width(1)) bitwiseor_5649 (
        .y(_T_4502),
        .a(_T_4499),
        .b(_T_4501)
    );
    wire _T_4504;
    wire [1:0] _WTEMP_749;
    PAD_SIGNED #(.width(1), .n(2)) s_pad_5650 (
        .y(_WTEMP_749),
        .in(1'sh0)
    );
    NEQ_SIGNED #(.width(2)) s_neq_5651 (
        .y(_T_4504),
        .a(_T_4497),
        .b(_WTEMP_749)
    );
    wire [25:0] _T_4505;
    ASSINT #(.width(26)) assint_5652 (
        .y(_T_4505),
        .in(_T_4495)
    );
    wire _T_4507;
    wire [25:0] _WTEMP_750;
    PAD_SIGNED #(.width(1), .n(26)) s_pad_5653 (
        .y(_WTEMP_750),
        .in(-1'sh1)
    );
    EQ_SIGNED #(.width(26)) s_eq_5654 (
        .y(_T_4507),
        .a(_T_4505),
        .b(_WTEMP_750)
    );
    wire [25:0] _T_4508;
    ASSINT #(.width(26)) assint_5655 (
        .y(_T_4508),
        .in(_T_4495)
    );
    wire _T_4510;
    wire [25:0] _WTEMP_751;
    PAD_SIGNED #(.width(2), .n(26)) s_pad_5656 (
        .y(_WTEMP_751),
        .in(-2'sh2)
    );
    EQ_SIGNED #(.width(26)) s_eq_5657 (
        .y(_T_4510),
        .a(_T_4508),
        .b(_WTEMP_751)
    );
    wire _T_4511;
    BITWISEOR #(.width(1)) bitwiseor_5658 (
        .y(_T_4511),
        .a(_T_4507),
        .b(_T_4510)
    );
    wire _T_4513;
    wire [1:0] _WTEMP_752;
    PAD_SIGNED #(.width(1), .n(2)) s_pad_5659 (
        .y(_WTEMP_752),
        .in(-1'sh1)
    );
    EQ_SIGNED #(.width(2)) s_eq_5660 (
        .y(_T_4513),
        .a(_T_4497),
        .b(_WTEMP_752)
    );
    wire _T_4514;
    BITS #(.width(2), .high(0), .low(0)) bits_5661 (
        .y(_T_4514),
        .in(_T_4497)
    );
    wire _T_4515;
    MUX_UNSIGNED #(.width(1)) u_mux_5662 (
        .y(_T_4515),
        .sel(_T_4511),
        .a(_T_4513),
        .b(_T_4514)
    );
    wire _T_4516;
    MUX_UNSIGNED #(.width(1)) u_mux_5663 (
        .y(_T_4516),
        .sel(_T_4502),
        .a(_T_4504),
        .b(_T_4515)
    );
    wire [38:0] _T_4517;
    BITS #(.width(64), .high(38), .low(0)) bits_5664 (
        .y(_T_4517),
        .in(_alu__io_adder_out)
    );
    wire [39:0] _T_4518;
    CAT #(.width_a(1), .width_b(39)) cat_5665 (
        .y(_T_4518),
        .a(_T_4516),
        .b(_T_4517)
    );
    wire [63:0] _T_4519;
    MUX_UNSIGNED #(.width(64)) u_mux_5666 (
        .y(_T_4519),
        .sel(_mem_ctrl_fp__q),
        .a(io_fpu_store_data),
        .b(_mem_reg_rs2__q)
    );
    wire _T_4520;
    BITWISEOR #(.width(1)) bitwiseor_5667 (
        .y(_T_4520),
        .a(killm_common),
        .b(mem_breakpoint)
    );
    wire _T_4521;
    BITWISEAND #(.width(1)) bitwiseand_5668 (
        .y(_T_4521),
        .a(_mem_ctrl_mem__q),
        .b(mem_xcpt)
    );
    wire _T_4523;
    EQ_UNSIGNED #(.width(1)) u_eq_5669 (
        .y(_T_4523),
        .a(io_dmem_s1_kill),
        .b(1'h0)
    );
    wire _T_4524;
    BITWISEAND #(.width(1)) bitwiseand_5670 (
        .y(_T_4524),
        .a(_T_4521),
        .b(_T_4523)
    );
    wire [1:0] _T_4525;
    CAT #(.width_a(1), .width_b(1)) cat_5671 (
        .y(_T_4525),
        .a(io_dmem_xcpt_pf_ld),
        .b(io_dmem_xcpt_pf_st)
    );
    wire [1:0] _T_4526;
    CAT #(.width_a(1), .width_b(1)) cat_5672 (
        .y(_T_4526),
        .a(io_dmem_xcpt_ma_ld),
        .b(io_dmem_xcpt_ma_st)
    );
    wire [3:0] _T_4527;
    CAT #(.width_a(2), .width_b(2)) cat_5673 (
        .y(_T_4527),
        .a(_T_4526),
        .b(_T_4525)
    );
    wire _T_4529;
    wire [3:0] _WTEMP_753;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_5674 (
        .y(_WTEMP_753),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_5675 (
        .y(_T_4529),
        .a(_T_4527),
        .b(_WTEMP_753)
    );
    wire _T_4530;
    BITWISEOR #(.width(1)) bitwiseor_5676 (
        .y(_T_4530),
        .a(_T_4529),
        .b(reset)
    );
    wire _T_4532;
    EQ_UNSIGNED #(.width(1)) u_eq_5677 (
        .y(_T_4532),
        .a(_T_4530),
        .b(1'h0)
    );
    wire _T_4533;
    assign _T_4533 = 1'h0;
    wire _T_4535;
    EQ_UNSIGNED #(.width(1)) u_eq_5678 (
        .y(_T_4535),
        .a(replay_wb_common),
        .b(1'h0)
    );
    wire _T_4536;
    assign _T_4536 = 1'h0;
    wire _T_4538;
    wire [1:0] _WTEMP_754;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_5679 (
        .y(_WTEMP_754),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(2)) u_neq_5680 (
        .y(_T_4538),
        .a(_csr__io_status_xs),
        .b(_WTEMP_754)
    );
    wire _T_4539;
    BITWISEAND #(.width(1)) bitwiseand_5681 (
        .y(_T_4539),
        .a(_wb_reg_xcpt__q),
        .b(_T_4538)
    );
    wire [6:0] _T_4558_funct;
    wire [4:0] _T_4558_rs2;
    wire [4:0] _T_4558_rs1;
    wire _T_4558_xd;
    wire _T_4558_xs1;
    wire _T_4558_xs2;
    wire [4:0] _T_4558_rd;
    wire [6:0] _T_4558_opcode;
    wire [31:0] _T_4568;
    wire [6:0] _T_4569;
    BITS #(.width(32), .high(6), .low(0)) bits_5682 (
        .y(_T_4569),
        .in(_T_4568)
    );
    wire [4:0] _T_4570;
    BITS #(.width(32), .high(11), .low(7)) bits_5683 (
        .y(_T_4570),
        .in(_T_4568)
    );
    wire _T_4571;
    BITS #(.width(32), .high(12), .low(12)) bits_5684 (
        .y(_T_4571),
        .in(_T_4568)
    );
    wire _T_4572;
    BITS #(.width(32), .high(13), .low(13)) bits_5685 (
        .y(_T_4572),
        .in(_T_4568)
    );
    wire _T_4573;
    BITS #(.width(32), .high(14), .low(14)) bits_5686 (
        .y(_T_4573),
        .in(_T_4568)
    );
    wire [4:0] _T_4574;
    BITS #(.width(32), .high(19), .low(15)) bits_5687 (
        .y(_T_4574),
        .in(_T_4568)
    );
    wire [4:0] _T_4575;
    BITS #(.width(32), .high(24), .low(20)) bits_5688 (
        .y(_T_4575),
        .in(_T_4568)
    );
    wire [6:0] _T_4576;
    BITS #(.width(32), .high(31), .low(25)) bits_5689 (
        .y(_T_4576),
        .in(_T_4568)
    );
    wire [31:0] _T_4577;
    BITS #(.width(64), .high(31), .low(0)) bits_5690 (
        .y(_T_4577),
        .in(_csr__io_time)
    );
    wire [4:0] _T_4579;
    wire [4:0] _WTEMP_755;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_5691 (
        .y(_WTEMP_755),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(5)) u_mux_5692 (
        .y(_T_4579),
        .sel(rf_wen),
        .a(rf_waddr),
        .b(_WTEMP_755)
    );
    wire [4:0] _T_4580;
    BITS #(.width(32), .high(19), .low(15)) bits_5693 (
        .y(_T_4580),
        .in(_wb_reg_inst__q)
    );
    wire [63:0] __T_4581__q;
    wire [63:0] __T_4581__d;
    DFF_POSCLK #(.width(64)) _T_4581 (
        .q(__T_4581__q),
        .d(__T_4581__d),
        .clk(clock)
    );
    wire [63:0] __T_4582__q;
    wire [63:0] __T_4582__d;
    DFF_POSCLK #(.width(64)) _T_4582 (
        .q(__T_4582__q),
        .d(__T_4582__d),
        .clk(clock)
    );
    wire [4:0] _T_4583;
    BITS #(.width(32), .high(24), .low(20)) bits_5694 (
        .y(_T_4583),
        .in(_wb_reg_inst__q)
    );
    wire [63:0] __T_4584__q;
    wire [63:0] __T_4584__d;
    DFF_POSCLK #(.width(64)) _T_4584 (
        .q(__T_4584__q),
        .d(__T_4584__d),
        .clk(clock)
    );
    wire [63:0] __T_4585__q;
    wire [63:0] __T_4585__d;
    DFF_POSCLK #(.width(64)) _T_4585 (
        .q(__T_4585__q),
        .d(__T_4585__d),
        .clk(clock)
    );
    wire _T_4587;
    EQ_UNSIGNED #(.width(1)) u_eq_5695 (
        .y(_T_4587),
        .a(reset),
        .b(1'h0)
    );
    assign _T_3331__T_4200_data = _node_389;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_5696 (
        .y(_T_3803_0),
        .in(1'h0)
    );
    assign _T_3803_1 = 3'h4;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_5697 (
        .y(_T_3803_2),
        .in(1'h1)
    );
    assign _T_3803_3 = 3'h5;
    assign __T_4154__d = _T_4153;
    MUX_UNSIGNED #(.width(32)) u_mux_5698 (
        .y(_WTEMP_736),
        .sel(_T_4268),
        .a(_T_4267),
        .b(_node_392)
    );
    MUX_UNSIGNED #(.width(32)) u_mux_5699 (
        .y(_WTEMP_739),
        .sel(_T_4373),
        .a(_T_4372),
        .b(_node_394)
    );
    assign _T_4558_funct = _T_4576;
    assign _T_4558_opcode = _T_4569;
    assign _T_4558_rd = _T_4570;
    assign _T_4558_rs1 = _T_4574;
    assign _T_4558_rs2 = _T_4575;
    assign _T_4558_xd = _T_4573;
    assign _T_4558_xs1 = _T_4572;
    assign _T_4558_xs2 = _T_4571;
    assign _T_4568 = _wb_reg_inst__q;
    assign __T_4581__d = ex_rs_0;
    assign __T_4582__d = __T_4581__q;
    assign __T_4584__d = ex_rs_1;
    assign __T_4585__d = __T_4584__q;
    assign _alu__clock = clock;
    assign _alu__io_dw = _ex_ctrl_alu_dw__q;
    assign _alu__io_fn = _ex_ctrl_alu_fn__q;
    assign _alu__io_in1 = _T_3713;
    assign _alu__io_in2 = _T_3712;
    assign _alu__reset = reset;
    assign _bpu__clock = clock;
    assign _bpu__io_bp_0_address = _csr__io_bp_0_address;
    assign _bpu__io_bp_0_control_action = _csr__io_bp_0_control_action;
    assign _bpu__io_bp_0_control_chain = _csr__io_bp_0_control_chain;
    assign _bpu__io_bp_0_control_dmode = _csr__io_bp_0_control_dmode;
    assign _bpu__io_bp_0_control_h = _csr__io_bp_0_control_h;
    assign _bpu__io_bp_0_control_m = _csr__io_bp_0_control_m;
    assign _bpu__io_bp_0_control_maskmax = _csr__io_bp_0_control_maskmax;
    assign _bpu__io_bp_0_control_r = _csr__io_bp_0_control_r;
    assign _bpu__io_bp_0_control_reserved = _csr__io_bp_0_control_reserved;
    assign _bpu__io_bp_0_control_s = _csr__io_bp_0_control_s;
    assign _bpu__io_bp_0_control_tmatch = _csr__io_bp_0_control_tmatch;
    assign _bpu__io_bp_0_control_ttype = _csr__io_bp_0_control_ttype;
    assign _bpu__io_bp_0_control_u = _csr__io_bp_0_control_u;
    assign _bpu__io_bp_0_control_w = _csr__io_bp_0_control_w;
    assign _bpu__io_bp_0_control_x = _csr__io_bp_0_control_x;
    assign _bpu__io_bp_0_control_zero = _csr__io_bp_0_control_zero;
    BITS #(.width(64), .high(38), .low(0)) bits_5700 (
        .y(_bpu__io_ea),
        .in(_mem_reg_wdata__q)
    );
    BITS #(.width(40), .high(38), .low(0)) bits_5701 (
        .y(_bpu__io_pc),
        .in(_ibuf__io_pc)
    );
    assign _bpu__io_status_debug = _csr__io_status_debug;
    assign _bpu__io_status_fs = _csr__io_status_fs;
    assign _bpu__io_status_hie = _csr__io_status_hie;
    assign _bpu__io_status_hpie = _csr__io_status_hpie;
    assign _bpu__io_status_hpp = _csr__io_status_hpp;
    assign _bpu__io_status_isa = _csr__io_status_isa;
    assign _bpu__io_status_mie = _csr__io_status_mie;
    assign _bpu__io_status_mpie = _csr__io_status_mpie;
    assign _bpu__io_status_mpp = _csr__io_status_mpp;
    assign _bpu__io_status_mprv = _csr__io_status_mprv;
    assign _bpu__io_status_mxr = _csr__io_status_mxr;
    assign _bpu__io_status_prv = _csr__io_status_prv;
    assign _bpu__io_status_pum = _csr__io_status_pum;
    assign _bpu__io_status_sd = _csr__io_status_sd;
    assign _bpu__io_status_sd_rv32 = _csr__io_status_sd_rv32;
    assign _bpu__io_status_sie = _csr__io_status_sie;
    assign _bpu__io_status_spie = _csr__io_status_spie;
    assign _bpu__io_status_spp = _csr__io_status_spp;
    assign _bpu__io_status_sxl = _csr__io_status_sxl;
    assign _bpu__io_status_tsr = _csr__io_status_tsr;
    assign _bpu__io_status_tvm = _csr__io_status_tvm;
    assign _bpu__io_status_tw = _csr__io_status_tw;
    assign _bpu__io_status_uie = _csr__io_status_uie;
    assign _bpu__io_status_upie = _csr__io_status_upie;
    assign _bpu__io_status_uxl = _csr__io_status_uxl;
    assign _bpu__io_status_xs = _csr__io_status_xs;
    assign _bpu__io_status_zero1 = _csr__io_status_zero1;
    assign _bpu__io_status_zero2 = _csr__io_status_zero2;
    assign _bpu__reset = reset;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_5702 (
        .y(bypass_mux_0),
        .in(1'h0)
    );
    assign bypass_mux_1 = _mem_reg_wdata__q;
    assign bypass_mux_2 = _wb_reg_wdata__q;
    assign bypass_mux_3 = io_dmem_resp_bits_data_word_bypass;
    assign _csr__clock = clock;
    assign _csr__io_badaddr = _T_4227;
    assign _csr__io_cause = _wb_reg_cause__q;
    assign _csr__io_decode_csr = _T_4203;
    assign _csr__io_exception = _wb_reg_xcpt__q;
    assign _csr__io_fcsr_flags_bits = io_fpu_fcsr_flags_bits;
    assign _csr__io_fcsr_flags_valid = io_fpu_fcsr_flags_valid;
    assign _csr__io_hartid = io_hartid;
    assign _csr__io_interrupts_debug = io_interrupts_debug;
    assign _csr__io_interrupts_meip = io_interrupts_meip;
    assign _csr__io_interrupts_msip = io_interrupts_msip;
    assign _csr__io_interrupts_mtip = io_interrupts_mtip;
    assign _csr__io_interrupts_seip = io_interrupts_seip;
    assign _csr__io_pc = _wb_reg_pc__q;
    assign _csr__io_retire = wb_valid;
    assign _csr__io_rocc_interrupt = io_rocc_interrupt;
    assign _csr__io_rw_addr = _T_4228;
    assign _csr__io_rw_cmd = _T_4230;
    assign _csr__io_rw_wdata = _wb_reg_wdata__q;
    assign _csr__reset = reset;
    assign ctrl_killd = _T_4429;
    assign _dcache_blocked__d = _T_4396;
    assign _div__clock = clock;
    assign _div__io_kill = _T_4155;
    assign _div__io_req_bits_dw = _ex_ctrl_alu_dw__q;
    assign _div__io_req_bits_fn = _ex_ctrl_alu_fn__q;
    assign _div__io_req_bits_in1 = ex_rs_0;
    assign _div__io_req_bits_in2 = ex_rs_1;
    assign _div__io_req_bits_tag = ex_waddr;
    assign _div__io_req_valid = _T_3714;
    MUX_UNSIGNED #(.width(1)) u_mux_5703 (
        .y(_div__io_resp_ready),
        .sel(_T_4183),
        .a(1'h0),
        .b(_T_4181)
    );
    assign _div__reset = reset;
    MUX_UNSIGNED #(.width(64)) u_mux_5704 (
        .y(_ex_cause__d),
        .sel(id_xcpt),
        .a(id_cause),
        .b(_ex_cause__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_5705 (
        .y(_ex_ctrl_alu_dw__d),
        .sel(_T_3729),
        .a(_node_366),
        .b(_ex_ctrl_alu_dw__q)
    );
    MUX_UNSIGNED #(.width(4)) u_mux_5706 (
        .y(_ex_ctrl_alu_fn__d),
        .sel(_T_3729),
        .a(_node_367),
        .b(_ex_ctrl_alu_fn__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_5707 (
        .y(_ex_ctrl_branch__d),
        .sel(_T_3729),
        .a(id_ctrl_branch),
        .b(_ex_ctrl_branch__q)
    );
    MUX_UNSIGNED #(.width(3)) u_mux_5708 (
        .y(_ex_ctrl_csr__d),
        .sel(_T_3729),
        .a(id_csr),
        .b(_ex_ctrl_csr__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_5709 (
        .y(_ex_ctrl_div__d),
        .sel(_T_3729),
        .a(id_ctrl_div),
        .b(_ex_ctrl_div__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_5710 (
        .y(_ex_ctrl_fence_i__d),
        .sel(_T_3729),
        .a(_node_368),
        .b(_ex_ctrl_fence_i__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_5711 (
        .y(_ex_ctrl_fp__d),
        .sel(_T_3729),
        .a(id_ctrl_fp),
        .b(_ex_ctrl_fp__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_5712 (
        .y(_ex_ctrl_jal__d),
        .sel(_T_3729),
        .a(id_ctrl_jal),
        .b(_ex_ctrl_jal__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_5713 (
        .y(_ex_ctrl_jalr__d),
        .sel(_T_3729),
        .a(id_ctrl_jalr),
        .b(_ex_ctrl_jalr__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_5714 (
        .y(_ex_ctrl_mem__d),
        .sel(_T_3729),
        .a(id_ctrl_mem),
        .b(_ex_ctrl_mem__q)
    );
    MUX_UNSIGNED #(.width(5)) u_mux_5715 (
        .y(_ex_ctrl_mem_cmd__d),
        .sel(_T_3729),
        .a(id_ctrl_mem_cmd),
        .b(_ex_ctrl_mem_cmd__q)
    );
    MUX_UNSIGNED #(.width(3)) u_mux_5716 (
        .y(_ex_ctrl_mem_type__d),
        .sel(_T_3729),
        .a(id_ctrl_mem_type),
        .b(_ex_ctrl_mem_type__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_5717 (
        .y(_ex_ctrl_rxs2__d),
        .sel(_T_3729),
        .a(id_ctrl_rxs2),
        .b(_ex_ctrl_rxs2__q)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_5718 (
        .y(_ex_ctrl_sel_alu1__d),
        .sel(_T_3729),
        .a(_node_369),
        .b(_ex_ctrl_sel_alu1__q)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_5719 (
        .y(_ex_ctrl_sel_alu2__d),
        .sel(_T_3729),
        .a(_node_370),
        .b(_ex_ctrl_sel_alu2__q)
    );
    MUX_UNSIGNED #(.width(3)) u_mux_5720 (
        .y(_ex_ctrl_sel_imm__d),
        .sel(_T_3729),
        .a(id_ctrl_sel_imm),
        .b(_ex_ctrl_sel_imm__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_5721 (
        .y(_ex_ctrl_wfd__d),
        .sel(_T_3729),
        .a(id_ctrl_wfd),
        .b(_ex_ctrl_wfd__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_5722 (
        .y(_ex_ctrl_wxd__d),
        .sel(_T_3729),
        .a(id_ctrl_wxd),
        .b(_ex_ctrl_wxd__q)
    );
    assign _ex_reg_btb_hit__d = _ibuf__io_inst_0_bits_btb_hit;
    MUX_UNSIGNED #(.width(7)) u_mux_5723 (
        .y(_ex_reg_btb_resp_bht_history__d),
        .sel(_ibuf__io_inst_0_bits_btb_hit),
        .a(_ibuf__io_btb_resp_bht_history),
        .b(_ex_reg_btb_resp_bht_history__q)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_5724 (
        .y(_ex_reg_btb_resp_bht_value__d),
        .sel(_ibuf__io_inst_0_bits_btb_hit),
        .a(_ibuf__io_btb_resp_bht_value),
        .b(_ex_reg_btb_resp_bht_value__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_5725 (
        .y(_ex_reg_btb_resp_bridx__d),
        .sel(_ibuf__io_inst_0_bits_btb_hit),
        .a(_ibuf__io_btb_resp_bridx),
        .b(_ex_reg_btb_resp_bridx__q)
    );
    MUX_UNSIGNED #(.width(6)) u_mux_5726 (
        .y(_ex_reg_btb_resp_entry__d),
        .sel(_ibuf__io_inst_0_bits_btb_hit),
        .a(_ibuf__io_btb_resp_entry),
        .b(_ex_reg_btb_resp_entry__q)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_5727 (
        .y(_ex_reg_btb_resp_mask__d),
        .sel(_ibuf__io_inst_0_bits_btb_hit),
        .a(_ibuf__io_btb_resp_mask),
        .b(_ex_reg_btb_resp_mask__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_5728 (
        .y(_ex_reg_btb_resp_taken__d),
        .sel(_ibuf__io_inst_0_bits_btb_hit),
        .a(_ibuf__io_btb_resp_taken),
        .b(_ex_reg_btb_resp_taken__q)
    );
    MUX_UNSIGNED #(.width(39)) u_mux_5729 (
        .y(_ex_reg_btb_resp_target__d),
        .sel(_ibuf__io_inst_0_bits_btb_hit),
        .a(_ibuf__io_btb_resp_target),
        .b(_ex_reg_btb_resp_target__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_5730 (
        .y(_ex_reg_flush_pipe__d),
        .sel(_T_3729),
        .a(_node_371),
        .b(_ex_reg_flush_pipe__q)
    );
    MUX_UNSIGNED #(.width(32)) u_mux_5731 (
        .y(_ex_reg_inst__d),
        .sel(_T_3780),
        .a(_ibuf__io_inst_0_bits_inst_bits),
        .b(_ex_reg_inst__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_5732 (
        .y(_ex_reg_load_use__d),
        .sel(_T_3729),
        .a(id_load_use),
        .b(_ex_reg_load_use__q)
    );
    MUX_UNSIGNED #(.width(40)) u_mux_5733 (
        .y(_ex_reg_pc__d),
        .sel(_T_3780),
        .a(_ibuf__io_pc),
        .b(_ex_reg_pc__q)
    );
    assign _ex_reg_replay__d = _T_3720;
    MUX_UNSIGNED #(.width(1)) u_mux_5734 (
        .y(_ex_reg_rs_bypass_0__d),
        .sel(_T_3729),
        .a(_T_3749),
        .b(_ex_reg_rs_bypass_0__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_5735 (
        .y(_ex_reg_rs_bypass_1__d),
        .sel(_T_3729),
        .a(_T_3764),
        .b(_ex_reg_rs_bypass_1__q)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_5736 (
        .y(_ex_reg_rs_lsb_0__d),
        .sel(_T_3729),
        .a(_node_372),
        .b(_ex_reg_rs_lsb_0__q)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_5737 (
        .y(_ex_reg_rs_lsb_1__d),
        .sel(_T_3729),
        .a(_node_373),
        .b(_ex_reg_rs_lsb_1__q)
    );
    MUX_UNSIGNED #(.width(62)) u_mux_5738 (
        .y(_ex_reg_rs_msb_0__d),
        .sel(_T_3729),
        .a(_node_374),
        .b(_ex_reg_rs_msb_0__q)
    );
    MUX_UNSIGNED #(.width(62)) u_mux_5739 (
        .y(_ex_reg_rs_msb_1__d),
        .sel(_T_3729),
        .a(_node_375),
        .b(_ex_reg_rs_msb_1__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_5740 (
        .y(_ex_reg_rvc__d),
        .sel(_T_3729),
        .a(_node_376),
        .b(_ex_reg_rvc__q)
    );
    assign _ex_reg_valid__d = _T_3716;
    assign _ex_reg_xcpt__d = _T_3723;
    assign _ex_reg_xcpt_interrupt__d = _T_3727;
    assign _ibuf__clock = clock;
    assign _ibuf__io_imem_bits_btb_bits_bht_history = io_imem_resp_bits_btb_bits_bht_history;
    assign _ibuf__io_imem_bits_btb_bits_bht_value = io_imem_resp_bits_btb_bits_bht_value;
    assign _ibuf__io_imem_bits_btb_bits_bridx = io_imem_resp_bits_btb_bits_bridx;
    assign _ibuf__io_imem_bits_btb_bits_entry = io_imem_resp_bits_btb_bits_entry;
    assign _ibuf__io_imem_bits_btb_bits_mask = io_imem_resp_bits_btb_bits_mask;
    assign _ibuf__io_imem_bits_btb_bits_taken = io_imem_resp_bits_btb_bits_taken;
    assign _ibuf__io_imem_bits_btb_bits_target = io_imem_resp_bits_btb_bits_target;
    assign _ibuf__io_imem_bits_btb_valid = io_imem_resp_bits_btb_valid;
    assign _ibuf__io_imem_bits_data = io_imem_resp_bits_data;
    assign _ibuf__io_imem_bits_mask = io_imem_resp_bits_mask;
    assign _ibuf__io_imem_bits_pc = io_imem_resp_bits_pc;
    assign _ibuf__io_imem_bits_replay = io_imem_resp_bits_replay;
    assign _ibuf__io_imem_bits_xcpt_if = io_imem_resp_bits_xcpt_if;
    assign _ibuf__io_imem_valid = io_imem_resp_valid;
    assign _ibuf__io_inst_0_ready = _T_4444;
    assign _ibuf__io_kill = take_pc;
    assign _ibuf__reset = reset;
    assign id_ctrl_alu_dw = _T_2997;
    assign id_ctrl_alu_fn = _T_3081;
    assign id_ctrl_amo = _T_3310;
    assign id_ctrl_branch = _T_2821;
    assign id_ctrl_csr = _T_3292;
    assign id_ctrl_div = _T_3236;
    assign id_ctrl_dp = _T_3326;
    assign id_ctrl_fence = _T_3304;
    assign id_ctrl_fence_i = _T_3298;
    assign id_ctrl_fp = _T_2814;
    assign id_ctrl_jal = _T_2827;
    assign id_ctrl_jalr = _T_2833;
    assign id_ctrl_legal = _T_2803;
    assign id_ctrl_mem = _T_3102;
    assign id_ctrl_mem_cmd = _T_3162;
    assign id_ctrl_mem_type = _T_3182;
    assign id_ctrl_rfs1 = _T_3198;
    assign id_ctrl_rfs2 = _T_3215;
    assign id_ctrl_rfs3 = _T_3217;
    assign id_ctrl_rocc = 1'h0;
    assign id_ctrl_rxs1 = _T_2880;
    assign id_ctrl_rxs2 = _T_2854;
    assign id_ctrl_sel_alu1 = _T_2950;
    assign id_ctrl_sel_alu2 = _T_2924;
    assign id_ctrl_sel_imm = _T_2986;
    assign id_ctrl_wfd = _T_3230;
    assign id_ctrl_wxd = _T_3272;
    assign id_load_use = _T_4325;
    assign _WTEMP_114 = _T_3512;
    MUX_UNSIGNED #(.width(64)) u_mux_5741 (
        .y(id_rs_0),
        .sel(rf_wen),
        .a(_node_390),
        .b(_T_3341)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_5742 (
        .y(id_rs_1),
        .sel(rf_wen),
        .a(_node_391),
        .b(_T_3351)
    );
    assign io_dmem_invalidate_lr = _wb_reg_xcpt__q;
    assign io_dmem_req_bits_addr = _T_4518;
    assign io_dmem_req_bits_cmd = _ex_ctrl_mem_cmd__q;
    assign io_dmem_req_bits_data = 64'h0;
    assign io_dmem_req_bits_phys = 1'h0;
    PAD_UNSIGNED #(.width(6), .n(7)) u_pad_5743 (
        .y(io_dmem_req_bits_tag),
        .in(ex_dcache_tag)
    );
    assign io_dmem_req_bits_typ = _ex_ctrl_mem_type__q;
    assign io_dmem_req_valid = _T_4493;
    assign io_dmem_s1_data = _T_4519;
    assign io_dmem_s1_kill = _T_4520;
    assign io_fpu_dmem_resp_data = io_dmem_resp_bits_data_word_bypass;
    assign io_fpu_dmem_resp_tag = dmem_resp_waddr;
    assign io_fpu_dmem_resp_type = io_dmem_resp_bits_typ;
    assign io_fpu_dmem_resp_val = _T_4492;
    assign io_fpu_fcsr_rm = _csr__io_fcsr_rm;
    assign io_fpu_fromint_data = ex_rs_0;
    assign io_fpu_inst = _ibuf__io_inst_0_bits_inst_bits;
    assign io_fpu_killm = killm_common;
    assign io_fpu_killx = ctrl_killx;
    assign io_fpu_valid = _T_4491;
    assign io_imem_bht_update_bits_mispredict = mem_misprediction;
    assign io_imem_bht_update_bits_pc = io_imem_btb_update_bits_pc;
    assign io_imem_bht_update_bits_prediction_bits_bht_history = io_imem_btb_update_bits_prediction_bits_bht_history;
    assign io_imem_bht_update_bits_prediction_bits_bht_value = io_imem_btb_update_bits_prediction_bits_bht_value;
    assign io_imem_bht_update_bits_prediction_bits_bridx = io_imem_btb_update_bits_prediction_bits_bridx;
    assign io_imem_bht_update_bits_prediction_bits_entry = io_imem_btb_update_bits_prediction_bits_entry;
    assign io_imem_bht_update_bits_prediction_bits_mask = io_imem_btb_update_bits_prediction_bits_mask;
    assign io_imem_bht_update_bits_prediction_bits_taken = io_imem_btb_update_bits_prediction_bits_taken;
    assign io_imem_bht_update_bits_prediction_bits_target = io_imem_btb_update_bits_prediction_bits_target;
    assign io_imem_bht_update_bits_prediction_valid = io_imem_btb_update_bits_prediction_valid;
    assign io_imem_bht_update_bits_taken = mem_br_taken;
    assign io_imem_bht_update_valid = _T_4483;
    BITS #(.width(40), .high(38), .low(0)) bits_5744 (
        .y(io_imem_btb_update_bits_br_pc),
        .in(_T_4475)
    );
    assign io_imem_btb_update_bits_isJump = _T_4464;
    assign io_imem_btb_update_bits_isReturn = _T_4470;
    assign io_imem_btb_update_bits_isValid = _T_4463;
    assign io_imem_btb_update_bits_pc = _T_4479;
    assign io_imem_btb_update_bits_prediction_bits_bht_history = _mem_reg_btb_resp_bht_history__q;
    assign io_imem_btb_update_bits_prediction_bits_bht_value = _mem_reg_btb_resp_bht_value__q;
    assign io_imem_btb_update_bits_prediction_bits_bridx = _mem_reg_btb_resp_bridx__q;
    assign io_imem_btb_update_bits_prediction_bits_entry = _mem_reg_btb_resp_entry__q;
    assign io_imem_btb_update_bits_prediction_bits_mask = _mem_reg_btb_resp_mask__q;
    assign io_imem_btb_update_bits_prediction_bits_taken = _mem_reg_btb_resp_taken__q;
    assign io_imem_btb_update_bits_prediction_bits_target = _mem_reg_btb_resp_target__q;
    assign io_imem_btb_update_bits_prediction_valid = _mem_reg_btb_hit__q;
    assign io_imem_btb_update_bits_taken = 1'h0;
    BITS #(.width(40), .high(38), .low(0)) bits_5745 (
        .y(io_imem_btb_update_bits_target),
        .in(io_imem_req_bits_pc)
    );
    assign io_imem_btb_update_valid = _T_4460;
    assign io_imem_flush_icache = _T_4441;
    assign io_imem_flush_tlb = _csr__io_fatc;
    assign io_imem_ras_update_bits_isCall = _T_4488;
    assign io_imem_ras_update_bits_isReturn = io_imem_btb_update_bits_isReturn;
    assign io_imem_ras_update_bits_prediction_bits_bht_history = io_imem_btb_update_bits_prediction_bits_bht_history;
    assign io_imem_ras_update_bits_prediction_bits_bht_value = io_imem_btb_update_bits_prediction_bits_bht_value;
    assign io_imem_ras_update_bits_prediction_bits_bridx = io_imem_btb_update_bits_prediction_bits_bridx;
    assign io_imem_ras_update_bits_prediction_bits_entry = io_imem_btb_update_bits_prediction_bits_entry;
    assign io_imem_ras_update_bits_prediction_bits_mask = io_imem_btb_update_bits_prediction_bits_mask;
    assign io_imem_ras_update_bits_prediction_bits_taken = io_imem_btb_update_bits_prediction_bits_taken;
    assign io_imem_ras_update_bits_prediction_bits_target = io_imem_btb_update_bits_prediction_bits_target;
    assign io_imem_ras_update_bits_prediction_valid = io_imem_btb_update_bits_prediction_valid;
    BITS #(.width(64), .high(38), .low(0)) bits_5746 (
        .y(io_imem_ras_update_bits_returnAddr),
        .in(mem_int_wdata)
    );
    assign io_imem_ras_update_valid = _T_4486;
    assign io_imem_req_bits_pc = _T_4437;
    assign io_imem_req_bits_speculative = _T_4431;
    assign io_imem_req_valid = take_pc;
    assign io_imem_resp_ready = _ibuf__io_imem_ready;
    assign io_ptw_invalidate = _csr__io_fatc;
    assign io_ptw_ptbr_asid = _csr__io_ptbr_asid;
    assign io_ptw_ptbr_mode = _csr__io_ptbr_mode;
    assign io_ptw_ptbr_ppn = _csr__io_ptbr_ppn;
    assign io_ptw_status_debug = _csr__io_status_debug;
    assign io_ptw_status_fs = _csr__io_status_fs;
    assign io_ptw_status_hie = _csr__io_status_hie;
    assign io_ptw_status_hpie = _csr__io_status_hpie;
    assign io_ptw_status_hpp = _csr__io_status_hpp;
    assign io_ptw_status_isa = _csr__io_status_isa;
    assign io_ptw_status_mie = _csr__io_status_mie;
    assign io_ptw_status_mpie = _csr__io_status_mpie;
    assign io_ptw_status_mpp = _csr__io_status_mpp;
    assign io_ptw_status_mprv = _csr__io_status_mprv;
    assign io_ptw_status_mxr = _csr__io_status_mxr;
    assign io_ptw_status_prv = _csr__io_status_prv;
    assign io_ptw_status_pum = _csr__io_status_pum;
    assign io_ptw_status_sd = _csr__io_status_sd;
    assign io_ptw_status_sd_rv32 = _csr__io_status_sd_rv32;
    assign io_ptw_status_sie = _csr__io_status_sie;
    assign io_ptw_status_spie = _csr__io_status_spie;
    assign io_ptw_status_spp = _csr__io_status_spp;
    assign io_ptw_status_sxl = _csr__io_status_sxl;
    assign io_ptw_status_tsr = _csr__io_status_tsr;
    assign io_ptw_status_tvm = _csr__io_status_tvm;
    assign io_ptw_status_tw = _csr__io_status_tw;
    assign io_ptw_status_uie = _csr__io_status_uie;
    assign io_ptw_status_upie = _csr__io_status_upie;
    assign io_ptw_status_uxl = _csr__io_status_uxl;
    assign io_ptw_status_xs = _csr__io_status_xs;
    assign io_ptw_status_zero1 = _csr__io_status_zero1;
    assign io_ptw_status_zero2 = _csr__io_status_zero2;
    assign io_rocc_cmd_bits_inst_funct = _T_4558_funct;
    assign io_rocc_cmd_bits_inst_opcode = _T_4558_opcode;
    assign io_rocc_cmd_bits_inst_rd = _T_4558_rd;
    assign io_rocc_cmd_bits_inst_rs1 = _T_4558_rs1;
    assign io_rocc_cmd_bits_inst_rs2 = _T_4558_rs2;
    assign io_rocc_cmd_bits_inst_xd = _T_4558_xd;
    assign io_rocc_cmd_bits_inst_xs1 = _T_4558_xs1;
    assign io_rocc_cmd_bits_inst_xs2 = _T_4558_xs2;
    assign io_rocc_cmd_bits_rs1 = _wb_reg_wdata__q;
    assign io_rocc_cmd_bits_rs2 = 64'h0;
    assign io_rocc_cmd_bits_status_debug = _csr__io_status_debug;
    assign io_rocc_cmd_bits_status_fs = _csr__io_status_fs;
    assign io_rocc_cmd_bits_status_hie = _csr__io_status_hie;
    assign io_rocc_cmd_bits_status_hpie = _csr__io_status_hpie;
    assign io_rocc_cmd_bits_status_hpp = _csr__io_status_hpp;
    assign io_rocc_cmd_bits_status_isa = _csr__io_status_isa;
    assign io_rocc_cmd_bits_status_mie = _csr__io_status_mie;
    assign io_rocc_cmd_bits_status_mpie = _csr__io_status_mpie;
    assign io_rocc_cmd_bits_status_mpp = _csr__io_status_mpp;
    assign io_rocc_cmd_bits_status_mprv = _csr__io_status_mprv;
    assign io_rocc_cmd_bits_status_mxr = _csr__io_status_mxr;
    assign io_rocc_cmd_bits_status_prv = _csr__io_status_prv;
    assign io_rocc_cmd_bits_status_pum = _csr__io_status_pum;
    assign io_rocc_cmd_bits_status_sd = _csr__io_status_sd;
    assign io_rocc_cmd_bits_status_sd_rv32 = _csr__io_status_sd_rv32;
    assign io_rocc_cmd_bits_status_sie = _csr__io_status_sie;
    assign io_rocc_cmd_bits_status_spie = _csr__io_status_spie;
    assign io_rocc_cmd_bits_status_spp = _csr__io_status_spp;
    assign io_rocc_cmd_bits_status_sxl = _csr__io_status_sxl;
    assign io_rocc_cmd_bits_status_tsr = _csr__io_status_tsr;
    assign io_rocc_cmd_bits_status_tvm = _csr__io_status_tvm;
    assign io_rocc_cmd_bits_status_tw = _csr__io_status_tw;
    assign io_rocc_cmd_bits_status_uie = _csr__io_status_uie;
    assign io_rocc_cmd_bits_status_upie = _csr__io_status_upie;
    assign io_rocc_cmd_bits_status_uxl = _csr__io_status_uxl;
    assign io_rocc_cmd_bits_status_xs = _csr__io_status_xs;
    assign io_rocc_cmd_bits_status_zero1 = _csr__io_status_zero1;
    assign io_rocc_cmd_bits_status_zero2 = _csr__io_status_zero2;
    assign io_rocc_cmd_valid = 1'h0;
    assign io_rocc_exception = _T_4539;
    assign io_rocc_mem_acquire = 1'h0;
    assign io_rocc_mem_ordered = 1'h0;
    assign io_rocc_mem_release = 1'h0;
    assign io_rocc_mem_replay_next = 1'h0;
    assign io_rocc_mem_req_ready = 1'h0;
    assign io_rocc_mem_resp_bits_addr = 40'h0;
    assign io_rocc_mem_resp_bits_cmd = 5'h0;
    assign io_rocc_mem_resp_bits_data = 64'h0;
    assign io_rocc_mem_resp_bits_data_word_bypass = 64'h0;
    assign io_rocc_mem_resp_bits_has_data = 1'h0;
    assign io_rocc_mem_resp_bits_replay = 1'h0;
    assign io_rocc_mem_resp_bits_store_data = 64'h0;
    assign io_rocc_mem_resp_bits_tag = 7'h0;
    assign io_rocc_mem_resp_bits_typ = 3'h0;
    assign io_rocc_mem_resp_valid = 1'h0;
    assign io_rocc_mem_s2_nack = 1'h0;
    assign io_rocc_mem_xcpt_ma_ld = 1'h0;
    assign io_rocc_mem_xcpt_ma_st = 1'h0;
    assign io_rocc_mem_xcpt_pf_ld = 1'h0;
    assign io_rocc_mem_xcpt_pf_st = 1'h0;
    assign io_rocc_resp_ready = 1'h0;
    MUX_UNSIGNED #(.width(5)) u_mux_5747 (
        .y(ll_waddr),
        .sel(_T_4183),
        .a(dmem_resp_waddr),
        .b(_div__io_resp_bits_tag)
    );
    assign ll_wdata = _div__io_resp_bits_data;
    MUX_UNSIGNED #(.width(1)) u_mux_5748 (
        .y(ll_wen),
        .sel(_T_4183),
        .a(1'h1),
        .b(_T_4182)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_5749 (
        .y(_mem_ctrl_branch__d),
        .sel(ex_pc_valid),
        .a(_ex_ctrl_branch__q),
        .b(_mem_ctrl_branch__q)
    );
    MUX_UNSIGNED #(.width(3)) u_mux_5750 (
        .y(_mem_ctrl_csr__d),
        .sel(ex_pc_valid),
        .a(_ex_ctrl_csr__q),
        .b(_mem_ctrl_csr__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_5751 (
        .y(_mem_ctrl_div__d),
        .sel(ex_pc_valid),
        .a(_ex_ctrl_div__q),
        .b(_mem_ctrl_div__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_5752 (
        .y(_mem_ctrl_fence_i__d),
        .sel(ex_pc_valid),
        .a(_ex_ctrl_fence_i__q),
        .b(_mem_ctrl_fence_i__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_5753 (
        .y(_mem_ctrl_fp__d),
        .sel(ex_pc_valid),
        .a(_ex_ctrl_fp__q),
        .b(_mem_ctrl_fp__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_5754 (
        .y(_mem_ctrl_jal__d),
        .sel(ex_pc_valid),
        .a(_ex_ctrl_jal__q),
        .b(_mem_ctrl_jal__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_5755 (
        .y(_mem_ctrl_jalr__d),
        .sel(ex_pc_valid),
        .a(_ex_ctrl_jalr__q),
        .b(_mem_ctrl_jalr__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_5756 (
        .y(_mem_ctrl_mem__d),
        .sel(ex_pc_valid),
        .a(_ex_ctrl_mem__q),
        .b(_mem_ctrl_mem__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_5757 (
        .y(_mem_ctrl_wfd__d),
        .sel(ex_pc_valid),
        .a(_ex_ctrl_wfd__q),
        .b(_mem_ctrl_wfd__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_5758 (
        .y(_mem_ctrl_wxd__d),
        .sel(ex_pc_valid),
        .a(_ex_ctrl_wxd__q),
        .b(_mem_ctrl_wxd__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_5759 (
        .y(_mem_reg_btb_hit__d),
        .sel(ex_pc_valid),
        .a(_ex_reg_btb_hit__q),
        .b(_mem_reg_btb_hit__q)
    );
    MUX_UNSIGNED #(.width(7)) u_mux_5760 (
        .y(_mem_reg_btb_resp_bht_history__d),
        .sel(ex_pc_valid),
        .a(_node_377),
        .b(_mem_reg_btb_resp_bht_history__q)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_5761 (
        .y(_mem_reg_btb_resp_bht_value__d),
        .sel(ex_pc_valid),
        .a(_node_378),
        .b(_mem_reg_btb_resp_bht_value__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_5762 (
        .y(_mem_reg_btb_resp_bridx__d),
        .sel(ex_pc_valid),
        .a(_node_379),
        .b(_mem_reg_btb_resp_bridx__q)
    );
    MUX_UNSIGNED #(.width(6)) u_mux_5763 (
        .y(_mem_reg_btb_resp_entry__d),
        .sel(ex_pc_valid),
        .a(_node_380),
        .b(_mem_reg_btb_resp_entry__q)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_5764 (
        .y(_mem_reg_btb_resp_mask__d),
        .sel(ex_pc_valid),
        .a(_node_381),
        .b(_mem_reg_btb_resp_mask__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_5765 (
        .y(_mem_reg_btb_resp_taken__d),
        .sel(ex_pc_valid),
        .a(_node_382),
        .b(_mem_reg_btb_resp_taken__q)
    );
    MUX_UNSIGNED #(.width(39)) u_mux_5766 (
        .y(_mem_reg_btb_resp_target__d),
        .sel(ex_pc_valid),
        .a(_node_383),
        .b(_mem_reg_btb_resp_target__q)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_5767 (
        .y(_mem_reg_cause__d),
        .sel(ex_xcpt),
        .a(_ex_cause__q),
        .b(_mem_reg_cause__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_5768 (
        .y(_mem_reg_flush_pipe__d),
        .sel(ex_pc_valid),
        .a(_ex_reg_flush_pipe__q),
        .b(_mem_reg_flush_pipe__q)
    );
    MUX_UNSIGNED #(.width(32)) u_mux_5769 (
        .y(_mem_reg_inst__d),
        .sel(ex_pc_valid),
        .a(_ex_reg_inst__q),
        .b(_mem_reg_inst__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_5770 (
        .y(_mem_reg_load__d),
        .sel(ex_pc_valid),
        .a(_T_4077),
        .b(_mem_reg_load__q)
    );
    MUX_UNSIGNED #(.width(40)) u_mux_5771 (
        .y(_mem_reg_pc__d),
        .sel(ex_pc_valid),
        .a(_ex_reg_pc__q),
        .b(_mem_reg_pc__q)
    );
    assign _mem_reg_replay__d = _T_4057;
    MUX_UNSIGNED #(.width(64)) u_mux_5772 (
        .y(_mem_reg_rs2__d),
        .sel(ex_pc_valid),
        .a(_node_384),
        .b(_mem_reg_rs2__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_5773 (
        .y(_mem_reg_rvc__d),
        .sel(ex_pc_valid),
        .a(_ex_reg_rvc__q),
        .b(_mem_reg_rvc__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_5774 (
        .y(_mem_reg_slow_bypass__d),
        .sel(ex_pc_valid),
        .a(ex_slow_bypass),
        .b(_mem_reg_slow_bypass__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_5775 (
        .y(_mem_reg_store__d),
        .sel(ex_pc_valid),
        .a(_T_4088),
        .b(_mem_reg_store__q)
    );
    assign _mem_reg_valid__d = _T_4054;
    MUX_UNSIGNED #(.width(64)) u_mux_5776 (
        .y(_mem_reg_wdata__d),
        .sel(ex_pc_valid),
        .a(_alu__io_out),
        .b(_mem_reg_wdata__q)
    );
    assign _mem_reg_xcpt__d = _T_4060;
    assign _mem_reg_xcpt_interrupt__d = _T_4063;
    assign _rocc_blocked__d = _T_4404;
    assign take_pc_id = 1'h0;
    assign take_pc_mem = _T_4052;
    assign take_pc_wb = _T_4175;
    MUX_UNSIGNED #(.width(3)) u_mux_5777 (
        .y(_wb_ctrl_csr__d),
        .sel(mem_pc_valid),
        .a(_mem_ctrl_csr__q),
        .b(_wb_ctrl_csr__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_5778 (
        .y(_wb_ctrl_div__d),
        .sel(mem_pc_valid),
        .a(_mem_ctrl_div__q),
        .b(_wb_ctrl_div__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_5779 (
        .y(_wb_ctrl_fence_i__d),
        .sel(mem_pc_valid),
        .a(_mem_ctrl_fence_i__q),
        .b(_wb_ctrl_fence_i__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_5780 (
        .y(_wb_ctrl_mem__d),
        .sel(mem_pc_valid),
        .a(_mem_ctrl_mem__q),
        .b(_wb_ctrl_mem__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_5781 (
        .y(_wb_ctrl_wfd__d),
        .sel(mem_pc_valid),
        .a(_mem_ctrl_wfd__q),
        .b(_wb_ctrl_wfd__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_5782 (
        .y(_wb_ctrl_wxd__d),
        .sel(mem_pc_valid),
        .a(_mem_ctrl_wxd__q),
        .b(_wb_ctrl_wxd__q)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_5783 (
        .y(_wb_reg_cause__d),
        .sel(mem_xcpt),
        .a(mem_cause),
        .b(_wb_reg_cause__q)
    );
    MUX_UNSIGNED #(.width(32)) u_mux_5784 (
        .y(_wb_reg_inst__d),
        .sel(mem_pc_valid),
        .a(_mem_reg_inst__q),
        .b(_wb_reg_inst__q)
    );
    MUX_UNSIGNED #(.width(40)) u_mux_5785 (
        .y(_wb_reg_pc__d),
        .sel(mem_pc_valid),
        .a(_mem_reg_pc__q),
        .b(_wb_reg_pc__q)
    );
    assign _wb_reg_replay__d = _T_4161;
    assign _wb_reg_valid__d = _T_4158;
    MUX_UNSIGNED #(.width(64)) u_mux_5786 (
        .y(_wb_reg_wdata__d),
        .sel(mem_pc_valid),
        .a(_T_4169),
        .b(_wb_reg_wdata__q)
    );
    assign _wb_reg_xcpt__d = _T_4164;
endmodule //RocketCore
module DFF_POSCLK(q, d, clk);
    parameter width = 4;
    output reg [width-1:0] q;
    input [width-1:0] d;
    input clk;
    always @(posedge clk) begin
        q <= d;
    end
endmodule // DFF_POSCLK
module BITWISEOR(y, a, b);
    parameter width = 4;
    output [width-1:0] y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a | b;
endmodule // BITWISEOR
module IBuf(
    input clock,
    input reset,
    output io_imem_ready,
    input io_imem_valid,
    input io_imem_bits_btb_valid,
    input io_imem_bits_btb_bits_taken,
    input [1:0] io_imem_bits_btb_bits_mask,
    input io_imem_bits_btb_bits_bridx,
    input [38:0] io_imem_bits_btb_bits_target,
    input [5:0] io_imem_bits_btb_bits_entry,
    input [6:0] io_imem_bits_btb_bits_bht_history,
    input [1:0] io_imem_bits_btb_bits_bht_value,
    input [39:0] io_imem_bits_pc,
    input [31:0] io_imem_bits_data,
    input [1:0] io_imem_bits_mask,
    input io_imem_bits_xcpt_if,
    input io_imem_bits_replay,
    input io_kill,
    output [39:0] io_pc,
    output io_btb_resp_taken,
    output [1:0] io_btb_resp_mask,
    output io_btb_resp_bridx,
    output [38:0] io_btb_resp_target,
    output [5:0] io_btb_resp_entry,
    output [6:0] io_btb_resp_bht_history,
    output [1:0] io_btb_resp_bht_value,
    input io_inst_0_ready,
    output io_inst_0_valid,
    output io_inst_0_bits_pf0,
    output io_inst_0_bits_pf1,
    output io_inst_0_bits_replay,
    output io_inst_0_bits_btb_hit,
    output io_inst_0_bits_rvc,
    output [31:0] io_inst_0_bits_inst_bits,
    output [4:0] io_inst_0_bits_inst_rd,
    output [4:0] io_inst_0_bits_inst_rs1,
    output [4:0] io_inst_0_bits_inst_rs2,
    output [4:0] io_inst_0_bits_inst_rs3,
    output [31:0] io_inst_0_bits_raw
);
    wire _nBufValid__q;
    wire _nBufValid__d;
    DFF_POSCLK #(.width(1)) nBufValid (
        .q(_nBufValid__q),
        .d(_nBufValid__d),
        .clk(clock)
    );
    wire _WTEMP_0;
    MUX_UNSIGNED #(.width(1)) u_mux_3 (
        .y(_nBufValid__d),
        .sel(reset),
        .a(1'h0),
        .b(_WTEMP_0)
    );
    wire _buf_btb_valid__q;
    wire _buf_btb_valid__d;
    DFF_POSCLK #(.width(1)) buf_btb_valid (
        .q(_buf_btb_valid__q),
        .d(_buf_btb_valid__d),
        .clk(clock)
    );
    wire _buf_btb_bits_taken__q;
    wire _buf_btb_bits_taken__d;
    DFF_POSCLK #(.width(1)) buf_btb_bits_taken (
        .q(_buf_btb_bits_taken__q),
        .d(_buf_btb_bits_taken__d),
        .clk(clock)
    );
    wire [1:0] _buf_btb_bits_mask__q;
    wire [1:0] _buf_btb_bits_mask__d;
    DFF_POSCLK #(.width(2)) buf_btb_bits_mask (
        .q(_buf_btb_bits_mask__q),
        .d(_buf_btb_bits_mask__d),
        .clk(clock)
    );
    wire _buf_btb_bits_bridx__q;
    wire _buf_btb_bits_bridx__d;
    DFF_POSCLK #(.width(1)) buf_btb_bits_bridx (
        .q(_buf_btb_bits_bridx__q),
        .d(_buf_btb_bits_bridx__d),
        .clk(clock)
    );
    wire [38:0] _buf_btb_bits_target__q;
    wire [38:0] _buf_btb_bits_target__d;
    DFF_POSCLK #(.width(39)) buf_btb_bits_target (
        .q(_buf_btb_bits_target__q),
        .d(_buf_btb_bits_target__d),
        .clk(clock)
    );
    wire [5:0] _buf_btb_bits_entry__q;
    wire [5:0] _buf_btb_bits_entry__d;
    DFF_POSCLK #(.width(6)) buf_btb_bits_entry (
        .q(_buf_btb_bits_entry__q),
        .d(_buf_btb_bits_entry__d),
        .clk(clock)
    );
    wire [6:0] _buf_btb_bits_bht_history__q;
    wire [6:0] _buf_btb_bits_bht_history__d;
    DFF_POSCLK #(.width(7)) buf_btb_bits_bht_history (
        .q(_buf_btb_bits_bht_history__q),
        .d(_buf_btb_bits_bht_history__d),
        .clk(clock)
    );
    wire [1:0] _buf_btb_bits_bht_value__q;
    wire [1:0] _buf_btb_bits_bht_value__d;
    DFF_POSCLK #(.width(2)) buf_btb_bits_bht_value (
        .q(_buf_btb_bits_bht_value__q),
        .d(_buf_btb_bits_bht_value__d),
        .clk(clock)
    );
    wire [39:0] _buf_pc__q;
    wire [39:0] _buf_pc__d;
    DFF_POSCLK #(.width(40)) buf_pc (
        .q(_buf_pc__q),
        .d(_buf_pc__d),
        .clk(clock)
    );
    wire [31:0] _buf_data__q;
    wire [31:0] _buf_data__d;
    DFF_POSCLK #(.width(32)) buf_data (
        .q(_buf_data__q),
        .d(_buf_data__d),
        .clk(clock)
    );
    wire [1:0] _buf_mask__q;
    wire [1:0] _buf_mask__d;
    DFF_POSCLK #(.width(2)) buf_mask (
        .q(_buf_mask__q),
        .d(_buf_mask__d),
        .clk(clock)
    );
    wire _buf_xcpt_if__q;
    wire _buf_xcpt_if__d;
    DFF_POSCLK #(.width(1)) buf_xcpt_if (
        .q(_buf_xcpt_if__q),
        .d(_buf_xcpt_if__d),
        .clk(clock)
    );
    wire _buf_replay__q;
    wire _buf_replay__d;
    DFF_POSCLK #(.width(1)) buf_replay (
        .q(_buf_replay__q),
        .d(_buf_replay__d),
        .clk(clock)
    );
    wire _ibufBTBHit__q;
    wire _ibufBTBHit__d;
    DFF_POSCLK #(.width(1)) ibufBTBHit (
        .q(_ibufBTBHit__q),
        .d(_ibufBTBHit__d),
        .clk(clock)
    );
    wire _ibufBTBResp_taken__q;
    wire _ibufBTBResp_taken__d;
    DFF_POSCLK #(.width(1)) ibufBTBResp_taken (
        .q(_ibufBTBResp_taken__q),
        .d(_ibufBTBResp_taken__d),
        .clk(clock)
    );
    wire [1:0] _ibufBTBResp_mask__q;
    wire [1:0] _ibufBTBResp_mask__d;
    DFF_POSCLK #(.width(2)) ibufBTBResp_mask (
        .q(_ibufBTBResp_mask__q),
        .d(_ibufBTBResp_mask__d),
        .clk(clock)
    );
    wire _ibufBTBResp_bridx__q;
    wire _ibufBTBResp_bridx__d;
    DFF_POSCLK #(.width(1)) ibufBTBResp_bridx (
        .q(_ibufBTBResp_bridx__q),
        .d(_ibufBTBResp_bridx__d),
        .clk(clock)
    );
    wire [38:0] _ibufBTBResp_target__q;
    wire [38:0] _ibufBTBResp_target__d;
    DFF_POSCLK #(.width(39)) ibufBTBResp_target (
        .q(_ibufBTBResp_target__q),
        .d(_ibufBTBResp_target__d),
        .clk(clock)
    );
    wire [5:0] _ibufBTBResp_entry__q;
    wire [5:0] _ibufBTBResp_entry__d;
    DFF_POSCLK #(.width(6)) ibufBTBResp_entry (
        .q(_ibufBTBResp_entry__q),
        .d(_ibufBTBResp_entry__d),
        .clk(clock)
    );
    wire [6:0] _ibufBTBResp_bht_history__q;
    wire [6:0] _ibufBTBResp_bht_history__d;
    DFF_POSCLK #(.width(7)) ibufBTBResp_bht_history (
        .q(_ibufBTBResp_bht_history__q),
        .d(_ibufBTBResp_bht_history__d),
        .clk(clock)
    );
    wire [1:0] _ibufBTBResp_bht_value__q;
    wire [1:0] _ibufBTBResp_bht_value__d;
    DFF_POSCLK #(.width(2)) ibufBTBResp_bht_value (
        .q(_ibufBTBResp_bht_value__q),
        .d(_ibufBTBResp_bht_value__d),
        .clk(clock)
    );
    wire pcWordBits;
    BITS #(.width(40), .high(1), .low(1)) bits_4 (
        .y(pcWordBits),
        .in(io_imem_bits_pc)
    );
    wire [1:0] nReady;
    wire _T_375;
    BITWISEAND #(.width(1)) bitwiseand_5 (
        .y(_T_375),
        .a(io_imem_bits_btb_valid),
        .b(io_imem_bits_btb_bits_taken)
    );
    wire [1:0] _T_377;
    ADD_UNSIGNED #(.width(1)) u_add_6 (
        .y(_T_377),
        .a(io_imem_bits_btb_bits_bridx),
        .b(1'h1)
    );
    wire [1:0] _T_379;
    MUX_UNSIGNED #(.width(2)) u_mux_7 (
        .y(_T_379),
        .sel(_T_375),
        .a(_T_377),
        .b(2'h2)
    );
    wire [2:0] _T_380;
    wire [1:0] _WTEMP_1;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_8 (
        .y(_WTEMP_1),
        .in(pcWordBits)
    );
    SUB_UNSIGNED #(.width(2)) u_sub_9 (
        .y(_T_380),
        .a(_T_379),
        .b(_WTEMP_1)
    );
    wire [2:0] _T_381;
    ASUINT #(.width(3)) asuint_10 (
        .y(_T_381),
        .in(_T_380)
    );
    wire [1:0] nIC;
    TAIL #(.width(3), .n(1)) tail_11 (
        .y(nIC),
        .in(_T_381)
    );
    wire [2:0] _T_382;
    wire [1:0] _WTEMP_2;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_12 (
        .y(_WTEMP_2),
        .in(_nBufValid__q)
    );
    SUB_UNSIGNED #(.width(2)) u_sub_13 (
        .y(_T_382),
        .a(nReady),
        .b(_WTEMP_2)
    );
    wire [2:0] _T_383;
    ASUINT #(.width(3)) asuint_14 (
        .y(_T_383),
        .in(_T_382)
    );
    wire [1:0] nICReady;
    TAIL #(.width(3), .n(1)) tail_15 (
        .y(nICReady),
        .in(_T_383)
    );
    wire [1:0] _T_385;
    wire [1:0] _WTEMP_3;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_16 (
        .y(_WTEMP_3),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_17 (
        .y(_T_385),
        .sel(io_imem_valid),
        .a(nIC),
        .b(_WTEMP_3)
    );
    wire [2:0] _T_386;
    wire [1:0] _WTEMP_4;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_18 (
        .y(_WTEMP_4),
        .in(_nBufValid__q)
    );
    ADD_UNSIGNED #(.width(2)) u_add_19 (
        .y(_T_386),
        .a(_T_385),
        .b(_WTEMP_4)
    );
    wire [1:0] nValid;
    TAIL #(.width(3), .n(1)) tail_20 (
        .y(nValid),
        .in(_T_386)
    );
    wire _T_387;
    wire [1:0] _WTEMP_5;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_21 (
        .y(_WTEMP_5),
        .in(_nBufValid__q)
    );
    GEQ_UNSIGNED #(.width(2)) u_geq_22 (
        .y(_T_387),
        .a(nReady),
        .b(_WTEMP_5)
    );
    wire _T_388;
    GEQ_UNSIGNED #(.width(2)) u_geq_23 (
        .y(_T_388),
        .a(nICReady),
        .b(nIC)
    );
    wire [2:0] _T_390;
    SUB_UNSIGNED #(.width(2)) u_sub_24 (
        .y(_T_390),
        .a(nIC),
        .b(nICReady)
    );
    wire [2:0] _T_391;
    ASUINT #(.width(3)) asuint_25 (
        .y(_T_391),
        .in(_T_390)
    );
    wire [1:0] _T_392;
    TAIL #(.width(3), .n(1)) tail_26 (
        .y(_T_392),
        .in(_T_391)
    );
    wire _T_393;
    wire [1:0] _WTEMP_6;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_27 (
        .y(_WTEMP_6),
        .in(1'h1)
    );
    GEQ_UNSIGNED #(.width(2)) u_geq_28 (
        .y(_T_393),
        .a(_WTEMP_6),
        .b(_T_392)
    );
    wire _T_394;
    BITWISEOR #(.width(1)) bitwiseor_29 (
        .y(_T_394),
        .a(_T_388),
        .b(_T_393)
    );
    wire _T_395;
    BITWISEAND #(.width(1)) bitwiseand_30 (
        .y(_T_395),
        .a(_T_387),
        .b(_T_394)
    );
    wire _T_396;
    wire [1:0] _WTEMP_7;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_31 (
        .y(_WTEMP_7),
        .in(_nBufValid__q)
    );
    GEQ_UNSIGNED #(.width(2)) u_geq_32 (
        .y(_T_396),
        .a(nReady),
        .b(_WTEMP_7)
    );
    wire [2:0] _T_398;
    wire [1:0] _WTEMP_8;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_33 (
        .y(_WTEMP_8),
        .in(_nBufValid__q)
    );
    SUB_UNSIGNED #(.width(2)) u_sub_34 (
        .y(_T_398),
        .a(_WTEMP_8),
        .b(nReady)
    );
    wire [2:0] _T_399;
    ASUINT #(.width(3)) asuint_35 (
        .y(_T_399),
        .in(_T_398)
    );
    wire [1:0] _T_400;
    TAIL #(.width(3), .n(1)) tail_36 (
        .y(_T_400),
        .in(_T_399)
    );
    wire [1:0] _T_401;
    wire [1:0] _WTEMP_9;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_37 (
        .y(_WTEMP_9),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_38 (
        .y(_T_401),
        .sel(_T_396),
        .a(_WTEMP_9),
        .b(_T_400)
    );
    wire _T_402;
    wire [1:0] _WTEMP_10;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_39 (
        .y(_WTEMP_10),
        .in(_nBufValid__q)
    );
    GEQ_UNSIGNED #(.width(2)) u_geq_40 (
        .y(_T_402),
        .a(nReady),
        .b(_WTEMP_10)
    );
    wire _T_403;
    BITWISEAND #(.width(1)) bitwiseand_41 (
        .y(_T_403),
        .a(io_imem_valid),
        .b(_T_402)
    );
    wire _T_404;
    LT_UNSIGNED #(.width(2)) u_lt_42 (
        .y(_T_404),
        .a(nICReady),
        .b(nIC)
    );
    wire _T_405;
    BITWISEAND #(.width(1)) bitwiseand_43 (
        .y(_T_405),
        .a(_T_403),
        .b(_T_404)
    );
    wire [2:0] _T_407;
    SUB_UNSIGNED #(.width(2)) u_sub_44 (
        .y(_T_407),
        .a(nIC),
        .b(nICReady)
    );
    wire [2:0] _T_408;
    ASUINT #(.width(3)) asuint_45 (
        .y(_T_408),
        .in(_T_407)
    );
    wire [1:0] _T_409;
    TAIL #(.width(3), .n(1)) tail_46 (
        .y(_T_409),
        .in(_T_408)
    );
    wire _T_410;
    wire [1:0] _WTEMP_11;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_47 (
        .y(_WTEMP_11),
        .in(1'h1)
    );
    GEQ_UNSIGNED #(.width(2)) u_geq_48 (
        .y(_T_410),
        .a(_WTEMP_11),
        .b(_T_409)
    );
    wire _T_411;
    BITWISEAND #(.width(1)) bitwiseand_49 (
        .y(_T_411),
        .a(_T_405),
        .b(_T_410)
    );
    wire [2:0] _T_412;
    wire [1:0] _WTEMP_12;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_50 (
        .y(_WTEMP_12),
        .in(pcWordBits)
    );
    ADD_UNSIGNED #(.width(2)) u_add_51 (
        .y(_T_412),
        .a(_WTEMP_12),
        .b(nICReady)
    );
    wire [1:0] _T_413;
    TAIL #(.width(3), .n(1)) tail_52 (
        .y(_T_413),
        .in(_T_412)
    );
    wire [2:0] _T_414;
    SUB_UNSIGNED #(.width(2)) u_sub_53 (
        .y(_T_414),
        .a(nIC),
        .b(nICReady)
    );
    wire [2:0] _T_415;
    ASUINT #(.width(3)) asuint_54 (
        .y(_T_415),
        .in(_T_414)
    );
    wire [1:0] _T_416;
    TAIL #(.width(3), .n(1)) tail_55 (
        .y(_T_416),
        .in(_T_415)
    );
    wire [15:0] _T_417;
    SHR_UNSIGNED #(.width(32), .n(16)) u_shr_56 (
        .y(_T_417),
        .in(io_imem_bits_data)
    );
    wire [31:0] _T_418;
    CAT #(.width_a(16), .width_b(16)) cat_57 (
        .y(_T_418),
        .a(_T_417),
        .b(_T_417)
    );
    wire [63:0] _T_419;
    CAT #(.width_a(32), .width_b(32)) cat_58 (
        .y(_T_419),
        .a(_T_418),
        .b(io_imem_bits_data)
    );
    wire [5:0] _T_420;
    SHL_UNSIGNED #(.width(2), .n(4)) u_shl_59 (
        .y(_T_420),
        .in(_T_413)
    );
    wire [63:0] _T_421;
    DSHR_UNSIGNED #(.width_in(64), .width_n(6)) u_dshr_60 (
        .y(_T_421),
        .in(_T_419),
        .n(_T_420)
    );
    wire [15:0] _T_422;
    BITS #(.width(64), .high(15), .low(0)) bits_61 (
        .y(_T_422),
        .in(_T_421)
    );
    wire [39:0] _T_423;
    assign _T_423 = 40'hFFFFFFFFFC;
    wire [39:0] _T_424;
    BITWISEAND #(.width(40)) bitwiseand_62 (
        .y(_T_424),
        .a(io_imem_bits_pc),
        .b(_T_423)
    );
    wire [2:0] _T_425;
    SHL_UNSIGNED #(.width(2), .n(1)) u_shl_63 (
        .y(_T_425),
        .in(nICReady)
    );
    wire [40:0] _T_426;
    wire [39:0] _WTEMP_13;
    PAD_UNSIGNED #(.width(3), .n(40)) u_pad_64 (
        .y(_WTEMP_13),
        .in(_T_425)
    );
    ADD_UNSIGNED #(.width(40)) u_add_65 (
        .y(_T_426),
        .a(io_imem_bits_pc),
        .b(_WTEMP_13)
    );
    wire [39:0] _T_427;
    TAIL #(.width(41), .n(1)) tail_66 (
        .y(_T_427),
        .in(_T_426)
    );
    wire [39:0] _T_428;
    BITWISEAND #(.width(40)) bitwiseand_67 (
        .y(_T_428),
        .a(_T_427),
        .b(40'h3)
    );
    wire [39:0] _T_429;
    BITWISEOR #(.width(40)) bitwiseor_68 (
        .y(_T_429),
        .a(_T_424),
        .b(_T_428)
    );
    wire [2:0] _T_430;
    wire [1:0] _WTEMP_14;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_69 (
        .y(_WTEMP_14),
        .in(io_imem_bits_btb_bits_bridx)
    );
    ADD_UNSIGNED #(.width(2)) u_add_70 (
        .y(_T_430),
        .a(_WTEMP_14),
        .b(nICReady)
    );
    wire [1:0] _T_431;
    TAIL #(.width(3), .n(1)) tail_71 (
        .y(_T_431),
        .in(_T_430)
    );
    wire [6:0] _node_0;
    MUX_UNSIGNED #(.width(7)) u_mux_72 (
        .y(_node_0),
        .sel(io_imem_bits_btb_valid),
        .a(io_imem_bits_btb_bits_bht_history),
        .b(_ibufBTBResp_bht_history__q)
    );
    wire [1:0] _node_1;
    MUX_UNSIGNED #(.width(2)) u_mux_73 (
        .y(_node_1),
        .sel(io_imem_bits_btb_valid),
        .a(io_imem_bits_btb_bits_bht_value),
        .b(_ibufBTBResp_bht_value__q)
    );
    wire [1:0] _node_2;
    wire [1:0] _WTEMP_15;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_74 (
        .y(_WTEMP_15),
        .in(_ibufBTBResp_bridx__q)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_75 (
        .y(_node_2),
        .sel(io_imem_bits_btb_valid),
        .a(_T_431),
        .b(_WTEMP_15)
    );
    wire [5:0] _node_3;
    MUX_UNSIGNED #(.width(6)) u_mux_76 (
        .y(_node_3),
        .sel(io_imem_bits_btb_valid),
        .a(io_imem_bits_btb_bits_entry),
        .b(_ibufBTBResp_entry__q)
    );
    wire [1:0] _node_4;
    MUX_UNSIGNED #(.width(2)) u_mux_77 (
        .y(_node_4),
        .sel(io_imem_bits_btb_valid),
        .a(io_imem_bits_btb_bits_mask),
        .b(_ibufBTBResp_mask__q)
    );
    wire _node_5;
    MUX_UNSIGNED #(.width(1)) u_mux_78 (
        .y(_node_5),
        .sel(io_imem_bits_btb_valid),
        .a(io_imem_bits_btb_bits_taken),
        .b(_ibufBTBResp_taken__q)
    );
    wire [38:0] _node_6;
    MUX_UNSIGNED #(.width(39)) u_mux_79 (
        .y(_node_6),
        .sel(io_imem_bits_btb_valid),
        .a(io_imem_bits_btb_bits_target),
        .b(_ibufBTBResp_target__q)
    );
    wire [1:0] _node_7;
    MUX_UNSIGNED #(.width(2)) u_mux_80 (
        .y(_node_7),
        .sel(_T_411),
        .a(_T_416),
        .b(_T_401)
    );
    wire [2:0] _T_434;
    wire [1:0] _WTEMP_16;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_81 (
        .y(_WTEMP_16),
        .in(_nBufValid__q)
    );
    ADD_UNSIGNED #(.width(2)) u_add_82 (
        .y(_T_434),
        .a(2'h2),
        .b(_WTEMP_16)
    );
    wire [1:0] _T_435;
    TAIL #(.width(3), .n(1)) tail_83 (
        .y(_T_435),
        .in(_T_434)
    );
    wire [2:0] _T_436;
    wire [1:0] _WTEMP_17;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_84 (
        .y(_WTEMP_17),
        .in(pcWordBits)
    );
    SUB_UNSIGNED #(.width(2)) u_sub_85 (
        .y(_T_436),
        .a(_T_435),
        .b(_WTEMP_17)
    );
    wire [2:0] _T_437;
    ASUINT #(.width(3)) asuint_86 (
        .y(_T_437),
        .in(_T_436)
    );
    wire [1:0] _T_438;
    TAIL #(.width(3), .n(1)) tail_87 (
        .y(_T_438),
        .in(_T_437)
    );
    wire [1:0] icShiftAmt;
    BITS #(.width(2), .high(1), .low(0)) bits_88 (
        .y(icShiftAmt),
        .in(_T_438)
    );
    wire [15:0] _T_439;
    BITS #(.width(32), .high(15), .low(0)) bits_89 (
        .y(_T_439),
        .in(io_imem_bits_data)
    );
    wire [31:0] _T_440;
    CAT #(.width_a(16), .width_b(16)) cat_90 (
        .y(_T_440),
        .a(_T_439),
        .b(_T_439)
    );
    wire [63:0] _T_441;
    CAT #(.width_a(32), .width_b(32)) cat_91 (
        .y(_T_441),
        .a(io_imem_bits_data),
        .b(_T_440)
    );
    wire [15:0] _T_442;
    SHR_UNSIGNED #(.width(64), .n(48)) u_shr_92 (
        .y(_T_442),
        .in(_T_441)
    );
    wire [31:0] _T_443;
    CAT #(.width_a(16), .width_b(16)) cat_93 (
        .y(_T_443),
        .a(_T_442),
        .b(_T_442)
    );
    wire [63:0] _T_444;
    CAT #(.width_a(32), .width_b(32)) cat_94 (
        .y(_T_444),
        .a(_T_443),
        .b(_T_443)
    );
    wire [127:0] _T_445;
    CAT #(.width_a(64), .width_b(64)) cat_95 (
        .y(_T_445),
        .a(_T_444),
        .b(_T_441)
    );
    wire [5:0] _T_446;
    SHL_UNSIGNED #(.width(2), .n(4)) u_shl_96 (
        .y(_T_446),
        .in(icShiftAmt)
    );
    wire [190:0] _T_447;
    DSHL_UNSIGNED #(.width_in(128), .width_n(6)) u_dshl_97 (
        .y(_T_447),
        .in(_T_445),
        .n(_T_446)
    );
    wire [31:0] icData;
    BITS #(.width(191), .high(95), .low(64)) bits_98 (
        .y(icData),
        .in(_T_447)
    );
    wire [31:0] _T_449;
    assign _T_449 = 32'hFFFFFFFF;
    wire [4:0] _T_450;
    SHL_UNSIGNED #(.width(1), .n(4)) u_shl_99 (
        .y(_T_450),
        .in(_nBufValid__q)
    );
    wire [62:0] _T_451;
    DSHL_UNSIGNED #(.width_in(32), .width_n(5)) u_dshl_100 (
        .y(_T_451),
        .in(_T_449),
        .n(_T_450)
    );
    wire [31:0] icMask;
    BITS #(.width(63), .high(31), .low(0)) bits_101 (
        .y(icMask),
        .in(_T_451)
    );
    wire [31:0] _T_452;
    BITWISEAND #(.width(32)) bitwiseand_102 (
        .y(_T_452),
        .a(icData),
        .b(icMask)
    );
    wire [31:0] _T_453;
    BITWISENOT #(.width(32)) bitwisenot_103 (
        .y(_T_453),
        .in(icMask)
    );
    wire [31:0] _T_454;
    BITWISEAND #(.width(32)) bitwiseand_104 (
        .y(_T_454),
        .a(_buf_data__q),
        .b(_T_453)
    );
    wire [31:0] inst;
    BITWISEOR #(.width(32)) bitwiseor_105 (
        .y(inst),
        .a(_T_452),
        .b(_T_454)
    );
    wire [3:0] _T_456;
    DSHL_UNSIGNED #(.width_in(1), .width_n(2)) u_dshl_106 (
        .y(_T_456),
        .in(1'h1),
        .n(nValid)
    );
    wire [4:0] _T_458;
    wire [3:0] _WTEMP_18;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_107 (
        .y(_WTEMP_18),
        .in(1'h1)
    );
    SUB_UNSIGNED #(.width(4)) u_sub_108 (
        .y(_T_458),
        .a(_T_456),
        .b(_WTEMP_18)
    );
    wire [4:0] _T_459;
    ASUINT #(.width(5)) asuint_109 (
        .y(_T_459),
        .in(_T_458)
    );
    wire [3:0] _T_460;
    TAIL #(.width(5), .n(1)) tail_110 (
        .y(_T_460),
        .in(_T_459)
    );
    wire [1:0] valid;
    BITS #(.width(4), .high(1), .low(0)) bits_111 (
        .y(valid),
        .in(_T_460)
    );
    wire [1:0] _T_462;
    DSHL_UNSIGNED #(.width_in(1), .width_n(1)) u_dshl_112 (
        .y(_T_462),
        .in(1'h1),
        .n(_nBufValid__q)
    );
    wire [2:0] _T_464;
    wire [1:0] _WTEMP_19;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_113 (
        .y(_WTEMP_19),
        .in(1'h1)
    );
    SUB_UNSIGNED #(.width(2)) u_sub_114 (
        .y(_T_464),
        .a(_T_462),
        .b(_WTEMP_19)
    );
    wire [2:0] _T_465;
    ASUINT #(.width(3)) asuint_115 (
        .y(_T_465),
        .in(_T_464)
    );
    wire [1:0] bufMask;
    TAIL #(.width(3), .n(1)) tail_116 (
        .y(bufMask),
        .in(_T_465)
    );
    wire [1:0] _T_467;
    wire [1:0] _WTEMP_20;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_117 (
        .y(_WTEMP_20),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_118 (
        .y(_T_467),
        .sel(_buf_xcpt_if__q),
        .a(bufMask),
        .b(_WTEMP_20)
    );
    wire [1:0] _T_468;
    BITWISENOT #(.width(2)) bitwisenot_119 (
        .y(_T_468),
        .in(bufMask)
    );
    wire [1:0] _T_470;
    wire [1:0] _WTEMP_21;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_120 (
        .y(_WTEMP_21),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_121 (
        .y(_T_470),
        .sel(io_imem_bits_xcpt_if),
        .a(_T_468),
        .b(_WTEMP_21)
    );
    wire [1:0] _T_471;
    BITWISEOR #(.width(2)) bitwiseor_122 (
        .y(_T_471),
        .a(_T_467),
        .b(_T_470)
    );
    wire [1:0] xcpt_if;
    BITWISEAND #(.width(2)) bitwiseand_123 (
        .y(xcpt_if),
        .a(valid),
        .b(_T_471)
    );
    wire [1:0] _T_473;
    wire [1:0] _WTEMP_22;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_124 (
        .y(_WTEMP_22),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_125 (
        .y(_T_473),
        .sel(_buf_replay__q),
        .a(bufMask),
        .b(_WTEMP_22)
    );
    wire [1:0] _T_474;
    BITWISENOT #(.width(2)) bitwisenot_126 (
        .y(_T_474),
        .in(bufMask)
    );
    wire [1:0] _T_476;
    wire [1:0] _WTEMP_23;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_127 (
        .y(_WTEMP_23),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_128 (
        .y(_T_476),
        .sel(io_imem_bits_replay),
        .a(_T_474),
        .b(_WTEMP_23)
    );
    wire [1:0] _T_477;
    BITWISEOR #(.width(2)) bitwiseor_129 (
        .y(_T_477),
        .a(_T_473),
        .b(_T_476)
    );
    wire [1:0] ic_replay;
    BITWISEAND #(.width(2)) bitwiseand_130 (
        .y(ic_replay),
        .a(valid),
        .b(_T_477)
    );
    wire [1:0] _T_479;
    DSHL_UNSIGNED #(.width_in(1), .width_n(1)) u_dshl_131 (
        .y(_T_479),
        .in(1'h1),
        .n(_ibufBTBResp_bridx__q)
    );
    wire [1:0] ibufBTBHitMask;
    wire [1:0] _WTEMP_24;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_132 (
        .y(_WTEMP_24),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_133 (
        .y(ibufBTBHitMask),
        .sel(_ibufBTBHit__q),
        .a(_T_479),
        .b(_WTEMP_24)
    );
    wire _T_482;
    EQ_UNSIGNED #(.width(1)) u_eq_134 (
        .y(_T_482),
        .a(io_imem_bits_btb_valid),
        .b(1'h0)
    );
    wire _T_483;
    GEQ_UNSIGNED #(.width(1)) u_geq_135 (
        .y(_T_483),
        .a(io_imem_bits_btb_bits_bridx),
        .b(pcWordBits)
    );
    wire _T_484;
    BITWISEOR #(.width(1)) bitwiseor_136 (
        .y(_T_484),
        .a(_T_482),
        .b(_T_483)
    );
    wire _T_485;
    BITWISEOR #(.width(1)) bitwiseor_137 (
        .y(_T_485),
        .a(_T_484),
        .b(reset)
    );
    wire _T_487;
    EQ_UNSIGNED #(.width(1)) u_eq_138 (
        .y(_T_487),
        .a(_T_485),
        .b(1'h0)
    );
    wire [1:0] _T_488;
    ADD_UNSIGNED #(.width(1)) u_add_139 (
        .y(_T_488),
        .a(io_imem_bits_btb_bits_bridx),
        .b(_nBufValid__q)
    );
    wire [2:0] _T_489;
    wire [1:0] _WTEMP_25;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_140 (
        .y(_WTEMP_25),
        .in(pcWordBits)
    );
    SUB_UNSIGNED #(.width(2)) u_sub_141 (
        .y(_T_489),
        .a(_T_488),
        .b(_WTEMP_25)
    );
    wire [2:0] _T_490;
    ASUINT #(.width(3)) asuint_142 (
        .y(_T_490),
        .in(_T_489)
    );
    wire [1:0] _T_491;
    TAIL #(.width(3), .n(1)) tail_143 (
        .y(_T_491),
        .in(_T_490)
    );
    wire [3:0] _T_493;
    DSHL_UNSIGNED #(.width_in(1), .width_n(2)) u_dshl_144 (
        .y(_T_493),
        .in(1'h1),
        .n(_T_491)
    );
    wire [3:0] icBTBHitMask;
    wire [3:0] _WTEMP_26;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_145 (
        .y(_WTEMP_26),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(4)) u_mux_146 (
        .y(icBTBHitMask),
        .sel(io_imem_bits_btb_valid),
        .a(_T_493),
        .b(_WTEMP_26)
    );
    wire [1:0] _T_495;
    BITWISEAND #(.width(2)) bitwiseand_147 (
        .y(_T_495),
        .a(ibufBTBHitMask),
        .b(bufMask)
    );
    wire [1:0] _T_496;
    BITWISENOT #(.width(2)) bitwisenot_148 (
        .y(_T_496),
        .in(bufMask)
    );
    wire [3:0] _T_497;
    wire [3:0] _WTEMP_27;
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_149 (
        .y(_WTEMP_27),
        .in(_T_496)
    );
    BITWISEAND #(.width(4)) bitwiseand_150 (
        .y(_T_497),
        .a(icBTBHitMask),
        .b(_WTEMP_27)
    );
    wire [3:0] btbHitMask;
    wire [3:0] _WTEMP_28;
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_151 (
        .y(_WTEMP_28),
        .in(_T_495)
    );
    BITWISEOR #(.width(4)) bitwiseor_152 (
        .y(btbHitMask),
        .a(_WTEMP_28),
        .b(_T_497)
    );
    wire [1:0] _T_498;
    BITWISEAND #(.width(2)) bitwiseand_153 (
        .y(_T_498),
        .a(ibufBTBHitMask),
        .b(bufMask)
    );
    wire _T_500;
    wire [1:0] _WTEMP_29;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_154 (
        .y(_WTEMP_29),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(2)) u_neq_155 (
        .y(_T_500),
        .a(_T_498),
        .b(_WTEMP_29)
    );
    wire _T_501_taken;
    MUX_UNSIGNED #(.width(1)) u_mux_156 (
        .y(_T_501_taken),
        .sel(_T_500),
        .a(_ibufBTBResp_taken__q),
        .b(io_imem_bits_btb_bits_taken)
    );
    wire [1:0] _T_501_mask;
    MUX_UNSIGNED #(.width(2)) u_mux_157 (
        .y(_T_501_mask),
        .sel(_T_500),
        .a(_ibufBTBResp_mask__q),
        .b(io_imem_bits_btb_bits_mask)
    );
    wire _T_501_bridx;
    MUX_UNSIGNED #(.width(1)) u_mux_158 (
        .y(_T_501_bridx),
        .sel(_T_500),
        .a(_ibufBTBResp_bridx__q),
        .b(io_imem_bits_btb_bits_bridx)
    );
    wire [38:0] _T_501_target;
    MUX_UNSIGNED #(.width(39)) u_mux_159 (
        .y(_T_501_target),
        .sel(_T_500),
        .a(_ibufBTBResp_target__q),
        .b(io_imem_bits_btb_bits_target)
    );
    wire [5:0] _T_501_entry;
    MUX_UNSIGNED #(.width(6)) u_mux_160 (
        .y(_T_501_entry),
        .sel(_T_500),
        .a(_ibufBTBResp_entry__q),
        .b(io_imem_bits_btb_bits_entry)
    );
    wire [6:0] _T_501_bht_history;
    MUX_UNSIGNED #(.width(7)) u_mux_161 (
        .y(_T_501_bht_history),
        .sel(_T_500),
        .a(_ibufBTBResp_bht_history__q),
        .b(io_imem_bits_btb_bits_bht_history)
    );
    wire [1:0] _T_501_bht_value;
    MUX_UNSIGNED #(.width(2)) u_mux_162 (
        .y(_T_501_bht_value),
        .sel(_T_500),
        .a(_ibufBTBResp_bht_value__q),
        .b(io_imem_bits_btb_bits_bht_value)
    );
    wire _T_511;
    GT_UNSIGNED #(.width(1)) u_gt_163 (
        .y(_T_511),
        .a(_nBufValid__q),
        .b(1'h0)
    );
    wire [39:0] _T_512;
    MUX_UNSIGNED #(.width(40)) u_mux_164 (
        .y(_T_512),
        .sel(_T_511),
        .a(_buf_pc__q),
        .b(io_imem_bits_pc)
    );
    wire _RVCExpander__clock;
    wire _RVCExpander__reset;
    wire [31:0] _RVCExpander__io_in;
    wire [31:0] _RVCExpander__io_out_bits;
    wire [4:0] _RVCExpander__io_out_rd;
    wire [4:0] _RVCExpander__io_out_rs1;
    wire [4:0] _RVCExpander__io_out_rs2;
    wire [4:0] _RVCExpander__io_out_rs3;
    wire _RVCExpander__io_rvc;
    RVCExpander RVCExpander (
        .clock(_RVCExpander__clock),
        .reset(_RVCExpander__reset),
        .io_in(_RVCExpander__io_in),
        .io_out_bits(_RVCExpander__io_out_bits),
        .io_out_rd(_RVCExpander__io_out_rd),
        .io_out_rs1(_RVCExpander__io_out_rs1),
        .io_out_rs2(_RVCExpander__io_out_rs2),
        .io_out_rs3(_RVCExpander__io_out_rs3),
        .io_rvc(_RVCExpander__io_rvc)
    );
    wire [1:0] _T_514;
    DSHR_UNSIGNED #(.width_in(2), .width_n(1)) u_dshr_1283 (
        .y(_T_514),
        .in(ic_replay),
        .n(1'h0)
    );
    wire _T_515;
    BITS #(.width(2), .high(0), .low(0)) bits_1284 (
        .y(_T_515),
        .in(_T_514)
    );
    wire _T_517;
    EQ_UNSIGNED #(.width(1)) u_eq_1285 (
        .y(_T_517),
        .a(_RVCExpander__io_rvc),
        .b(1'h0)
    );
    wire [3:0] _T_518;
    DSHR_UNSIGNED #(.width_in(4), .width_n(1)) u_dshr_1286 (
        .y(_T_518),
        .in(btbHitMask),
        .n(1'h0)
    );
    wire _T_519;
    BITS #(.width(4), .high(0), .low(0)) bits_1287 (
        .y(_T_519),
        .in(_T_518)
    );
    wire [1:0] _T_521;
    assign _T_521 = 2'h1;
    wire _T_522;
    assign _T_522 = 1'h1;
    wire [1:0] _T_523;
    DSHR_UNSIGNED #(.width_in(2), .width_n(1)) u_dshr_1288 (
        .y(_T_523),
        .in(ic_replay),
        .n(_T_522)
    );
    wire _T_524;
    BITS #(.width(2), .high(0), .low(0)) bits_1289 (
        .y(_T_524),
        .in(_T_523)
    );
    wire _T_525;
    BITWISEOR #(.width(1)) bitwiseor_1290 (
        .y(_T_525),
        .a(_T_519),
        .b(_T_524)
    );
    wire _T_526;
    BITWISEAND #(.width(1)) bitwiseand_1291 (
        .y(_T_526),
        .a(_T_517),
        .b(_T_525)
    );
    wire _T_527;
    BITWISEOR #(.width(1)) bitwiseor_1292 (
        .y(_T_527),
        .a(_T_515),
        .b(_T_526)
    );
    wire [1:0] _T_528;
    DSHR_UNSIGNED #(.width_in(2), .width_n(1)) u_dshr_1293 (
        .y(_T_528),
        .in(valid),
        .n(1'h0)
    );
    wire _T_529;
    BITS #(.width(2), .high(0), .low(0)) bits_1294 (
        .y(_T_529),
        .in(_T_528)
    );
    wire [1:0] _T_531;
    assign _T_531 = 2'h1;
    wire _T_532;
    assign _T_532 = 1'h1;
    wire [1:0] _T_533;
    DSHR_UNSIGNED #(.width_in(2), .width_n(1)) u_dshr_1295 (
        .y(_T_533),
        .in(valid),
        .n(_T_532)
    );
    wire _T_534;
    BITS #(.width(2), .high(0), .low(0)) bits_1296 (
        .y(_T_534),
        .in(_T_533)
    );
    wire _T_535;
    BITWISEOR #(.width(1)) bitwiseor_1297 (
        .y(_T_535),
        .a(_RVCExpander__io_rvc),
        .b(_T_534)
    );
    wire [1:0] _T_537;
    assign _T_537 = 2'h1;
    wire _T_538;
    assign _T_538 = 1'h1;
    wire [1:0] _T_539;
    DSHR_UNSIGNED #(.width_in(2), .width_n(1)) u_dshr_1298 (
        .y(_T_539),
        .in(xcpt_if),
        .n(_T_538)
    );
    wire _T_540;
    BITS #(.width(2), .high(0), .low(0)) bits_1299 (
        .y(_T_540),
        .in(_T_539)
    );
    wire _T_541;
    BITWISEOR #(.width(1)) bitwiseor_1300 (
        .y(_T_541),
        .a(_T_535),
        .b(_T_540)
    );
    wire _T_542;
    BITWISEOR #(.width(1)) bitwiseor_1301 (
        .y(_T_542),
        .a(_T_541),
        .b(_T_527)
    );
    wire _T_543;
    BITWISEAND #(.width(1)) bitwiseand_1302 (
        .y(_T_543),
        .a(_T_529),
        .b(_T_542)
    );
    wire [1:0] _T_544;
    DSHR_UNSIGNED #(.width_in(2), .width_n(1)) u_dshr_1303 (
        .y(_T_544),
        .in(xcpt_if),
        .n(1'h0)
    );
    wire _T_545;
    BITS #(.width(2), .high(0), .low(0)) bits_1304 (
        .y(_T_545),
        .in(_T_544)
    );
    wire _T_547;
    EQ_UNSIGNED #(.width(1)) u_eq_1305 (
        .y(_T_547),
        .a(_RVCExpander__io_rvc),
        .b(1'h0)
    );
    wire [1:0] _T_549;
    assign _T_549 = 2'h1;
    wire _T_550;
    assign _T_550 = 1'h1;
    wire [1:0] _T_551;
    DSHR_UNSIGNED #(.width_in(2), .width_n(1)) u_dshr_1306 (
        .y(_T_551),
        .in(xcpt_if),
        .n(_T_550)
    );
    wire _T_552;
    BITS #(.width(2), .high(0), .low(0)) bits_1307 (
        .y(_T_552),
        .in(_T_551)
    );
    wire _T_553;
    BITWISEAND #(.width(1)) bitwiseand_1308 (
        .y(_T_553),
        .a(_T_547),
        .b(_T_552)
    );
    wire [3:0] _T_554;
    DSHR_UNSIGNED #(.width_in(4), .width_n(1)) u_dshr_1309 (
        .y(_T_554),
        .in(btbHitMask),
        .n(1'h0)
    );
    wire _T_555;
    BITS #(.width(4), .high(0), .low(0)) bits_1310 (
        .y(_T_555),
        .in(_T_554)
    );
    wire _T_557;
    EQ_UNSIGNED #(.width(1)) u_eq_1311 (
        .y(_T_557),
        .a(_RVCExpander__io_rvc),
        .b(1'h0)
    );
    wire [1:0] _T_559;
    assign _T_559 = 2'h1;
    wire _T_560;
    assign _T_560 = 1'h1;
    wire [3:0] _T_561;
    DSHR_UNSIGNED #(.width_in(4), .width_n(1)) u_dshr_1312 (
        .y(_T_561),
        .in(btbHitMask),
        .n(_T_560)
    );
    wire _T_562;
    BITS #(.width(4), .high(0), .low(0)) bits_1313 (
        .y(_T_562),
        .in(_T_561)
    );
    wire _T_563;
    BITWISEAND #(.width(1)) bitwiseand_1314 (
        .y(_T_563),
        .a(_T_557),
        .b(_T_562)
    );
    wire _T_564;
    BITWISEOR #(.width(1)) bitwiseor_1315 (
        .y(_T_564),
        .a(_T_555),
        .b(_T_563)
    );
    wire _T_565;
    BITWISEAND #(.width(1)) bitwiseand_1316 (
        .y(_T_565),
        .a(io_inst_0_ready),
        .b(io_inst_0_valid)
    );
    wire [1:0] _T_567;
    assign _T_567 = 2'h1;
    wire _T_568;
    assign _T_568 = 1'h1;
    wire [2:0] _T_570;
    assign _T_570 = 3'h2;
    wire [1:0] _T_571;
    assign _T_571 = 2'h2;
    wire [1:0] _T_572;
    wire [1:0] _WTEMP_106;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_1317 (
        .y(_WTEMP_106),
        .in(_T_568)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_1318 (
        .y(_T_572),
        .sel(_RVCExpander__io_rvc),
        .a(_WTEMP_106),
        .b(_T_571)
    );
    wire [1:0] _T_574;
    assign _T_574 = 2'h1;
    wire _T_575;
    assign _T_575 = 1'h1;
    wire [2:0] _T_577;
    assign _T_577 = 3'h2;
    wire [1:0] _T_578;
    assign _T_578 = 2'h2;
    wire [1:0] _T_579;
    wire [1:0] _WTEMP_107;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_1319 (
        .y(_WTEMP_107),
        .in(_T_575)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_1320 (
        .y(_T_579),
        .sel(_RVCExpander__io_rvc),
        .a(_WTEMP_107),
        .b(_T_578)
    );
    wire [15:0] _T_580;
    SHR_UNSIGNED #(.width(32), .n(16)) u_shr_1321 (
        .y(_T_580),
        .in(inst)
    );
    wire _T_581;
    SHR_UNSIGNED #(.width(32), .n(32)) u_shr_1322 (
        .y(_T_581),
        .in(inst)
    );
    wire [15:0] _T_582;
    wire [15:0] _WTEMP_108;
    PAD_UNSIGNED #(.width(1), .n(16)) u_pad_1323 (
        .y(_WTEMP_108),
        .in(_T_581)
    );
    MUX_UNSIGNED #(.width(16)) u_mux_1324 (
        .y(_T_582),
        .sel(_RVCExpander__io_rvc),
        .a(_T_580),
        .b(_WTEMP_108)
    );
    assign _RVCExpander__clock = clock;
    assign _RVCExpander__io_in = inst;
    assign _RVCExpander__reset = reset;
    MUX_UNSIGNED #(.width(7)) u_mux_1325 (
        .y(_buf_btb_bits_bht_history__d),
        .sel(_T_411),
        .a(io_imem_bits_btb_bits_bht_history),
        .b(_buf_btb_bits_bht_history__q)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_1326 (
        .y(_buf_btb_bits_bht_value__d),
        .sel(_T_411),
        .a(io_imem_bits_btb_bits_bht_value),
        .b(_buf_btb_bits_bht_value__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_1327 (
        .y(_buf_btb_bits_bridx__d),
        .sel(_T_411),
        .a(io_imem_bits_btb_bits_bridx),
        .b(_buf_btb_bits_bridx__q)
    );
    MUX_UNSIGNED #(.width(6)) u_mux_1328 (
        .y(_buf_btb_bits_entry__d),
        .sel(_T_411),
        .a(io_imem_bits_btb_bits_entry),
        .b(_buf_btb_bits_entry__q)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_1329 (
        .y(_buf_btb_bits_mask__d),
        .sel(_T_411),
        .a(io_imem_bits_btb_bits_mask),
        .b(_buf_btb_bits_mask__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_1330 (
        .y(_buf_btb_bits_taken__d),
        .sel(_T_411),
        .a(io_imem_bits_btb_bits_taken),
        .b(_buf_btb_bits_taken__q)
    );
    MUX_UNSIGNED #(.width(39)) u_mux_1331 (
        .y(_buf_btb_bits_target__d),
        .sel(_T_411),
        .a(io_imem_bits_btb_bits_target),
        .b(_buf_btb_bits_target__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_1332 (
        .y(_buf_btb_valid__d),
        .sel(_T_411),
        .a(io_imem_bits_btb_valid),
        .b(_buf_btb_valid__q)
    );
    wire [31:0] _WTEMP_109;
    PAD_UNSIGNED #(.width(16), .n(32)) u_pad_1333 (
        .y(_WTEMP_109),
        .in(_T_422)
    );
    MUX_UNSIGNED #(.width(32)) u_mux_1334 (
        .y(_buf_data__d),
        .sel(_T_411),
        .a(_WTEMP_109),
        .b(_buf_data__q)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_1335 (
        .y(_buf_mask__d),
        .sel(_T_411),
        .a(io_imem_bits_mask),
        .b(_buf_mask__q)
    );
    MUX_UNSIGNED #(.width(40)) u_mux_1336 (
        .y(_buf_pc__d),
        .sel(_T_411),
        .a(_T_429),
        .b(_buf_pc__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_1337 (
        .y(_buf_replay__d),
        .sel(_T_411),
        .a(io_imem_bits_replay),
        .b(_buf_replay__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_1338 (
        .y(_buf_xcpt_if__d),
        .sel(_T_411),
        .a(io_imem_bits_xcpt_if),
        .b(_buf_xcpt_if__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_1339 (
        .y(_ibufBTBHit__d),
        .sel(_T_411),
        .a(io_imem_bits_btb_valid),
        .b(_ibufBTBHit__q)
    );
    MUX_UNSIGNED #(.width(7)) u_mux_1340 (
        .y(_ibufBTBResp_bht_history__d),
        .sel(_T_411),
        .a(_node_0),
        .b(_ibufBTBResp_bht_history__q)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_1341 (
        .y(_ibufBTBResp_bht_value__d),
        .sel(_T_411),
        .a(_node_1),
        .b(_ibufBTBResp_bht_value__q)
    );
    wire [1:0] _WTEMP_110;
    BITS #(.width(2), .high(0), .low(0)) bits_1342 (
        .y(_ibufBTBResp_bridx__d),
        .in(_WTEMP_110)
    );
    wire [1:0] _WTEMP_111;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_1343 (
        .y(_WTEMP_111),
        .in(_ibufBTBResp_bridx__q)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_1344 (
        .y(_WTEMP_110),
        .sel(_T_411),
        .a(_node_2),
        .b(_WTEMP_111)
    );
    MUX_UNSIGNED #(.width(6)) u_mux_1345 (
        .y(_ibufBTBResp_entry__d),
        .sel(_T_411),
        .a(_node_3),
        .b(_ibufBTBResp_entry__q)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_1346 (
        .y(_ibufBTBResp_mask__d),
        .sel(_T_411),
        .a(_node_4),
        .b(_ibufBTBResp_mask__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_1347 (
        .y(_ibufBTBResp_taken__d),
        .sel(_T_411),
        .a(_node_5),
        .b(_ibufBTBResp_taken__q)
    );
    MUX_UNSIGNED #(.width(39)) u_mux_1348 (
        .y(_ibufBTBResp_target__d),
        .sel(_T_411),
        .a(_node_6),
        .b(_ibufBTBResp_target__q)
    );
    assign io_btb_resp_bht_history = _T_501_bht_history;
    assign io_btb_resp_bht_value = _T_501_bht_value;
    assign io_btb_resp_bridx = _T_501_bridx;
    assign io_btb_resp_entry = _T_501_entry;
    assign io_btb_resp_mask = _T_501_mask;
    assign io_btb_resp_taken = _T_501_taken;
    assign io_btb_resp_target = _T_501_target;
    assign io_imem_ready = _T_395;
    assign io_inst_0_bits_btb_hit = _T_564;
    assign io_inst_0_bits_inst_bits = _RVCExpander__io_out_bits;
    assign io_inst_0_bits_inst_rd = _RVCExpander__io_out_rd;
    assign io_inst_0_bits_inst_rs1 = _RVCExpander__io_out_rs1;
    assign io_inst_0_bits_inst_rs2 = _RVCExpander__io_out_rs2;
    assign io_inst_0_bits_inst_rs3 = _RVCExpander__io_out_rs3;
    assign io_inst_0_bits_pf0 = _T_545;
    assign io_inst_0_bits_pf1 = _T_553;
    assign io_inst_0_bits_raw = inst;
    assign io_inst_0_bits_replay = _T_527;
    assign io_inst_0_bits_rvc = _RVCExpander__io_rvc;
    assign io_inst_0_valid = _T_543;
    assign io_pc = _T_512;
    wire [1:0] _WTEMP_112;
    wire [1:0] _WTEMP_113;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_1349 (
        .y(_WTEMP_113),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_1350 (
        .y(_WTEMP_112),
        .sel(io_kill),
        .a(_WTEMP_113),
        .b(_node_7)
    );
    BITS #(.width(2), .high(0), .low(0)) bits_1351 (
        .y(_WTEMP_0),
        .in(_WTEMP_112)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_1352 (
        .y(nReady),
        .sel(_T_565),
        .a(_T_572),
        .b(2'h0)
    );
endmodule //IBuf
module MUX_UNSIGNED(y, sel, a, b);
    parameter width = 4;
    output [width-1:0] y;
    input sel;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = sel ? a : b;
endmodule // MUX_UNSIGNED
module BITS(y, in);
    parameter width = 4;
    parameter high = 2;
    parameter low = 0;
    output [high-low:0] y;
    input [width-1:0] in;
    assign y = in[high:low];
endmodule // BITS
module BITWISEAND(y, a, b);
    parameter width = 4;
    output [width-1:0] y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a & b;
endmodule // BITWISEAND
module ADD_UNSIGNED(y, a, b);
    parameter width = 4;
    output [width:0] y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a + b;
endmodule // ADD_UNSIGNED
module PAD_UNSIGNED(y, in);
    parameter width = 4;
    parameter n = 4;
    output [(n > width ? n : width)-1:0] y;
    input [width-1:0] in;
    assign y = (n > width) ? {{(n - width){1'b0}}, in} : in;
endmodule // PAD_UNSIGNED
module SUB_UNSIGNED(y, a, b);
    parameter width = 4;
    output [width:0] y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a - b;
endmodule // SUB_UNSIGNED
module ASUINT(y, in);
    parameter width = 4;
    output [width-1:0] y;
    input [width-1:0] in;
    assign y = $unsigned(in);
endmodule // ASUINT
module TAIL(y, in);
    parameter width = 4;
    parameter n = 2;
    output [width-n-1:0] y;
    input [width-1:0] in;
    assign y = in[width-n-1:0];
endmodule // TAIL
module GEQ_UNSIGNED(y, a, b);
    parameter width = 4;
    output y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a >= b;
endmodule // GEQ_UNSIGNED
module LT_UNSIGNED(y, a, b);
    parameter width = 4;
    output y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a < b;
endmodule // LT_UNSIGNED
module SHR_UNSIGNED(y, in);
    parameter width = 4;
    parameter n = 2;
    output [(n < width ? (width-n-1) : 0):0] y;
    input [width-1:0] in;
    assign y = n < width ? in[width-1:n] : 1'b0;
endmodule // SHR_UNSIGNED
module CAT(y, a, b);
    parameter width_a = 4;
    parameter width_b = 4;
    output [width_a+width_b-1:0] y;
    input [width_a-1:0] a;
    input [width_b-1:0] b;
    assign y = {a, b};
endmodule // CAT
module SHL_UNSIGNED(y, in);
    parameter width = 4;
    parameter n = 4;
    output [width+n-1:0] y;
    input [width-1:0] in;
    wire [width+n-1:0] temp;
    assign temp = {{n{1'b0}}, in};
    assign y = temp << n;
endmodule // SHL_UNSIGNED
module DSHR_UNSIGNED(y, in, n);
    parameter width_in = 4;
    parameter width_n = 2;
    output [width_in-1:0] y;
    input [width_in-1:0] in;
    input [width_n-1:0] n;
    assign y = in >> n;
endmodule // DSHR_UNSIGNED
module DSHL_UNSIGNED(y, in, n);
    parameter width_in = 4;
    parameter width_n = 2;
    output [(width_in+2**width_n-1)-1:0] y;
    input [width_in-1:0] in;
    input [width_n-1:0] n;
    wire [(width_in+2**width_n-1)-1:0] temp;
    assign temp = {{(2**width_n-1){1'b0}}, in};
    assign y = temp << n;
endmodule // DSHL_UNSIGNED
module BITWISENOT(y, in);
    parameter width = 4;
    output [width-1:0] y;
    input [width-1:0] in;
    assign y = ~in;
endmodule // BITWISENOT
module EQ_UNSIGNED(y, a, b);
    parameter width = 4;
    output y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a == b;
endmodule // EQ_UNSIGNED
module NEQ_UNSIGNED(y, a, b);
    parameter width = 4;
    output y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a != b;
endmodule // NEQ_UNSIGNED
module GT_UNSIGNED(y, a, b);
    parameter width = 4;
    output y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a > b;
endmodule // GT_UNSIGNED
module RVCExpander(
    input clock,
    input reset,
    input [31:0] io_in,
    output [31:0] io_out_bits,
    output [4:0] io_out_rd,
    output [4:0] io_out_rs1,
    output [4:0] io_out_rs2,
    output [4:0] io_out_rs3,
    output io_rvc
);
    wire [1:0] _T_12;
    BITS #(.width(32), .high(1), .low(0)) bits_165 (
        .y(_T_12),
        .in(io_in)
    );
    wire _T_14;
    NEQ_UNSIGNED #(.width(2)) u_neq_166 (
        .y(_T_14),
        .a(_T_12),
        .b(2'h3)
    );
    wire [7:0] _T_15;
    BITS #(.width(32), .high(12), .low(5)) bits_167 (
        .y(_T_15),
        .in(io_in)
    );
    wire _T_17;
    wire [7:0] _WTEMP_30;
    PAD_UNSIGNED #(.width(1), .n(8)) u_pad_168 (
        .y(_WTEMP_30),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(8)) u_neq_169 (
        .y(_T_17),
        .a(_T_15),
        .b(_WTEMP_30)
    );
    wire [6:0] _T_20;
    MUX_UNSIGNED #(.width(7)) u_mux_170 (
        .y(_T_20),
        .sel(_T_17),
        .a(7'h13),
        .b(7'h1F)
    );
    wire [3:0] _T_21;
    BITS #(.width(32), .high(10), .low(7)) bits_171 (
        .y(_T_21),
        .in(io_in)
    );
    wire [1:0] _T_22;
    BITS #(.width(32), .high(12), .low(11)) bits_172 (
        .y(_T_22),
        .in(io_in)
    );
    wire _T_23;
    BITS #(.width(32), .high(5), .low(5)) bits_173 (
        .y(_T_23),
        .in(io_in)
    );
    wire _T_24;
    BITS #(.width(32), .high(6), .low(6)) bits_174 (
        .y(_T_24),
        .in(io_in)
    );
    wire [2:0] _T_26;
    CAT #(.width_a(1), .width_b(2)) cat_175 (
        .y(_T_26),
        .a(_T_24),
        .b(2'h0)
    );
    wire [5:0] _T_27;
    CAT #(.width_a(4), .width_b(2)) cat_176 (
        .y(_T_27),
        .a(_T_21),
        .b(_T_22)
    );
    wire [6:0] _T_28;
    CAT #(.width_a(6), .width_b(1)) cat_177 (
        .y(_T_28),
        .a(_T_27),
        .b(_T_23)
    );
    wire [9:0] _T_29;
    CAT #(.width_a(7), .width_b(3)) cat_178 (
        .y(_T_29),
        .a(_T_28),
        .b(_T_26)
    );
    wire [2:0] _T_33;
    BITS #(.width(32), .high(4), .low(2)) bits_179 (
        .y(_T_33),
        .in(io_in)
    );
    wire [4:0] _T_34;
    CAT #(.width_a(2), .width_b(3)) cat_180 (
        .y(_T_34),
        .a(2'h1),
        .b(_T_33)
    );
    wire [11:0] _T_35;
    CAT #(.width_a(5), .width_b(7)) cat_181 (
        .y(_T_35),
        .a(_T_34),
        .b(_T_20)
    );
    wire [14:0] _T_36;
    CAT #(.width_a(10), .width_b(5)) cat_182 (
        .y(_T_36),
        .a(_T_29),
        .b(5'h2)
    );
    wire [17:0] _T_37;
    CAT #(.width_a(15), .width_b(3)) cat_183 (
        .y(_T_37),
        .a(_T_36),
        .b(3'h0)
    );
    wire [29:0] _T_38;
    CAT #(.width_a(18), .width_b(12)) cat_184 (
        .y(_T_38),
        .a(_T_37),
        .b(_T_35)
    );
    wire [2:0] _T_40;
    BITS #(.width(32), .high(4), .low(2)) bits_185 (
        .y(_T_40),
        .in(io_in)
    );
    wire [4:0] _T_41;
    CAT #(.width_a(2), .width_b(3)) cat_186 (
        .y(_T_41),
        .a(2'h1),
        .b(_T_40)
    );
    wire [2:0] _T_44;
    BITS #(.width(32), .high(4), .low(2)) bits_187 (
        .y(_T_44),
        .in(io_in)
    );
    wire [4:0] _T_45;
    CAT #(.width_a(2), .width_b(3)) cat_188 (
        .y(_T_45),
        .a(2'h1),
        .b(_T_44)
    );
    wire [4:0] _T_46;
    BITS #(.width(32), .high(31), .low(27)) bits_189 (
        .y(_T_46),
        .in(io_in)
    );
    wire [31:0] _T_53_bits;
    wire [4:0] _T_53_rd;
    wire [4:0] _T_53_rs1;
    wire [4:0] _T_53_rs2;
    wire [4:0] _T_53_rs3;
    wire [1:0] _T_59;
    BITS #(.width(32), .high(6), .low(5)) bits_190 (
        .y(_T_59),
        .in(io_in)
    );
    wire [2:0] _T_60;
    BITS #(.width(32), .high(12), .low(10)) bits_191 (
        .y(_T_60),
        .in(io_in)
    );
    wire [4:0] _T_62;
    CAT #(.width_a(2), .width_b(3)) cat_192 (
        .y(_T_62),
        .a(_T_59),
        .b(_T_60)
    );
    wire [7:0] _T_63;
    CAT #(.width_a(5), .width_b(3)) cat_193 (
        .y(_T_63),
        .a(_T_62),
        .b(3'h0)
    );
    wire [2:0] _T_65;
    BITS #(.width(32), .high(9), .low(7)) bits_194 (
        .y(_T_65),
        .in(io_in)
    );
    wire [4:0] _T_66;
    CAT #(.width_a(2), .width_b(3)) cat_195 (
        .y(_T_66),
        .a(2'h1),
        .b(_T_65)
    );
    wire [2:0] _T_69;
    BITS #(.width(32), .high(4), .low(2)) bits_196 (
        .y(_T_69),
        .in(io_in)
    );
    wire [4:0] _T_70;
    CAT #(.width_a(2), .width_b(3)) cat_197 (
        .y(_T_70),
        .a(2'h1),
        .b(_T_69)
    );
    wire [11:0] _T_72;
    CAT #(.width_a(5), .width_b(7)) cat_198 (
        .y(_T_72),
        .a(_T_70),
        .b(7'h7)
    );
    wire [12:0] _T_73;
    CAT #(.width_a(8), .width_b(5)) cat_199 (
        .y(_T_73),
        .a(_T_63),
        .b(_T_66)
    );
    wire [15:0] _T_74;
    CAT #(.width_a(13), .width_b(3)) cat_200 (
        .y(_T_74),
        .a(_T_73),
        .b(3'h3)
    );
    wire [27:0] _T_75;
    CAT #(.width_a(16), .width_b(12)) cat_201 (
        .y(_T_75),
        .a(_T_74),
        .b(_T_72)
    );
    wire [2:0] _T_77;
    BITS #(.width(32), .high(4), .low(2)) bits_202 (
        .y(_T_77),
        .in(io_in)
    );
    wire [4:0] _T_78;
    CAT #(.width_a(2), .width_b(3)) cat_203 (
        .y(_T_78),
        .a(2'h1),
        .b(_T_77)
    );
    wire [2:0] _T_80;
    BITS #(.width(32), .high(9), .low(7)) bits_204 (
        .y(_T_80),
        .in(io_in)
    );
    wire [4:0] _T_81;
    CAT #(.width_a(2), .width_b(3)) cat_205 (
        .y(_T_81),
        .a(2'h1),
        .b(_T_80)
    );
    wire [2:0] _T_83;
    BITS #(.width(32), .high(4), .low(2)) bits_206 (
        .y(_T_83),
        .in(io_in)
    );
    wire [4:0] _T_84;
    CAT #(.width_a(2), .width_b(3)) cat_207 (
        .y(_T_84),
        .a(2'h1),
        .b(_T_83)
    );
    wire [4:0] _T_85;
    BITS #(.width(32), .high(31), .low(27)) bits_208 (
        .y(_T_85),
        .in(io_in)
    );
    wire [31:0] _T_92_bits;
    wire [4:0] _T_92_rd;
    wire [4:0] _T_92_rs1;
    wire [4:0] _T_92_rs2;
    wire [4:0] _T_92_rs3;
    wire _T_98;
    BITS #(.width(32), .high(5), .low(5)) bits_209 (
        .y(_T_98),
        .in(io_in)
    );
    wire [2:0] _T_99;
    BITS #(.width(32), .high(12), .low(10)) bits_210 (
        .y(_T_99),
        .in(io_in)
    );
    wire _T_100;
    BITS #(.width(32), .high(6), .low(6)) bits_211 (
        .y(_T_100),
        .in(io_in)
    );
    wire [2:0] _T_102;
    CAT #(.width_a(1), .width_b(2)) cat_212 (
        .y(_T_102),
        .a(_T_100),
        .b(2'h0)
    );
    wire [3:0] _T_103;
    CAT #(.width_a(1), .width_b(3)) cat_213 (
        .y(_T_103),
        .a(_T_98),
        .b(_T_99)
    );
    wire [6:0] _T_104;
    CAT #(.width_a(4), .width_b(3)) cat_214 (
        .y(_T_104),
        .a(_T_103),
        .b(_T_102)
    );
    wire [2:0] _T_106;
    BITS #(.width(32), .high(9), .low(7)) bits_215 (
        .y(_T_106),
        .in(io_in)
    );
    wire [4:0] _T_107;
    CAT #(.width_a(2), .width_b(3)) cat_216 (
        .y(_T_107),
        .a(2'h1),
        .b(_T_106)
    );
    wire [2:0] _T_110;
    BITS #(.width(32), .high(4), .low(2)) bits_217 (
        .y(_T_110),
        .in(io_in)
    );
    wire [4:0] _T_111;
    CAT #(.width_a(2), .width_b(3)) cat_218 (
        .y(_T_111),
        .a(2'h1),
        .b(_T_110)
    );
    wire [11:0] _T_113;
    CAT #(.width_a(5), .width_b(7)) cat_219 (
        .y(_T_113),
        .a(_T_111),
        .b(7'h3)
    );
    wire [11:0] _T_114;
    CAT #(.width_a(7), .width_b(5)) cat_220 (
        .y(_T_114),
        .a(_T_104),
        .b(_T_107)
    );
    wire [14:0] _T_115;
    CAT #(.width_a(12), .width_b(3)) cat_221 (
        .y(_T_115),
        .a(_T_114),
        .b(3'h2)
    );
    wire [26:0] _T_116;
    CAT #(.width_a(15), .width_b(12)) cat_222 (
        .y(_T_116),
        .a(_T_115),
        .b(_T_113)
    );
    wire [2:0] _T_118;
    BITS #(.width(32), .high(4), .low(2)) bits_223 (
        .y(_T_118),
        .in(io_in)
    );
    wire [4:0] _T_119;
    CAT #(.width_a(2), .width_b(3)) cat_224 (
        .y(_T_119),
        .a(2'h1),
        .b(_T_118)
    );
    wire [2:0] _T_121;
    BITS #(.width(32), .high(9), .low(7)) bits_225 (
        .y(_T_121),
        .in(io_in)
    );
    wire [4:0] _T_122;
    CAT #(.width_a(2), .width_b(3)) cat_226 (
        .y(_T_122),
        .a(2'h1),
        .b(_T_121)
    );
    wire [2:0] _T_124;
    BITS #(.width(32), .high(4), .low(2)) bits_227 (
        .y(_T_124),
        .in(io_in)
    );
    wire [4:0] _T_125;
    CAT #(.width_a(2), .width_b(3)) cat_228 (
        .y(_T_125),
        .a(2'h1),
        .b(_T_124)
    );
    wire [4:0] _T_126;
    BITS #(.width(32), .high(31), .low(27)) bits_229 (
        .y(_T_126),
        .in(io_in)
    );
    wire [31:0] _T_133_bits;
    wire [4:0] _T_133_rd;
    wire [4:0] _T_133_rs1;
    wire [4:0] _T_133_rs2;
    wire [4:0] _T_133_rs3;
    wire [1:0] _T_139;
    BITS #(.width(32), .high(6), .low(5)) bits_230 (
        .y(_T_139),
        .in(io_in)
    );
    wire [2:0] _T_140;
    BITS #(.width(32), .high(12), .low(10)) bits_231 (
        .y(_T_140),
        .in(io_in)
    );
    wire [4:0] _T_142;
    CAT #(.width_a(2), .width_b(3)) cat_232 (
        .y(_T_142),
        .a(_T_139),
        .b(_T_140)
    );
    wire [7:0] _T_143;
    CAT #(.width_a(5), .width_b(3)) cat_233 (
        .y(_T_143),
        .a(_T_142),
        .b(3'h0)
    );
    wire [2:0] _T_145;
    BITS #(.width(32), .high(9), .low(7)) bits_234 (
        .y(_T_145),
        .in(io_in)
    );
    wire [4:0] _T_146;
    CAT #(.width_a(2), .width_b(3)) cat_235 (
        .y(_T_146),
        .a(2'h1),
        .b(_T_145)
    );
    wire [2:0] _T_149;
    BITS #(.width(32), .high(4), .low(2)) bits_236 (
        .y(_T_149),
        .in(io_in)
    );
    wire [4:0] _T_150;
    CAT #(.width_a(2), .width_b(3)) cat_237 (
        .y(_T_150),
        .a(2'h1),
        .b(_T_149)
    );
    wire [11:0] _T_152;
    CAT #(.width_a(5), .width_b(7)) cat_238 (
        .y(_T_152),
        .a(_T_150),
        .b(7'h3)
    );
    wire [12:0] _T_153;
    CAT #(.width_a(8), .width_b(5)) cat_239 (
        .y(_T_153),
        .a(_T_143),
        .b(_T_146)
    );
    wire [15:0] _T_154;
    CAT #(.width_a(13), .width_b(3)) cat_240 (
        .y(_T_154),
        .a(_T_153),
        .b(3'h3)
    );
    wire [27:0] _T_155;
    CAT #(.width_a(16), .width_b(12)) cat_241 (
        .y(_T_155),
        .a(_T_154),
        .b(_T_152)
    );
    wire [2:0] _T_157;
    BITS #(.width(32), .high(4), .low(2)) bits_242 (
        .y(_T_157),
        .in(io_in)
    );
    wire [4:0] _T_158;
    CAT #(.width_a(2), .width_b(3)) cat_243 (
        .y(_T_158),
        .a(2'h1),
        .b(_T_157)
    );
    wire [2:0] _T_160;
    BITS #(.width(32), .high(9), .low(7)) bits_244 (
        .y(_T_160),
        .in(io_in)
    );
    wire [4:0] _T_161;
    CAT #(.width_a(2), .width_b(3)) cat_245 (
        .y(_T_161),
        .a(2'h1),
        .b(_T_160)
    );
    wire [2:0] _T_163;
    BITS #(.width(32), .high(4), .low(2)) bits_246 (
        .y(_T_163),
        .in(io_in)
    );
    wire [4:0] _T_164;
    CAT #(.width_a(2), .width_b(3)) cat_247 (
        .y(_T_164),
        .a(2'h1),
        .b(_T_163)
    );
    wire [4:0] _T_165;
    BITS #(.width(32), .high(31), .low(27)) bits_248 (
        .y(_T_165),
        .in(io_in)
    );
    wire [31:0] _T_172_bits;
    wire [4:0] _T_172_rd;
    wire [4:0] _T_172_rs1;
    wire [4:0] _T_172_rs2;
    wire [4:0] _T_172_rs3;
    wire _T_178;
    BITS #(.width(32), .high(5), .low(5)) bits_249 (
        .y(_T_178),
        .in(io_in)
    );
    wire [2:0] _T_179;
    BITS #(.width(32), .high(12), .low(10)) bits_250 (
        .y(_T_179),
        .in(io_in)
    );
    wire _T_180;
    BITS #(.width(32), .high(6), .low(6)) bits_251 (
        .y(_T_180),
        .in(io_in)
    );
    wire [2:0] _T_182;
    CAT #(.width_a(1), .width_b(2)) cat_252 (
        .y(_T_182),
        .a(_T_180),
        .b(2'h0)
    );
    wire [3:0] _T_183;
    CAT #(.width_a(1), .width_b(3)) cat_253 (
        .y(_T_183),
        .a(_T_178),
        .b(_T_179)
    );
    wire [6:0] _T_184;
    CAT #(.width_a(4), .width_b(3)) cat_254 (
        .y(_T_184),
        .a(_T_183),
        .b(_T_182)
    );
    wire [1:0] _T_185;
    SHR_UNSIGNED #(.width(7), .n(5)) u_shr_255 (
        .y(_T_185),
        .in(_T_184)
    );
    wire [2:0] _T_187;
    BITS #(.width(32), .high(4), .low(2)) bits_256 (
        .y(_T_187),
        .in(io_in)
    );
    wire [4:0] _T_188;
    CAT #(.width_a(2), .width_b(3)) cat_257 (
        .y(_T_188),
        .a(2'h1),
        .b(_T_187)
    );
    wire [2:0] _T_190;
    BITS #(.width(32), .high(9), .low(7)) bits_258 (
        .y(_T_190),
        .in(io_in)
    );
    wire [4:0] _T_191;
    CAT #(.width_a(2), .width_b(3)) cat_259 (
        .y(_T_191),
        .a(2'h1),
        .b(_T_190)
    );
    wire _T_193;
    BITS #(.width(32), .high(5), .low(5)) bits_260 (
        .y(_T_193),
        .in(io_in)
    );
    wire [2:0] _T_194;
    BITS #(.width(32), .high(12), .low(10)) bits_261 (
        .y(_T_194),
        .in(io_in)
    );
    wire _T_195;
    BITS #(.width(32), .high(6), .low(6)) bits_262 (
        .y(_T_195),
        .in(io_in)
    );
    wire [2:0] _T_197;
    CAT #(.width_a(1), .width_b(2)) cat_263 (
        .y(_T_197),
        .a(_T_195),
        .b(2'h0)
    );
    wire [3:0] _T_198;
    CAT #(.width_a(1), .width_b(3)) cat_264 (
        .y(_T_198),
        .a(_T_193),
        .b(_T_194)
    );
    wire [6:0] _T_199;
    CAT #(.width_a(4), .width_b(3)) cat_265 (
        .y(_T_199),
        .a(_T_198),
        .b(_T_197)
    );
    wire [4:0] _T_200;
    BITS #(.width(7), .high(4), .low(0)) bits_266 (
        .y(_T_200),
        .in(_T_199)
    );
    wire [7:0] _T_202;
    CAT #(.width_a(3), .width_b(5)) cat_267 (
        .y(_T_202),
        .a(3'h2),
        .b(_T_200)
    );
    wire [14:0] _T_203;
    CAT #(.width_a(8), .width_b(7)) cat_268 (
        .y(_T_203),
        .a(_T_202),
        .b(7'h2F)
    );
    wire [6:0] _T_204;
    CAT #(.width_a(2), .width_b(5)) cat_269 (
        .y(_T_204),
        .a(_T_185),
        .b(_T_188)
    );
    wire [11:0] _T_205;
    CAT #(.width_a(7), .width_b(5)) cat_270 (
        .y(_T_205),
        .a(_T_204),
        .b(_T_191)
    );
    wire [26:0] _T_206;
    CAT #(.width_a(12), .width_b(15)) cat_271 (
        .y(_T_206),
        .a(_T_205),
        .b(_T_203)
    );
    wire [2:0] _T_208;
    BITS #(.width(32), .high(4), .low(2)) bits_272 (
        .y(_T_208),
        .in(io_in)
    );
    wire [4:0] _T_209;
    CAT #(.width_a(2), .width_b(3)) cat_273 (
        .y(_T_209),
        .a(2'h1),
        .b(_T_208)
    );
    wire [2:0] _T_211;
    BITS #(.width(32), .high(9), .low(7)) bits_274 (
        .y(_T_211),
        .in(io_in)
    );
    wire [4:0] _T_212;
    CAT #(.width_a(2), .width_b(3)) cat_275 (
        .y(_T_212),
        .a(2'h1),
        .b(_T_211)
    );
    wire [2:0] _T_214;
    BITS #(.width(32), .high(4), .low(2)) bits_276 (
        .y(_T_214),
        .in(io_in)
    );
    wire [4:0] _T_215;
    CAT #(.width_a(2), .width_b(3)) cat_277 (
        .y(_T_215),
        .a(2'h1),
        .b(_T_214)
    );
    wire [4:0] _T_216;
    BITS #(.width(32), .high(31), .low(27)) bits_278 (
        .y(_T_216),
        .in(io_in)
    );
    wire [31:0] _T_223_bits;
    wire [4:0] _T_223_rd;
    wire [4:0] _T_223_rs1;
    wire [4:0] _T_223_rs2;
    wire [4:0] _T_223_rs3;
    wire [1:0] _T_229;
    BITS #(.width(32), .high(6), .low(5)) bits_279 (
        .y(_T_229),
        .in(io_in)
    );
    wire [2:0] _T_230;
    BITS #(.width(32), .high(12), .low(10)) bits_280 (
        .y(_T_230),
        .in(io_in)
    );
    wire [4:0] _T_232;
    CAT #(.width_a(2), .width_b(3)) cat_281 (
        .y(_T_232),
        .a(_T_229),
        .b(_T_230)
    );
    wire [7:0] _T_233;
    CAT #(.width_a(5), .width_b(3)) cat_282 (
        .y(_T_233),
        .a(_T_232),
        .b(3'h0)
    );
    wire [2:0] _T_234;
    SHR_UNSIGNED #(.width(8), .n(5)) u_shr_283 (
        .y(_T_234),
        .in(_T_233)
    );
    wire [2:0] _T_236;
    BITS #(.width(32), .high(4), .low(2)) bits_284 (
        .y(_T_236),
        .in(io_in)
    );
    wire [4:0] _T_237;
    CAT #(.width_a(2), .width_b(3)) cat_285 (
        .y(_T_237),
        .a(2'h1),
        .b(_T_236)
    );
    wire [2:0] _T_239;
    BITS #(.width(32), .high(9), .low(7)) bits_286 (
        .y(_T_239),
        .in(io_in)
    );
    wire [4:0] _T_240;
    CAT #(.width_a(2), .width_b(3)) cat_287 (
        .y(_T_240),
        .a(2'h1),
        .b(_T_239)
    );
    wire [1:0] _T_242;
    BITS #(.width(32), .high(6), .low(5)) bits_288 (
        .y(_T_242),
        .in(io_in)
    );
    wire [2:0] _T_243;
    BITS #(.width(32), .high(12), .low(10)) bits_289 (
        .y(_T_243),
        .in(io_in)
    );
    wire [4:0] _T_245;
    CAT #(.width_a(2), .width_b(3)) cat_290 (
        .y(_T_245),
        .a(_T_242),
        .b(_T_243)
    );
    wire [7:0] _T_246;
    CAT #(.width_a(5), .width_b(3)) cat_291 (
        .y(_T_246),
        .a(_T_245),
        .b(3'h0)
    );
    wire [4:0] _T_247;
    BITS #(.width(8), .high(4), .low(0)) bits_292 (
        .y(_T_247),
        .in(_T_246)
    );
    wire [7:0] _T_249;
    CAT #(.width_a(3), .width_b(5)) cat_293 (
        .y(_T_249),
        .a(3'h3),
        .b(_T_247)
    );
    wire [14:0] _T_250;
    CAT #(.width_a(8), .width_b(7)) cat_294 (
        .y(_T_250),
        .a(_T_249),
        .b(7'h27)
    );
    wire [7:0] _T_251;
    CAT #(.width_a(3), .width_b(5)) cat_295 (
        .y(_T_251),
        .a(_T_234),
        .b(_T_237)
    );
    wire [12:0] _T_252;
    CAT #(.width_a(8), .width_b(5)) cat_296 (
        .y(_T_252),
        .a(_T_251),
        .b(_T_240)
    );
    wire [27:0] _T_253;
    CAT #(.width_a(13), .width_b(15)) cat_297 (
        .y(_T_253),
        .a(_T_252),
        .b(_T_250)
    );
    wire [2:0] _T_255;
    BITS #(.width(32), .high(4), .low(2)) bits_298 (
        .y(_T_255),
        .in(io_in)
    );
    wire [4:0] _T_256;
    CAT #(.width_a(2), .width_b(3)) cat_299 (
        .y(_T_256),
        .a(2'h1),
        .b(_T_255)
    );
    wire [2:0] _T_258;
    BITS #(.width(32), .high(9), .low(7)) bits_300 (
        .y(_T_258),
        .in(io_in)
    );
    wire [4:0] _T_259;
    CAT #(.width_a(2), .width_b(3)) cat_301 (
        .y(_T_259),
        .a(2'h1),
        .b(_T_258)
    );
    wire [2:0] _T_261;
    BITS #(.width(32), .high(4), .low(2)) bits_302 (
        .y(_T_261),
        .in(io_in)
    );
    wire [4:0] _T_262;
    CAT #(.width_a(2), .width_b(3)) cat_303 (
        .y(_T_262),
        .a(2'h1),
        .b(_T_261)
    );
    wire [4:0] _T_263;
    BITS #(.width(32), .high(31), .low(27)) bits_304 (
        .y(_T_263),
        .in(io_in)
    );
    wire [31:0] _T_270_bits;
    wire [4:0] _T_270_rd;
    wire [4:0] _T_270_rs1;
    wire [4:0] _T_270_rs2;
    wire [4:0] _T_270_rs3;
    wire _T_276;
    BITS #(.width(32), .high(5), .low(5)) bits_305 (
        .y(_T_276),
        .in(io_in)
    );
    wire [2:0] _T_277;
    BITS #(.width(32), .high(12), .low(10)) bits_306 (
        .y(_T_277),
        .in(io_in)
    );
    wire _T_278;
    BITS #(.width(32), .high(6), .low(6)) bits_307 (
        .y(_T_278),
        .in(io_in)
    );
    wire [2:0] _T_280;
    CAT #(.width_a(1), .width_b(2)) cat_308 (
        .y(_T_280),
        .a(_T_278),
        .b(2'h0)
    );
    wire [3:0] _T_281;
    CAT #(.width_a(1), .width_b(3)) cat_309 (
        .y(_T_281),
        .a(_T_276),
        .b(_T_277)
    );
    wire [6:0] _T_282;
    CAT #(.width_a(4), .width_b(3)) cat_310 (
        .y(_T_282),
        .a(_T_281),
        .b(_T_280)
    );
    wire [1:0] _T_283;
    SHR_UNSIGNED #(.width(7), .n(5)) u_shr_311 (
        .y(_T_283),
        .in(_T_282)
    );
    wire [2:0] _T_285;
    BITS #(.width(32), .high(4), .low(2)) bits_312 (
        .y(_T_285),
        .in(io_in)
    );
    wire [4:0] _T_286;
    CAT #(.width_a(2), .width_b(3)) cat_313 (
        .y(_T_286),
        .a(2'h1),
        .b(_T_285)
    );
    wire [2:0] _T_288;
    BITS #(.width(32), .high(9), .low(7)) bits_314 (
        .y(_T_288),
        .in(io_in)
    );
    wire [4:0] _T_289;
    CAT #(.width_a(2), .width_b(3)) cat_315 (
        .y(_T_289),
        .a(2'h1),
        .b(_T_288)
    );
    wire _T_291;
    BITS #(.width(32), .high(5), .low(5)) bits_316 (
        .y(_T_291),
        .in(io_in)
    );
    wire [2:0] _T_292;
    BITS #(.width(32), .high(12), .low(10)) bits_317 (
        .y(_T_292),
        .in(io_in)
    );
    wire _T_293;
    BITS #(.width(32), .high(6), .low(6)) bits_318 (
        .y(_T_293),
        .in(io_in)
    );
    wire [2:0] _T_295;
    CAT #(.width_a(1), .width_b(2)) cat_319 (
        .y(_T_295),
        .a(_T_293),
        .b(2'h0)
    );
    wire [3:0] _T_296;
    CAT #(.width_a(1), .width_b(3)) cat_320 (
        .y(_T_296),
        .a(_T_291),
        .b(_T_292)
    );
    wire [6:0] _T_297;
    CAT #(.width_a(4), .width_b(3)) cat_321 (
        .y(_T_297),
        .a(_T_296),
        .b(_T_295)
    );
    wire [4:0] _T_298;
    BITS #(.width(7), .high(4), .low(0)) bits_322 (
        .y(_T_298),
        .in(_T_297)
    );
    wire [7:0] _T_300;
    CAT #(.width_a(3), .width_b(5)) cat_323 (
        .y(_T_300),
        .a(3'h2),
        .b(_T_298)
    );
    wire [14:0] _T_301;
    CAT #(.width_a(8), .width_b(7)) cat_324 (
        .y(_T_301),
        .a(_T_300),
        .b(7'h23)
    );
    wire [6:0] _T_302;
    CAT #(.width_a(2), .width_b(5)) cat_325 (
        .y(_T_302),
        .a(_T_283),
        .b(_T_286)
    );
    wire [11:0] _T_303;
    CAT #(.width_a(7), .width_b(5)) cat_326 (
        .y(_T_303),
        .a(_T_302),
        .b(_T_289)
    );
    wire [26:0] _T_304;
    CAT #(.width_a(12), .width_b(15)) cat_327 (
        .y(_T_304),
        .a(_T_303),
        .b(_T_301)
    );
    wire [2:0] _T_306;
    BITS #(.width(32), .high(4), .low(2)) bits_328 (
        .y(_T_306),
        .in(io_in)
    );
    wire [4:0] _T_307;
    CAT #(.width_a(2), .width_b(3)) cat_329 (
        .y(_T_307),
        .a(2'h1),
        .b(_T_306)
    );
    wire [2:0] _T_309;
    BITS #(.width(32), .high(9), .low(7)) bits_330 (
        .y(_T_309),
        .in(io_in)
    );
    wire [4:0] _T_310;
    CAT #(.width_a(2), .width_b(3)) cat_331 (
        .y(_T_310),
        .a(2'h1),
        .b(_T_309)
    );
    wire [2:0] _T_312;
    BITS #(.width(32), .high(4), .low(2)) bits_332 (
        .y(_T_312),
        .in(io_in)
    );
    wire [4:0] _T_313;
    CAT #(.width_a(2), .width_b(3)) cat_333 (
        .y(_T_313),
        .a(2'h1),
        .b(_T_312)
    );
    wire [4:0] _T_314;
    BITS #(.width(32), .high(31), .low(27)) bits_334 (
        .y(_T_314),
        .in(io_in)
    );
    wire [31:0] _T_321_bits;
    wire [4:0] _T_321_rd;
    wire [4:0] _T_321_rs1;
    wire [4:0] _T_321_rs2;
    wire [4:0] _T_321_rs3;
    wire [1:0] _T_327;
    BITS #(.width(32), .high(6), .low(5)) bits_335 (
        .y(_T_327),
        .in(io_in)
    );
    wire [2:0] _T_328;
    BITS #(.width(32), .high(12), .low(10)) bits_336 (
        .y(_T_328),
        .in(io_in)
    );
    wire [4:0] _T_330;
    CAT #(.width_a(2), .width_b(3)) cat_337 (
        .y(_T_330),
        .a(_T_327),
        .b(_T_328)
    );
    wire [7:0] _T_331;
    CAT #(.width_a(5), .width_b(3)) cat_338 (
        .y(_T_331),
        .a(_T_330),
        .b(3'h0)
    );
    wire [2:0] _T_332;
    SHR_UNSIGNED #(.width(8), .n(5)) u_shr_339 (
        .y(_T_332),
        .in(_T_331)
    );
    wire [2:0] _T_334;
    BITS #(.width(32), .high(4), .low(2)) bits_340 (
        .y(_T_334),
        .in(io_in)
    );
    wire [4:0] _T_335;
    CAT #(.width_a(2), .width_b(3)) cat_341 (
        .y(_T_335),
        .a(2'h1),
        .b(_T_334)
    );
    wire [2:0] _T_337;
    BITS #(.width(32), .high(9), .low(7)) bits_342 (
        .y(_T_337),
        .in(io_in)
    );
    wire [4:0] _T_338;
    CAT #(.width_a(2), .width_b(3)) cat_343 (
        .y(_T_338),
        .a(2'h1),
        .b(_T_337)
    );
    wire [1:0] _T_340;
    BITS #(.width(32), .high(6), .low(5)) bits_344 (
        .y(_T_340),
        .in(io_in)
    );
    wire [2:0] _T_341;
    BITS #(.width(32), .high(12), .low(10)) bits_345 (
        .y(_T_341),
        .in(io_in)
    );
    wire [4:0] _T_343;
    CAT #(.width_a(2), .width_b(3)) cat_346 (
        .y(_T_343),
        .a(_T_340),
        .b(_T_341)
    );
    wire [7:0] _T_344;
    CAT #(.width_a(5), .width_b(3)) cat_347 (
        .y(_T_344),
        .a(_T_343),
        .b(3'h0)
    );
    wire [4:0] _T_345;
    BITS #(.width(8), .high(4), .low(0)) bits_348 (
        .y(_T_345),
        .in(_T_344)
    );
    wire [7:0] _T_347;
    CAT #(.width_a(3), .width_b(5)) cat_349 (
        .y(_T_347),
        .a(3'h3),
        .b(_T_345)
    );
    wire [14:0] _T_348;
    CAT #(.width_a(8), .width_b(7)) cat_350 (
        .y(_T_348),
        .a(_T_347),
        .b(7'h23)
    );
    wire [7:0] _T_349;
    CAT #(.width_a(3), .width_b(5)) cat_351 (
        .y(_T_349),
        .a(_T_332),
        .b(_T_335)
    );
    wire [12:0] _T_350;
    CAT #(.width_a(8), .width_b(5)) cat_352 (
        .y(_T_350),
        .a(_T_349),
        .b(_T_338)
    );
    wire [27:0] _T_351;
    CAT #(.width_a(13), .width_b(15)) cat_353 (
        .y(_T_351),
        .a(_T_350),
        .b(_T_348)
    );
    wire [2:0] _T_353;
    BITS #(.width(32), .high(4), .low(2)) bits_354 (
        .y(_T_353),
        .in(io_in)
    );
    wire [4:0] _T_354;
    CAT #(.width_a(2), .width_b(3)) cat_355 (
        .y(_T_354),
        .a(2'h1),
        .b(_T_353)
    );
    wire [2:0] _T_356;
    BITS #(.width(32), .high(9), .low(7)) bits_356 (
        .y(_T_356),
        .in(io_in)
    );
    wire [4:0] _T_357;
    CAT #(.width_a(2), .width_b(3)) cat_357 (
        .y(_T_357),
        .a(2'h1),
        .b(_T_356)
    );
    wire [2:0] _T_359;
    BITS #(.width(32), .high(4), .low(2)) bits_358 (
        .y(_T_359),
        .in(io_in)
    );
    wire [4:0] _T_360;
    CAT #(.width_a(2), .width_b(3)) cat_359 (
        .y(_T_360),
        .a(2'h1),
        .b(_T_359)
    );
    wire [4:0] _T_361;
    BITS #(.width(32), .high(31), .low(27)) bits_360 (
        .y(_T_361),
        .in(io_in)
    );
    wire [31:0] _T_368_bits;
    wire [4:0] _T_368_rd;
    wire [4:0] _T_368_rs1;
    wire [4:0] _T_368_rs2;
    wire [4:0] _T_368_rs3;
    wire _T_374;
    BITS #(.width(32), .high(12), .low(12)) bits_361 (
        .y(_T_374),
        .in(io_in)
    );
    wire _T_375;
    BITS #(.width(1), .high(0), .low(0)) bits_362 (
        .y(_T_375),
        .in(_T_374)
    );
    wire [6:0] _T_378;
    MUX_UNSIGNED #(.width(7)) u_mux_363 (
        .y(_T_378),
        .sel(_T_375),
        .a(7'h7F),
        .b(7'h0)
    );
    wire [4:0] _T_379;
    BITS #(.width(32), .high(6), .low(2)) bits_364 (
        .y(_T_379),
        .in(io_in)
    );
    wire [11:0] _T_380;
    CAT #(.width_a(7), .width_b(5)) cat_365 (
        .y(_T_380),
        .a(_T_378),
        .b(_T_379)
    );
    wire [4:0] _T_381;
    BITS #(.width(32), .high(11), .low(7)) bits_366 (
        .y(_T_381),
        .in(io_in)
    );
    wire [4:0] _T_383;
    BITS #(.width(32), .high(11), .low(7)) bits_367 (
        .y(_T_383),
        .in(io_in)
    );
    wire [11:0] _T_385;
    CAT #(.width_a(5), .width_b(7)) cat_368 (
        .y(_T_385),
        .a(_T_383),
        .b(7'h13)
    );
    wire [16:0] _T_386;
    CAT #(.width_a(12), .width_b(5)) cat_369 (
        .y(_T_386),
        .a(_T_380),
        .b(_T_381)
    );
    wire [19:0] _T_387;
    CAT #(.width_a(17), .width_b(3)) cat_370 (
        .y(_T_387),
        .a(_T_386),
        .b(3'h0)
    );
    wire [31:0] _T_388;
    CAT #(.width_a(20), .width_b(12)) cat_371 (
        .y(_T_388),
        .a(_T_387),
        .b(_T_385)
    );
    wire [4:0] _T_389;
    BITS #(.width(32), .high(11), .low(7)) bits_372 (
        .y(_T_389),
        .in(io_in)
    );
    wire [4:0] _T_390;
    BITS #(.width(32), .high(11), .low(7)) bits_373 (
        .y(_T_390),
        .in(io_in)
    );
    wire [2:0] _T_392;
    BITS #(.width(32), .high(4), .low(2)) bits_374 (
        .y(_T_392),
        .in(io_in)
    );
    wire [4:0] _T_393;
    CAT #(.width_a(2), .width_b(3)) cat_375 (
        .y(_T_393),
        .a(2'h1),
        .b(_T_392)
    );
    wire [4:0] _T_394;
    BITS #(.width(32), .high(31), .low(27)) bits_376 (
        .y(_T_394),
        .in(io_in)
    );
    wire [31:0] _T_401_bits;
    wire [4:0] _T_401_rd;
    wire [4:0] _T_401_rs1;
    wire [4:0] _T_401_rs2;
    wire [4:0] _T_401_rs3;
    wire [4:0] _T_407;
    BITS #(.width(32), .high(11), .low(7)) bits_377 (
        .y(_T_407),
        .in(io_in)
    );
    wire _T_409;
    wire [4:0] _WTEMP_31;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_378 (
        .y(_WTEMP_31),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(5)) u_neq_379 (
        .y(_T_409),
        .a(_T_407),
        .b(_WTEMP_31)
    );
    wire [6:0] _T_412;
    MUX_UNSIGNED #(.width(7)) u_mux_380 (
        .y(_T_412),
        .sel(_T_409),
        .a(7'h1B),
        .b(7'h1F)
    );
    wire _T_413;
    BITS #(.width(32), .high(12), .low(12)) bits_381 (
        .y(_T_413),
        .in(io_in)
    );
    wire _T_414;
    BITS #(.width(1), .high(0), .low(0)) bits_382 (
        .y(_T_414),
        .in(_T_413)
    );
    wire [6:0] _T_417;
    MUX_UNSIGNED #(.width(7)) u_mux_383 (
        .y(_T_417),
        .sel(_T_414),
        .a(7'h7F),
        .b(7'h0)
    );
    wire [4:0] _T_418;
    BITS #(.width(32), .high(6), .low(2)) bits_384 (
        .y(_T_418),
        .in(io_in)
    );
    wire [11:0] _T_419;
    CAT #(.width_a(7), .width_b(5)) cat_385 (
        .y(_T_419),
        .a(_T_417),
        .b(_T_418)
    );
    wire [4:0] _T_420;
    BITS #(.width(32), .high(11), .low(7)) bits_386 (
        .y(_T_420),
        .in(io_in)
    );
    wire [4:0] _T_422;
    BITS #(.width(32), .high(11), .low(7)) bits_387 (
        .y(_T_422),
        .in(io_in)
    );
    wire [11:0] _T_423;
    CAT #(.width_a(5), .width_b(7)) cat_388 (
        .y(_T_423),
        .a(_T_422),
        .b(_T_412)
    );
    wire [16:0] _T_424;
    CAT #(.width_a(12), .width_b(5)) cat_389 (
        .y(_T_424),
        .a(_T_419),
        .b(_T_420)
    );
    wire [19:0] _T_425;
    CAT #(.width_a(17), .width_b(3)) cat_390 (
        .y(_T_425),
        .a(_T_424),
        .b(3'h0)
    );
    wire [31:0] _T_426;
    CAT #(.width_a(20), .width_b(12)) cat_391 (
        .y(_T_426),
        .a(_T_425),
        .b(_T_423)
    );
    wire [4:0] _T_427;
    BITS #(.width(32), .high(11), .low(7)) bits_392 (
        .y(_T_427),
        .in(io_in)
    );
    wire [4:0] _T_428;
    BITS #(.width(32), .high(11), .low(7)) bits_393 (
        .y(_T_428),
        .in(io_in)
    );
    wire [2:0] _T_430;
    BITS #(.width(32), .high(4), .low(2)) bits_394 (
        .y(_T_430),
        .in(io_in)
    );
    wire [4:0] _T_431;
    CAT #(.width_a(2), .width_b(3)) cat_395 (
        .y(_T_431),
        .a(2'h1),
        .b(_T_430)
    );
    wire [4:0] _T_432;
    BITS #(.width(32), .high(31), .low(27)) bits_396 (
        .y(_T_432),
        .in(io_in)
    );
    wire [31:0] _T_439_bits;
    wire [4:0] _T_439_rd;
    wire [4:0] _T_439_rs1;
    wire [4:0] _T_439_rs2;
    wire [4:0] _T_439_rs3;
    wire _T_445;
    BITS #(.width(32), .high(12), .low(12)) bits_397 (
        .y(_T_445),
        .in(io_in)
    );
    wire _T_446;
    BITS #(.width(1), .high(0), .low(0)) bits_398 (
        .y(_T_446),
        .in(_T_445)
    );
    wire [6:0] _T_449;
    MUX_UNSIGNED #(.width(7)) u_mux_399 (
        .y(_T_449),
        .sel(_T_446),
        .a(7'h7F),
        .b(7'h0)
    );
    wire [4:0] _T_450;
    BITS #(.width(32), .high(6), .low(2)) bits_400 (
        .y(_T_450),
        .in(io_in)
    );
    wire [11:0] _T_451;
    CAT #(.width_a(7), .width_b(5)) cat_401 (
        .y(_T_451),
        .a(_T_449),
        .b(_T_450)
    );
    wire [4:0] _T_454;
    BITS #(.width(32), .high(11), .low(7)) bits_402 (
        .y(_T_454),
        .in(io_in)
    );
    wire [11:0] _T_456;
    CAT #(.width_a(5), .width_b(7)) cat_403 (
        .y(_T_456),
        .a(_T_454),
        .b(7'h13)
    );
    wire [16:0] _T_457;
    CAT #(.width_a(12), .width_b(5)) cat_404 (
        .y(_T_457),
        .a(_T_451),
        .b(5'h0)
    );
    wire [19:0] _T_458;
    CAT #(.width_a(17), .width_b(3)) cat_405 (
        .y(_T_458),
        .a(_T_457),
        .b(3'h0)
    );
    wire [31:0] _T_459;
    CAT #(.width_a(20), .width_b(12)) cat_406 (
        .y(_T_459),
        .a(_T_458),
        .b(_T_456)
    );
    wire [4:0] _T_460;
    BITS #(.width(32), .high(11), .low(7)) bits_407 (
        .y(_T_460),
        .in(io_in)
    );
    wire [2:0] _T_463;
    BITS #(.width(32), .high(4), .low(2)) bits_408 (
        .y(_T_463),
        .in(io_in)
    );
    wire [4:0] _T_464;
    CAT #(.width_a(2), .width_b(3)) cat_409 (
        .y(_T_464),
        .a(2'h1),
        .b(_T_463)
    );
    wire [4:0] _T_465;
    BITS #(.width(32), .high(31), .low(27)) bits_410 (
        .y(_T_465),
        .in(io_in)
    );
    wire [31:0] _T_472_bits;
    wire [4:0] _T_472_rd;
    wire [4:0] _T_472_rs1;
    wire [4:0] _T_472_rs2;
    wire [4:0] _T_472_rs3;
    wire _T_478;
    BITS #(.width(32), .high(12), .low(12)) bits_411 (
        .y(_T_478),
        .in(io_in)
    );
    wire _T_479;
    BITS #(.width(1), .high(0), .low(0)) bits_412 (
        .y(_T_479),
        .in(_T_478)
    );
    wire [6:0] _T_482;
    MUX_UNSIGNED #(.width(7)) u_mux_413 (
        .y(_T_482),
        .sel(_T_479),
        .a(7'h7F),
        .b(7'h0)
    );
    wire [4:0] _T_483;
    BITS #(.width(32), .high(6), .low(2)) bits_414 (
        .y(_T_483),
        .in(io_in)
    );
    wire [11:0] _T_484;
    CAT #(.width_a(7), .width_b(5)) cat_415 (
        .y(_T_484),
        .a(_T_482),
        .b(_T_483)
    );
    wire _T_486;
    wire [11:0] _WTEMP_32;
    PAD_UNSIGNED #(.width(1), .n(12)) u_pad_416 (
        .y(_WTEMP_32),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(12)) u_neq_417 (
        .y(_T_486),
        .a(_T_484),
        .b(_WTEMP_32)
    );
    wire [6:0] _T_489;
    MUX_UNSIGNED #(.width(7)) u_mux_418 (
        .y(_T_489),
        .sel(_T_486),
        .a(7'h37),
        .b(7'h3F)
    );
    wire _T_490;
    BITS #(.width(32), .high(12), .low(12)) bits_419 (
        .y(_T_490),
        .in(io_in)
    );
    wire _T_491;
    BITS #(.width(1), .high(0), .low(0)) bits_420 (
        .y(_T_491),
        .in(_T_490)
    );
    wire [14:0] _T_494;
    MUX_UNSIGNED #(.width(15)) u_mux_421 (
        .y(_T_494),
        .sel(_T_491),
        .a(15'h7FFF),
        .b(15'h0)
    );
    wire [4:0] _T_495;
    BITS #(.width(32), .high(6), .low(2)) bits_422 (
        .y(_T_495),
        .in(io_in)
    );
    wire [19:0] _T_497;
    CAT #(.width_a(15), .width_b(5)) cat_423 (
        .y(_T_497),
        .a(_T_494),
        .b(_T_495)
    );
    wire [31:0] _T_498;
    CAT #(.width_a(20), .width_b(12)) cat_424 (
        .y(_T_498),
        .a(_T_497),
        .b(12'h0)
    );
    wire [19:0] _T_499;
    BITS #(.width(32), .high(31), .low(12)) bits_425 (
        .y(_T_499),
        .in(_T_498)
    );
    wire [4:0] _T_500;
    BITS #(.width(32), .high(11), .low(7)) bits_426 (
        .y(_T_500),
        .in(io_in)
    );
    wire [24:0] _T_501;
    CAT #(.width_a(20), .width_b(5)) cat_427 (
        .y(_T_501),
        .a(_T_499),
        .b(_T_500)
    );
    wire [31:0] _T_502;
    CAT #(.width_a(25), .width_b(7)) cat_428 (
        .y(_T_502),
        .a(_T_501),
        .b(_T_489)
    );
    wire [4:0] _T_503;
    BITS #(.width(32), .high(11), .low(7)) bits_429 (
        .y(_T_503),
        .in(io_in)
    );
    wire [4:0] _T_504;
    BITS #(.width(32), .high(11), .low(7)) bits_430 (
        .y(_T_504),
        .in(io_in)
    );
    wire [2:0] _T_506;
    BITS #(.width(32), .high(4), .low(2)) bits_431 (
        .y(_T_506),
        .in(io_in)
    );
    wire [4:0] _T_507;
    CAT #(.width_a(2), .width_b(3)) cat_432 (
        .y(_T_507),
        .a(2'h1),
        .b(_T_506)
    );
    wire [4:0] _T_508;
    BITS #(.width(32), .high(31), .low(27)) bits_433 (
        .y(_T_508),
        .in(io_in)
    );
    wire [31:0] _T_515_bits;
    wire [4:0] _T_515_rd;
    wire [4:0] _T_515_rs1;
    wire [4:0] _T_515_rs2;
    wire [4:0] _T_515_rs3;
    wire [4:0] _T_521;
    BITS #(.width(32), .high(11), .low(7)) bits_434 (
        .y(_T_521),
        .in(io_in)
    );
    wire _T_523;
    EQ_UNSIGNED #(.width(5)) u_eq_435 (
        .y(_T_523),
        .a(_T_521),
        .b(5'h0)
    );
    wire [4:0] _T_524;
    BITS #(.width(32), .high(11), .low(7)) bits_436 (
        .y(_T_524),
        .in(io_in)
    );
    wire _T_526;
    EQ_UNSIGNED #(.width(5)) u_eq_437 (
        .y(_T_526),
        .a(_T_524),
        .b(5'h2)
    );
    wire _T_527;
    BITWISEOR #(.width(1)) bitwiseor_438 (
        .y(_T_527),
        .a(_T_523),
        .b(_T_526)
    );
    wire _T_528;
    BITS #(.width(32), .high(12), .low(12)) bits_439 (
        .y(_T_528),
        .in(io_in)
    );
    wire _T_529;
    BITS #(.width(1), .high(0), .low(0)) bits_440 (
        .y(_T_529),
        .in(_T_528)
    );
    wire [6:0] _T_532;
    MUX_UNSIGNED #(.width(7)) u_mux_441 (
        .y(_T_532),
        .sel(_T_529),
        .a(7'h7F),
        .b(7'h0)
    );
    wire [4:0] _T_533;
    BITS #(.width(32), .high(6), .low(2)) bits_442 (
        .y(_T_533),
        .in(io_in)
    );
    wire [11:0] _T_534;
    CAT #(.width_a(7), .width_b(5)) cat_443 (
        .y(_T_534),
        .a(_T_532),
        .b(_T_533)
    );
    wire _T_536;
    wire [11:0] _WTEMP_33;
    PAD_UNSIGNED #(.width(1), .n(12)) u_pad_444 (
        .y(_WTEMP_33),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(12)) u_neq_445 (
        .y(_T_536),
        .a(_T_534),
        .b(_WTEMP_33)
    );
    wire [6:0] _T_539;
    MUX_UNSIGNED #(.width(7)) u_mux_446 (
        .y(_T_539),
        .sel(_T_536),
        .a(7'h13),
        .b(7'h1F)
    );
    wire _T_540;
    BITS #(.width(32), .high(12), .low(12)) bits_447 (
        .y(_T_540),
        .in(io_in)
    );
    wire _T_541;
    BITS #(.width(1), .high(0), .low(0)) bits_448 (
        .y(_T_541),
        .in(_T_540)
    );
    wire [2:0] _T_544;
    MUX_UNSIGNED #(.width(3)) u_mux_449 (
        .y(_T_544),
        .sel(_T_541),
        .a(3'h7),
        .b(3'h0)
    );
    wire [1:0] _T_545;
    BITS #(.width(32), .high(4), .low(3)) bits_450 (
        .y(_T_545),
        .in(io_in)
    );
    wire _T_546;
    BITS #(.width(32), .high(5), .low(5)) bits_451 (
        .y(_T_546),
        .in(io_in)
    );
    wire _T_547;
    BITS #(.width(32), .high(2), .low(2)) bits_452 (
        .y(_T_547),
        .in(io_in)
    );
    wire _T_548;
    BITS #(.width(32), .high(6), .low(6)) bits_453 (
        .y(_T_548),
        .in(io_in)
    );
    wire [1:0] _T_550;
    CAT #(.width_a(1), .width_b(1)) cat_454 (
        .y(_T_550),
        .a(_T_547),
        .b(_T_548)
    );
    wire [5:0] _T_551;
    CAT #(.width_a(2), .width_b(4)) cat_455 (
        .y(_T_551),
        .a(_T_550),
        .b(4'h0)
    );
    wire [4:0] _T_552;
    CAT #(.width_a(3), .width_b(2)) cat_456 (
        .y(_T_552),
        .a(_T_544),
        .b(_T_545)
    );
    wire [5:0] _T_553;
    CAT #(.width_a(5), .width_b(1)) cat_457 (
        .y(_T_553),
        .a(_T_552),
        .b(_T_546)
    );
    wire [11:0] _T_554;
    CAT #(.width_a(6), .width_b(6)) cat_458 (
        .y(_T_554),
        .a(_T_553),
        .b(_T_551)
    );
    wire [4:0] _T_555;
    BITS #(.width(32), .high(11), .low(7)) bits_459 (
        .y(_T_555),
        .in(io_in)
    );
    wire [4:0] _T_557;
    BITS #(.width(32), .high(11), .low(7)) bits_460 (
        .y(_T_557),
        .in(io_in)
    );
    wire [11:0] _T_558;
    CAT #(.width_a(5), .width_b(7)) cat_461 (
        .y(_T_558),
        .a(_T_557),
        .b(_T_539)
    );
    wire [16:0] _T_559;
    CAT #(.width_a(12), .width_b(5)) cat_462 (
        .y(_T_559),
        .a(_T_554),
        .b(_T_555)
    );
    wire [19:0] _T_560;
    CAT #(.width_a(17), .width_b(3)) cat_463 (
        .y(_T_560),
        .a(_T_559),
        .b(3'h0)
    );
    wire [31:0] _T_561;
    CAT #(.width_a(20), .width_b(12)) cat_464 (
        .y(_T_561),
        .a(_T_560),
        .b(_T_558)
    );
    wire [4:0] _T_562;
    BITS #(.width(32), .high(11), .low(7)) bits_465 (
        .y(_T_562),
        .in(io_in)
    );
    wire [4:0] _T_563;
    BITS #(.width(32), .high(11), .low(7)) bits_466 (
        .y(_T_563),
        .in(io_in)
    );
    wire [2:0] _T_565;
    BITS #(.width(32), .high(4), .low(2)) bits_467 (
        .y(_T_565),
        .in(io_in)
    );
    wire [4:0] _T_566;
    CAT #(.width_a(2), .width_b(3)) cat_468 (
        .y(_T_566),
        .a(2'h1),
        .b(_T_565)
    );
    wire [4:0] _T_567;
    BITS #(.width(32), .high(31), .low(27)) bits_469 (
        .y(_T_567),
        .in(io_in)
    );
    wire [31:0] _T_574_bits;
    wire [4:0] _T_574_rd;
    wire [4:0] _T_574_rs1;
    wire [4:0] _T_574_rs2;
    wire [4:0] _T_574_rs3;
    wire [31:0] _T_580_bits;
    MUX_UNSIGNED #(.width(32)) u_mux_470 (
        .y(_T_580_bits),
        .sel(_T_527),
        .a(_T_574_bits),
        .b(_T_515_bits)
    );
    wire [4:0] _T_580_rd;
    MUX_UNSIGNED #(.width(5)) u_mux_471 (
        .y(_T_580_rd),
        .sel(_T_527),
        .a(_T_574_rd),
        .b(_T_515_rd)
    );
    wire [4:0] _T_580_rs1;
    MUX_UNSIGNED #(.width(5)) u_mux_472 (
        .y(_T_580_rs1),
        .sel(_T_527),
        .a(_T_574_rs1),
        .b(_T_515_rs1)
    );
    wire [4:0] _T_580_rs2;
    MUX_UNSIGNED #(.width(5)) u_mux_473 (
        .y(_T_580_rs2),
        .sel(_T_527),
        .a(_T_574_rs2),
        .b(_T_515_rs2)
    );
    wire [4:0] _T_580_rs3;
    MUX_UNSIGNED #(.width(5)) u_mux_474 (
        .y(_T_580_rs3),
        .sel(_T_527),
        .a(_T_574_rs3),
        .b(_T_515_rs3)
    );
    wire _T_586;
    BITS #(.width(32), .high(12), .low(12)) bits_475 (
        .y(_T_586),
        .in(io_in)
    );
    wire [4:0] _T_587;
    BITS #(.width(32), .high(6), .low(2)) bits_476 (
        .y(_T_587),
        .in(io_in)
    );
    wire [5:0] _T_588;
    CAT #(.width_a(1), .width_b(5)) cat_477 (
        .y(_T_588),
        .a(_T_586),
        .b(_T_587)
    );
    wire [2:0] _T_590;
    BITS #(.width(32), .high(9), .low(7)) bits_478 (
        .y(_T_590),
        .in(io_in)
    );
    wire [4:0] _T_591;
    CAT #(.width_a(2), .width_b(3)) cat_479 (
        .y(_T_591),
        .a(2'h1),
        .b(_T_590)
    );
    wire [2:0] _T_594;
    BITS #(.width(32), .high(9), .low(7)) bits_480 (
        .y(_T_594),
        .in(io_in)
    );
    wire [4:0] _T_595;
    CAT #(.width_a(2), .width_b(3)) cat_481 (
        .y(_T_595),
        .a(2'h1),
        .b(_T_594)
    );
    wire [11:0] _T_597;
    CAT #(.width_a(5), .width_b(7)) cat_482 (
        .y(_T_597),
        .a(_T_595),
        .b(7'h13)
    );
    wire [10:0] _T_598;
    CAT #(.width_a(6), .width_b(5)) cat_483 (
        .y(_T_598),
        .a(_T_588),
        .b(_T_591)
    );
    wire [13:0] _T_599;
    CAT #(.width_a(11), .width_b(3)) cat_484 (
        .y(_T_599),
        .a(_T_598),
        .b(3'h5)
    );
    wire [25:0] _T_600;
    CAT #(.width_a(14), .width_b(12)) cat_485 (
        .y(_T_600),
        .a(_T_599),
        .b(_T_597)
    );
    wire _T_601;
    BITS #(.width(32), .high(12), .low(12)) bits_486 (
        .y(_T_601),
        .in(io_in)
    );
    wire [4:0] _T_602;
    BITS #(.width(32), .high(6), .low(2)) bits_487 (
        .y(_T_602),
        .in(io_in)
    );
    wire [5:0] _T_603;
    CAT #(.width_a(1), .width_b(5)) cat_488 (
        .y(_T_603),
        .a(_T_601),
        .b(_T_602)
    );
    wire [2:0] _T_605;
    BITS #(.width(32), .high(9), .low(7)) bits_489 (
        .y(_T_605),
        .in(io_in)
    );
    wire [4:0] _T_606;
    CAT #(.width_a(2), .width_b(3)) cat_490 (
        .y(_T_606),
        .a(2'h1),
        .b(_T_605)
    );
    wire [2:0] _T_609;
    BITS #(.width(32), .high(9), .low(7)) bits_491 (
        .y(_T_609),
        .in(io_in)
    );
    wire [4:0] _T_610;
    CAT #(.width_a(2), .width_b(3)) cat_492 (
        .y(_T_610),
        .a(2'h1),
        .b(_T_609)
    );
    wire [11:0] _T_612;
    CAT #(.width_a(5), .width_b(7)) cat_493 (
        .y(_T_612),
        .a(_T_610),
        .b(7'h13)
    );
    wire [10:0] _T_613;
    CAT #(.width_a(6), .width_b(5)) cat_494 (
        .y(_T_613),
        .a(_T_603),
        .b(_T_606)
    );
    wire [13:0] _T_614;
    CAT #(.width_a(11), .width_b(3)) cat_495 (
        .y(_T_614),
        .a(_T_613),
        .b(3'h5)
    );
    wire [25:0] _T_615;
    CAT #(.width_a(14), .width_b(12)) cat_496 (
        .y(_T_615),
        .a(_T_614),
        .b(_T_612)
    );
    wire [30:0] _T_617;
    wire [30:0] _WTEMP_34;
    PAD_UNSIGNED #(.width(26), .n(31)) u_pad_497 (
        .y(_WTEMP_34),
        .in(_T_615)
    );
    BITWISEOR #(.width(31)) bitwiseor_498 (
        .y(_T_617),
        .a(_WTEMP_34),
        .b(31'h40000000)
    );
    wire _T_618;
    BITS #(.width(32), .high(12), .low(12)) bits_499 (
        .y(_T_618),
        .in(io_in)
    );
    wire _T_619;
    BITS #(.width(1), .high(0), .low(0)) bits_500 (
        .y(_T_619),
        .in(_T_618)
    );
    wire [6:0] _T_622;
    MUX_UNSIGNED #(.width(7)) u_mux_501 (
        .y(_T_622),
        .sel(_T_619),
        .a(7'h7F),
        .b(7'h0)
    );
    wire [4:0] _T_623;
    BITS #(.width(32), .high(6), .low(2)) bits_502 (
        .y(_T_623),
        .in(io_in)
    );
    wire [11:0] _T_624;
    CAT #(.width_a(7), .width_b(5)) cat_503 (
        .y(_T_624),
        .a(_T_622),
        .b(_T_623)
    );
    wire [2:0] _T_626;
    BITS #(.width(32), .high(9), .low(7)) bits_504 (
        .y(_T_626),
        .in(io_in)
    );
    wire [4:0] _T_627;
    CAT #(.width_a(2), .width_b(3)) cat_505 (
        .y(_T_627),
        .a(2'h1),
        .b(_T_626)
    );
    wire [2:0] _T_630;
    BITS #(.width(32), .high(9), .low(7)) bits_506 (
        .y(_T_630),
        .in(io_in)
    );
    wire [4:0] _T_631;
    CAT #(.width_a(2), .width_b(3)) cat_507 (
        .y(_T_631),
        .a(2'h1),
        .b(_T_630)
    );
    wire [11:0] _T_633;
    CAT #(.width_a(5), .width_b(7)) cat_508 (
        .y(_T_633),
        .a(_T_631),
        .b(7'h13)
    );
    wire [16:0] _T_634;
    CAT #(.width_a(12), .width_b(5)) cat_509 (
        .y(_T_634),
        .a(_T_624),
        .b(_T_627)
    );
    wire [19:0] _T_635;
    CAT #(.width_a(17), .width_b(3)) cat_510 (
        .y(_T_635),
        .a(_T_634),
        .b(3'h7)
    );
    wire [31:0] _T_636;
    CAT #(.width_a(20), .width_b(12)) cat_511 (
        .y(_T_636),
        .a(_T_635),
        .b(_T_633)
    );
    wire _T_645;
    BITS #(.width(32), .high(12), .low(12)) bits_512 (
        .y(_T_645),
        .in(io_in)
    );
    wire [1:0] _T_646;
    BITS #(.width(32), .high(6), .low(5)) bits_513 (
        .y(_T_646),
        .in(io_in)
    );
    wire [2:0] _T_647;
    CAT #(.width_a(1), .width_b(2)) cat_514 (
        .y(_T_647),
        .a(_T_645),
        .b(_T_646)
    );
    wire [2:0] _T_649;
    wire [2:0] _WTEMP_35;
    PAD_UNSIGNED #(.width(2), .n(3)) u_pad_515 (
        .y(_WTEMP_35),
        .in(2'h3)
    );
    BITWISEAND #(.width(3)) bitwiseand_516 (
        .y(_T_649),
        .a(_T_647),
        .b(_WTEMP_35)
    );
    wire _T_651;
    GEQ_UNSIGNED #(.width(3)) u_geq_517 (
        .y(_T_651),
        .a(_T_647),
        .b(3'h4)
    );
    wire [2:0] _T_653;
    wire [2:0] _WTEMP_36;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_518 (
        .y(_WTEMP_36),
        .in(1'h1)
    );
    BITWISEAND #(.width(3)) bitwiseand_519 (
        .y(_T_653),
        .a(_T_649),
        .b(_WTEMP_36)
    );
    wire _T_655;
    wire [2:0] _WTEMP_37;
    PAD_UNSIGNED #(.width(2), .n(3)) u_pad_520 (
        .y(_WTEMP_37),
        .in(2'h2)
    );
    GEQ_UNSIGNED #(.width(3)) u_geq_521 (
        .y(_T_655),
        .a(_T_649),
        .b(_WTEMP_37)
    );
    wire [2:0] _T_657;
    assign _T_657 = 3'h0;
    wire _T_659;
    wire [2:0] _WTEMP_38;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_522 (
        .y(_WTEMP_38),
        .in(1'h1)
    );
    GEQ_UNSIGNED #(.width(3)) u_geq_523 (
        .y(_T_659),
        .a(_T_653),
        .b(_WTEMP_38)
    );
    wire [1:0] _T_660;
    MUX_UNSIGNED #(.width(2)) u_mux_524 (
        .y(_T_660),
        .sel(_T_659),
        .a(2'h3),
        .b(2'h2)
    );
    wire [2:0] _T_662;
    assign _T_662 = 3'h0;
    wire _T_664;
    wire [2:0] _WTEMP_39;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_525 (
        .y(_WTEMP_39),
        .in(1'h1)
    );
    GEQ_UNSIGNED #(.width(3)) u_geq_526 (
        .y(_T_664),
        .a(_T_653),
        .b(_WTEMP_39)
    );
    wire _T_665;
    assign _T_665 = 1'h0;
    wire [1:0] _T_666;
    wire [1:0] _WTEMP_40;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_527 (
        .y(_WTEMP_40),
        .in(_T_665)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_528 (
        .y(_T_666),
        .sel(_T_655),
        .a(_T_660),
        .b(_WTEMP_40)
    );
    wire [2:0] _T_668;
    wire [2:0] _WTEMP_41;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_529 (
        .y(_WTEMP_41),
        .in(1'h1)
    );
    BITWISEAND #(.width(3)) bitwiseand_530 (
        .y(_T_668),
        .a(_T_649),
        .b(_WTEMP_41)
    );
    wire _T_670;
    wire [2:0] _WTEMP_42;
    PAD_UNSIGNED #(.width(2), .n(3)) u_pad_531 (
        .y(_WTEMP_42),
        .in(2'h2)
    );
    GEQ_UNSIGNED #(.width(3)) u_geq_532 (
        .y(_T_670),
        .a(_T_649),
        .b(_WTEMP_42)
    );
    wire [2:0] _T_672;
    assign _T_672 = 3'h0;
    wire _T_674;
    wire [2:0] _WTEMP_43;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_533 (
        .y(_WTEMP_43),
        .in(1'h1)
    );
    GEQ_UNSIGNED #(.width(3)) u_geq_534 (
        .y(_T_674),
        .a(_T_668),
        .b(_WTEMP_43)
    );
    wire [2:0] _T_675;
    MUX_UNSIGNED #(.width(3)) u_mux_535 (
        .y(_T_675),
        .sel(_T_674),
        .a(3'h7),
        .b(3'h6)
    );
    wire [2:0] _T_677;
    assign _T_677 = 3'h0;
    wire _T_679;
    wire [2:0] _WTEMP_44;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_536 (
        .y(_WTEMP_44),
        .in(1'h1)
    );
    GEQ_UNSIGNED #(.width(3)) u_geq_537 (
        .y(_T_679),
        .a(_T_668),
        .b(_WTEMP_44)
    );
    wire [2:0] _T_680;
    wire [2:0] _WTEMP_45;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_538 (
        .y(_WTEMP_45),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(3)) u_mux_539 (
        .y(_T_680),
        .sel(_T_679),
        .a(3'h4),
        .b(_WTEMP_45)
    );
    wire [2:0] _T_681;
    MUX_UNSIGNED #(.width(3)) u_mux_540 (
        .y(_T_681),
        .sel(_T_670),
        .a(_T_675),
        .b(_T_680)
    );
    wire [2:0] _T_682;
    wire [2:0] _WTEMP_46;
    PAD_UNSIGNED #(.width(2), .n(3)) u_pad_541 (
        .y(_WTEMP_46),
        .in(_T_666)
    );
    MUX_UNSIGNED #(.width(3)) u_mux_542 (
        .y(_T_682),
        .sel(_T_651),
        .a(_WTEMP_46),
        .b(_T_681)
    );
    wire [1:0] _T_683;
    BITS #(.width(32), .high(6), .low(5)) bits_543 (
        .y(_T_683),
        .in(io_in)
    );
    wire _T_685;
    wire [1:0] _WTEMP_47;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_544 (
        .y(_WTEMP_47),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(2)) u_eq_545 (
        .y(_T_685),
        .a(_T_683),
        .b(_WTEMP_47)
    );
    wire [30:0] _T_688;
    wire [30:0] _WTEMP_48;
    PAD_UNSIGNED #(.width(1), .n(31)) u_pad_546 (
        .y(_WTEMP_48),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(31)) u_mux_547 (
        .y(_T_688),
        .sel(_T_685),
        .a(31'h40000000),
        .b(_WTEMP_48)
    );
    wire _T_689;
    BITS #(.width(32), .high(12), .low(12)) bits_548 (
        .y(_T_689),
        .in(io_in)
    );
    wire [6:0] _T_692;
    MUX_UNSIGNED #(.width(7)) u_mux_549 (
        .y(_T_692),
        .sel(_T_689),
        .a(7'h3B),
        .b(7'h33)
    );
    wire [2:0] _T_694;
    BITS #(.width(32), .high(4), .low(2)) bits_550 (
        .y(_T_694),
        .in(io_in)
    );
    wire [4:0] _T_695;
    CAT #(.width_a(2), .width_b(3)) cat_551 (
        .y(_T_695),
        .a(2'h1),
        .b(_T_694)
    );
    wire [2:0] _T_697;
    BITS #(.width(32), .high(9), .low(7)) bits_552 (
        .y(_T_697),
        .in(io_in)
    );
    wire [4:0] _T_698;
    CAT #(.width_a(2), .width_b(3)) cat_553 (
        .y(_T_698),
        .a(2'h1),
        .b(_T_697)
    );
    wire [2:0] _T_700;
    BITS #(.width(32), .high(9), .low(7)) bits_554 (
        .y(_T_700),
        .in(io_in)
    );
    wire [4:0] _T_701;
    CAT #(.width_a(2), .width_b(3)) cat_555 (
        .y(_T_701),
        .a(2'h1),
        .b(_T_700)
    );
    wire [11:0] _T_702;
    CAT #(.width_a(5), .width_b(7)) cat_556 (
        .y(_T_702),
        .a(_T_701),
        .b(_T_692)
    );
    wire [9:0] _T_703;
    CAT #(.width_a(5), .width_b(5)) cat_557 (
        .y(_T_703),
        .a(_T_695),
        .b(_T_698)
    );
    wire [12:0] _T_704;
    CAT #(.width_a(10), .width_b(3)) cat_558 (
        .y(_T_704),
        .a(_T_703),
        .b(_T_682)
    );
    wire [24:0] _T_705;
    CAT #(.width_a(13), .width_b(12)) cat_559 (
        .y(_T_705),
        .a(_T_704),
        .b(_T_702)
    );
    wire [30:0] _T_706;
    wire [30:0] _WTEMP_49;
    PAD_UNSIGNED #(.width(25), .n(31)) u_pad_560 (
        .y(_WTEMP_49),
        .in(_T_705)
    );
    BITWISEOR #(.width(31)) bitwiseor_561 (
        .y(_T_706),
        .a(_WTEMP_49),
        .b(_T_688)
    );
    wire [1:0] _T_707;
    BITS #(.width(32), .high(11), .low(10)) bits_562 (
        .y(_T_707),
        .in(io_in)
    );
    wire [1:0] _T_709;
    wire [1:0] _WTEMP_50;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_563 (
        .y(_WTEMP_50),
        .in(1'h1)
    );
    BITWISEAND #(.width(2)) bitwiseand_564 (
        .y(_T_709),
        .a(_T_707),
        .b(_WTEMP_50)
    );
    wire _T_711;
    GEQ_UNSIGNED #(.width(2)) u_geq_565 (
        .y(_T_711),
        .a(_T_707),
        .b(2'h2)
    );
    wire [1:0] _T_713;
    assign _T_713 = 2'h0;
    wire _T_715;
    wire [1:0] _WTEMP_51;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_566 (
        .y(_WTEMP_51),
        .in(1'h1)
    );
    GEQ_UNSIGNED #(.width(2)) u_geq_567 (
        .y(_T_715),
        .a(_T_709),
        .b(_WTEMP_51)
    );
    wire [31:0] _T_716;
    wire [31:0] _WTEMP_52;
    PAD_UNSIGNED #(.width(31), .n(32)) u_pad_568 (
        .y(_WTEMP_52),
        .in(_T_706)
    );
    MUX_UNSIGNED #(.width(32)) u_mux_569 (
        .y(_T_716),
        .sel(_T_715),
        .a(_WTEMP_52),
        .b(_T_636)
    );
    wire [1:0] _T_718;
    assign _T_718 = 2'h0;
    wire _T_720;
    wire [1:0] _WTEMP_53;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_570 (
        .y(_WTEMP_53),
        .in(1'h1)
    );
    GEQ_UNSIGNED #(.width(2)) u_geq_571 (
        .y(_T_720),
        .a(_T_709),
        .b(_WTEMP_53)
    );
    wire [30:0] _T_721;
    wire [30:0] _WTEMP_54;
    PAD_UNSIGNED #(.width(26), .n(31)) u_pad_572 (
        .y(_WTEMP_54),
        .in(_T_600)
    );
    MUX_UNSIGNED #(.width(31)) u_mux_573 (
        .y(_T_721),
        .sel(_T_720),
        .a(_T_617),
        .b(_WTEMP_54)
    );
    wire [31:0] _T_722;
    wire [31:0] _WTEMP_55;
    PAD_UNSIGNED #(.width(31), .n(32)) u_pad_574 (
        .y(_WTEMP_55),
        .in(_T_721)
    );
    MUX_UNSIGNED #(.width(32)) u_mux_575 (
        .y(_T_722),
        .sel(_T_711),
        .a(_T_716),
        .b(_WTEMP_55)
    );
    wire [2:0] _T_724;
    BITS #(.width(32), .high(9), .low(7)) bits_576 (
        .y(_T_724),
        .in(io_in)
    );
    wire [4:0] _T_725;
    CAT #(.width_a(2), .width_b(3)) cat_577 (
        .y(_T_725),
        .a(2'h1),
        .b(_T_724)
    );
    wire [2:0] _T_727;
    BITS #(.width(32), .high(9), .low(7)) bits_578 (
        .y(_T_727),
        .in(io_in)
    );
    wire [4:0] _T_728;
    CAT #(.width_a(2), .width_b(3)) cat_579 (
        .y(_T_728),
        .a(2'h1),
        .b(_T_727)
    );
    wire [2:0] _T_730;
    BITS #(.width(32), .high(4), .low(2)) bits_580 (
        .y(_T_730),
        .in(io_in)
    );
    wire [4:0] _T_731;
    CAT #(.width_a(2), .width_b(3)) cat_581 (
        .y(_T_731),
        .a(2'h1),
        .b(_T_730)
    );
    wire [4:0] _T_732;
    BITS #(.width(32), .high(31), .low(27)) bits_582 (
        .y(_T_732),
        .in(io_in)
    );
    wire [31:0] _T_739_bits;
    wire [4:0] _T_739_rd;
    wire [4:0] _T_739_rs1;
    wire [4:0] _T_739_rs2;
    wire [4:0] _T_739_rs3;
    wire _T_745;
    BITS #(.width(32), .high(12), .low(12)) bits_583 (
        .y(_T_745),
        .in(io_in)
    );
    wire _T_746;
    BITS #(.width(1), .high(0), .low(0)) bits_584 (
        .y(_T_746),
        .in(_T_745)
    );
    wire [9:0] _T_749;
    MUX_UNSIGNED #(.width(10)) u_mux_585 (
        .y(_T_749),
        .sel(_T_746),
        .a(10'h3FF),
        .b(10'h0)
    );
    wire _T_750;
    BITS #(.width(32), .high(8), .low(8)) bits_586 (
        .y(_T_750),
        .in(io_in)
    );
    wire [1:0] _T_751;
    BITS #(.width(32), .high(10), .low(9)) bits_587 (
        .y(_T_751),
        .in(io_in)
    );
    wire _T_752;
    BITS #(.width(32), .high(6), .low(6)) bits_588 (
        .y(_T_752),
        .in(io_in)
    );
    wire _T_753;
    BITS #(.width(32), .high(7), .low(7)) bits_589 (
        .y(_T_753),
        .in(io_in)
    );
    wire _T_754;
    BITS #(.width(32), .high(2), .low(2)) bits_590 (
        .y(_T_754),
        .in(io_in)
    );
    wire _T_755;
    BITS #(.width(32), .high(11), .low(11)) bits_591 (
        .y(_T_755),
        .in(io_in)
    );
    wire [2:0] _T_756;
    BITS #(.width(32), .high(5), .low(3)) bits_592 (
        .y(_T_756),
        .in(io_in)
    );
    wire [3:0] _T_758;
    CAT #(.width_a(3), .width_b(1)) cat_593 (
        .y(_T_758),
        .a(_T_756),
        .b(1'h0)
    );
    wire [1:0] _T_759;
    CAT #(.width_a(1), .width_b(1)) cat_594 (
        .y(_T_759),
        .a(_T_754),
        .b(_T_755)
    );
    wire [5:0] _T_760;
    CAT #(.width_a(2), .width_b(4)) cat_595 (
        .y(_T_760),
        .a(_T_759),
        .b(_T_758)
    );
    wire [1:0] _T_761;
    CAT #(.width_a(1), .width_b(1)) cat_596 (
        .y(_T_761),
        .a(_T_752),
        .b(_T_753)
    );
    wire [10:0] _T_762;
    CAT #(.width_a(10), .width_b(1)) cat_597 (
        .y(_T_762),
        .a(_T_749),
        .b(_T_750)
    );
    wire [12:0] _T_763;
    CAT #(.width_a(11), .width_b(2)) cat_598 (
        .y(_T_763),
        .a(_T_762),
        .b(_T_751)
    );
    wire [14:0] _T_764;
    CAT #(.width_a(13), .width_b(2)) cat_599 (
        .y(_T_764),
        .a(_T_763),
        .b(_T_761)
    );
    wire [20:0] _T_765;
    CAT #(.width_a(15), .width_b(6)) cat_600 (
        .y(_T_765),
        .a(_T_764),
        .b(_T_760)
    );
    wire _T_766;
    BITS #(.width(21), .high(20), .low(20)) bits_601 (
        .y(_T_766),
        .in(_T_765)
    );
    wire _T_767;
    BITS #(.width(32), .high(12), .low(12)) bits_602 (
        .y(_T_767),
        .in(io_in)
    );
    wire _T_768;
    BITS #(.width(1), .high(0), .low(0)) bits_603 (
        .y(_T_768),
        .in(_T_767)
    );
    wire [9:0] _T_771;
    MUX_UNSIGNED #(.width(10)) u_mux_604 (
        .y(_T_771),
        .sel(_T_768),
        .a(10'h3FF),
        .b(10'h0)
    );
    wire _T_772;
    BITS #(.width(32), .high(8), .low(8)) bits_605 (
        .y(_T_772),
        .in(io_in)
    );
    wire [1:0] _T_773;
    BITS #(.width(32), .high(10), .low(9)) bits_606 (
        .y(_T_773),
        .in(io_in)
    );
    wire _T_774;
    BITS #(.width(32), .high(6), .low(6)) bits_607 (
        .y(_T_774),
        .in(io_in)
    );
    wire _T_775;
    BITS #(.width(32), .high(7), .low(7)) bits_608 (
        .y(_T_775),
        .in(io_in)
    );
    wire _T_776;
    BITS #(.width(32), .high(2), .low(2)) bits_609 (
        .y(_T_776),
        .in(io_in)
    );
    wire _T_777;
    BITS #(.width(32), .high(11), .low(11)) bits_610 (
        .y(_T_777),
        .in(io_in)
    );
    wire [2:0] _T_778;
    BITS #(.width(32), .high(5), .low(3)) bits_611 (
        .y(_T_778),
        .in(io_in)
    );
    wire [3:0] _T_780;
    CAT #(.width_a(3), .width_b(1)) cat_612 (
        .y(_T_780),
        .a(_T_778),
        .b(1'h0)
    );
    wire [1:0] _T_781;
    CAT #(.width_a(1), .width_b(1)) cat_613 (
        .y(_T_781),
        .a(_T_776),
        .b(_T_777)
    );
    wire [5:0] _T_782;
    CAT #(.width_a(2), .width_b(4)) cat_614 (
        .y(_T_782),
        .a(_T_781),
        .b(_T_780)
    );
    wire [1:0] _T_783;
    CAT #(.width_a(1), .width_b(1)) cat_615 (
        .y(_T_783),
        .a(_T_774),
        .b(_T_775)
    );
    wire [10:0] _T_784;
    CAT #(.width_a(10), .width_b(1)) cat_616 (
        .y(_T_784),
        .a(_T_771),
        .b(_T_772)
    );
    wire [12:0] _T_785;
    CAT #(.width_a(11), .width_b(2)) cat_617 (
        .y(_T_785),
        .a(_T_784),
        .b(_T_773)
    );
    wire [14:0] _T_786;
    CAT #(.width_a(13), .width_b(2)) cat_618 (
        .y(_T_786),
        .a(_T_785),
        .b(_T_783)
    );
    wire [20:0] _T_787;
    CAT #(.width_a(15), .width_b(6)) cat_619 (
        .y(_T_787),
        .a(_T_786),
        .b(_T_782)
    );
    wire [9:0] _T_788;
    BITS #(.width(21), .high(10), .low(1)) bits_620 (
        .y(_T_788),
        .in(_T_787)
    );
    wire _T_789;
    BITS #(.width(32), .high(12), .low(12)) bits_621 (
        .y(_T_789),
        .in(io_in)
    );
    wire _T_790;
    BITS #(.width(1), .high(0), .low(0)) bits_622 (
        .y(_T_790),
        .in(_T_789)
    );
    wire [9:0] _T_793;
    MUX_UNSIGNED #(.width(10)) u_mux_623 (
        .y(_T_793),
        .sel(_T_790),
        .a(10'h3FF),
        .b(10'h0)
    );
    wire _T_794;
    BITS #(.width(32), .high(8), .low(8)) bits_624 (
        .y(_T_794),
        .in(io_in)
    );
    wire [1:0] _T_795;
    BITS #(.width(32), .high(10), .low(9)) bits_625 (
        .y(_T_795),
        .in(io_in)
    );
    wire _T_796;
    BITS #(.width(32), .high(6), .low(6)) bits_626 (
        .y(_T_796),
        .in(io_in)
    );
    wire _T_797;
    BITS #(.width(32), .high(7), .low(7)) bits_627 (
        .y(_T_797),
        .in(io_in)
    );
    wire _T_798;
    BITS #(.width(32), .high(2), .low(2)) bits_628 (
        .y(_T_798),
        .in(io_in)
    );
    wire _T_799;
    BITS #(.width(32), .high(11), .low(11)) bits_629 (
        .y(_T_799),
        .in(io_in)
    );
    wire [2:0] _T_800;
    BITS #(.width(32), .high(5), .low(3)) bits_630 (
        .y(_T_800),
        .in(io_in)
    );
    wire [3:0] _T_802;
    CAT #(.width_a(3), .width_b(1)) cat_631 (
        .y(_T_802),
        .a(_T_800),
        .b(1'h0)
    );
    wire [1:0] _T_803;
    CAT #(.width_a(1), .width_b(1)) cat_632 (
        .y(_T_803),
        .a(_T_798),
        .b(_T_799)
    );
    wire [5:0] _T_804;
    CAT #(.width_a(2), .width_b(4)) cat_633 (
        .y(_T_804),
        .a(_T_803),
        .b(_T_802)
    );
    wire [1:0] _T_805;
    CAT #(.width_a(1), .width_b(1)) cat_634 (
        .y(_T_805),
        .a(_T_796),
        .b(_T_797)
    );
    wire [10:0] _T_806;
    CAT #(.width_a(10), .width_b(1)) cat_635 (
        .y(_T_806),
        .a(_T_793),
        .b(_T_794)
    );
    wire [12:0] _T_807;
    CAT #(.width_a(11), .width_b(2)) cat_636 (
        .y(_T_807),
        .a(_T_806),
        .b(_T_795)
    );
    wire [14:0] _T_808;
    CAT #(.width_a(13), .width_b(2)) cat_637 (
        .y(_T_808),
        .a(_T_807),
        .b(_T_805)
    );
    wire [20:0] _T_809;
    CAT #(.width_a(15), .width_b(6)) cat_638 (
        .y(_T_809),
        .a(_T_808),
        .b(_T_804)
    );
    wire _T_810;
    BITS #(.width(21), .high(11), .low(11)) bits_639 (
        .y(_T_810),
        .in(_T_809)
    );
    wire _T_811;
    BITS #(.width(32), .high(12), .low(12)) bits_640 (
        .y(_T_811),
        .in(io_in)
    );
    wire _T_812;
    BITS #(.width(1), .high(0), .low(0)) bits_641 (
        .y(_T_812),
        .in(_T_811)
    );
    wire [9:0] _T_815;
    MUX_UNSIGNED #(.width(10)) u_mux_642 (
        .y(_T_815),
        .sel(_T_812),
        .a(10'h3FF),
        .b(10'h0)
    );
    wire _T_816;
    BITS #(.width(32), .high(8), .low(8)) bits_643 (
        .y(_T_816),
        .in(io_in)
    );
    wire [1:0] _T_817;
    BITS #(.width(32), .high(10), .low(9)) bits_644 (
        .y(_T_817),
        .in(io_in)
    );
    wire _T_818;
    BITS #(.width(32), .high(6), .low(6)) bits_645 (
        .y(_T_818),
        .in(io_in)
    );
    wire _T_819;
    BITS #(.width(32), .high(7), .low(7)) bits_646 (
        .y(_T_819),
        .in(io_in)
    );
    wire _T_820;
    BITS #(.width(32), .high(2), .low(2)) bits_647 (
        .y(_T_820),
        .in(io_in)
    );
    wire _T_821;
    BITS #(.width(32), .high(11), .low(11)) bits_648 (
        .y(_T_821),
        .in(io_in)
    );
    wire [2:0] _T_822;
    BITS #(.width(32), .high(5), .low(3)) bits_649 (
        .y(_T_822),
        .in(io_in)
    );
    wire [3:0] _T_824;
    CAT #(.width_a(3), .width_b(1)) cat_650 (
        .y(_T_824),
        .a(_T_822),
        .b(1'h0)
    );
    wire [1:0] _T_825;
    CAT #(.width_a(1), .width_b(1)) cat_651 (
        .y(_T_825),
        .a(_T_820),
        .b(_T_821)
    );
    wire [5:0] _T_826;
    CAT #(.width_a(2), .width_b(4)) cat_652 (
        .y(_T_826),
        .a(_T_825),
        .b(_T_824)
    );
    wire [1:0] _T_827;
    CAT #(.width_a(1), .width_b(1)) cat_653 (
        .y(_T_827),
        .a(_T_818),
        .b(_T_819)
    );
    wire [10:0] _T_828;
    CAT #(.width_a(10), .width_b(1)) cat_654 (
        .y(_T_828),
        .a(_T_815),
        .b(_T_816)
    );
    wire [12:0] _T_829;
    CAT #(.width_a(11), .width_b(2)) cat_655 (
        .y(_T_829),
        .a(_T_828),
        .b(_T_817)
    );
    wire [14:0] _T_830;
    CAT #(.width_a(13), .width_b(2)) cat_656 (
        .y(_T_830),
        .a(_T_829),
        .b(_T_827)
    );
    wire [20:0] _T_831;
    CAT #(.width_a(15), .width_b(6)) cat_657 (
        .y(_T_831),
        .a(_T_830),
        .b(_T_826)
    );
    wire [7:0] _T_832;
    BITS #(.width(21), .high(19), .low(12)) bits_658 (
        .y(_T_832),
        .in(_T_831)
    );
    wire [12:0] _T_835;
    CAT #(.width_a(8), .width_b(5)) cat_659 (
        .y(_T_835),
        .a(_T_832),
        .b(5'h0)
    );
    wire [19:0] _T_836;
    CAT #(.width_a(13), .width_b(7)) cat_660 (
        .y(_T_836),
        .a(_T_835),
        .b(7'h6F)
    );
    wire [10:0] _T_837;
    CAT #(.width_a(1), .width_b(10)) cat_661 (
        .y(_T_837),
        .a(_T_766),
        .b(_T_788)
    );
    wire [11:0] _T_838;
    CAT #(.width_a(11), .width_b(1)) cat_662 (
        .y(_T_838),
        .a(_T_837),
        .b(_T_810)
    );
    wire [31:0] _T_839;
    CAT #(.width_a(12), .width_b(20)) cat_663 (
        .y(_T_839),
        .a(_T_838),
        .b(_T_836)
    );
    wire [2:0] _T_842;
    BITS #(.width(32), .high(9), .low(7)) bits_664 (
        .y(_T_842),
        .in(io_in)
    );
    wire [4:0] _T_843;
    CAT #(.width_a(2), .width_b(3)) cat_665 (
        .y(_T_843),
        .a(2'h1),
        .b(_T_842)
    );
    wire [2:0] _T_845;
    BITS #(.width(32), .high(4), .low(2)) bits_666 (
        .y(_T_845),
        .in(io_in)
    );
    wire [4:0] _T_846;
    CAT #(.width_a(2), .width_b(3)) cat_667 (
        .y(_T_846),
        .a(2'h1),
        .b(_T_845)
    );
    wire [4:0] _T_847;
    BITS #(.width(32), .high(31), .low(27)) bits_668 (
        .y(_T_847),
        .in(io_in)
    );
    wire [31:0] _T_854_bits;
    wire [4:0] _T_854_rd;
    wire [4:0] _T_854_rs1;
    wire [4:0] _T_854_rs2;
    wire [4:0] _T_854_rs3;
    wire _T_860;
    BITS #(.width(32), .high(12), .low(12)) bits_669 (
        .y(_T_860),
        .in(io_in)
    );
    wire _T_861;
    BITS #(.width(1), .high(0), .low(0)) bits_670 (
        .y(_T_861),
        .in(_T_860)
    );
    wire [4:0] _T_864;
    MUX_UNSIGNED #(.width(5)) u_mux_671 (
        .y(_T_864),
        .sel(_T_861),
        .a(5'h1F),
        .b(5'h0)
    );
    wire [1:0] _T_865;
    BITS #(.width(32), .high(6), .low(5)) bits_672 (
        .y(_T_865),
        .in(io_in)
    );
    wire _T_866;
    BITS #(.width(32), .high(2), .low(2)) bits_673 (
        .y(_T_866),
        .in(io_in)
    );
    wire [1:0] _T_867;
    BITS #(.width(32), .high(11), .low(10)) bits_674 (
        .y(_T_867),
        .in(io_in)
    );
    wire [1:0] _T_868;
    BITS #(.width(32), .high(4), .low(3)) bits_675 (
        .y(_T_868),
        .in(io_in)
    );
    wire [3:0] _T_870;
    CAT #(.width_a(2), .width_b(2)) cat_676 (
        .y(_T_870),
        .a(_T_867),
        .b(_T_868)
    );
    wire [4:0] _T_871;
    CAT #(.width_a(4), .width_b(1)) cat_677 (
        .y(_T_871),
        .a(_T_870),
        .b(1'h0)
    );
    wire [6:0] _T_872;
    CAT #(.width_a(5), .width_b(2)) cat_678 (
        .y(_T_872),
        .a(_T_864),
        .b(_T_865)
    );
    wire [7:0] _T_873;
    CAT #(.width_a(7), .width_b(1)) cat_679 (
        .y(_T_873),
        .a(_T_872),
        .b(_T_866)
    );
    wire [12:0] _T_874;
    CAT #(.width_a(8), .width_b(5)) cat_680 (
        .y(_T_874),
        .a(_T_873),
        .b(_T_871)
    );
    wire _T_875;
    BITS #(.width(13), .high(12), .low(12)) bits_681 (
        .y(_T_875),
        .in(_T_874)
    );
    wire _T_876;
    BITS #(.width(32), .high(12), .low(12)) bits_682 (
        .y(_T_876),
        .in(io_in)
    );
    wire _T_877;
    BITS #(.width(1), .high(0), .low(0)) bits_683 (
        .y(_T_877),
        .in(_T_876)
    );
    wire [4:0] _T_880;
    MUX_UNSIGNED #(.width(5)) u_mux_684 (
        .y(_T_880),
        .sel(_T_877),
        .a(5'h1F),
        .b(5'h0)
    );
    wire [1:0] _T_881;
    BITS #(.width(32), .high(6), .low(5)) bits_685 (
        .y(_T_881),
        .in(io_in)
    );
    wire _T_882;
    BITS #(.width(32), .high(2), .low(2)) bits_686 (
        .y(_T_882),
        .in(io_in)
    );
    wire [1:0] _T_883;
    BITS #(.width(32), .high(11), .low(10)) bits_687 (
        .y(_T_883),
        .in(io_in)
    );
    wire [1:0] _T_884;
    BITS #(.width(32), .high(4), .low(3)) bits_688 (
        .y(_T_884),
        .in(io_in)
    );
    wire [3:0] _T_886;
    CAT #(.width_a(2), .width_b(2)) cat_689 (
        .y(_T_886),
        .a(_T_883),
        .b(_T_884)
    );
    wire [4:0] _T_887;
    CAT #(.width_a(4), .width_b(1)) cat_690 (
        .y(_T_887),
        .a(_T_886),
        .b(1'h0)
    );
    wire [6:0] _T_888;
    CAT #(.width_a(5), .width_b(2)) cat_691 (
        .y(_T_888),
        .a(_T_880),
        .b(_T_881)
    );
    wire [7:0] _T_889;
    CAT #(.width_a(7), .width_b(1)) cat_692 (
        .y(_T_889),
        .a(_T_888),
        .b(_T_882)
    );
    wire [12:0] _T_890;
    CAT #(.width_a(8), .width_b(5)) cat_693 (
        .y(_T_890),
        .a(_T_889),
        .b(_T_887)
    );
    wire [5:0] _T_891;
    BITS #(.width(13), .high(10), .low(5)) bits_694 (
        .y(_T_891),
        .in(_T_890)
    );
    wire [2:0] _T_894;
    BITS #(.width(32), .high(9), .low(7)) bits_695 (
        .y(_T_894),
        .in(io_in)
    );
    wire [4:0] _T_895;
    CAT #(.width_a(2), .width_b(3)) cat_696 (
        .y(_T_895),
        .a(2'h1),
        .b(_T_894)
    );
    wire _T_897;
    BITS #(.width(32), .high(12), .low(12)) bits_697 (
        .y(_T_897),
        .in(io_in)
    );
    wire _T_898;
    BITS #(.width(1), .high(0), .low(0)) bits_698 (
        .y(_T_898),
        .in(_T_897)
    );
    wire [4:0] _T_901;
    MUX_UNSIGNED #(.width(5)) u_mux_699 (
        .y(_T_901),
        .sel(_T_898),
        .a(5'h1F),
        .b(5'h0)
    );
    wire [1:0] _T_902;
    BITS #(.width(32), .high(6), .low(5)) bits_700 (
        .y(_T_902),
        .in(io_in)
    );
    wire _T_903;
    BITS #(.width(32), .high(2), .low(2)) bits_701 (
        .y(_T_903),
        .in(io_in)
    );
    wire [1:0] _T_904;
    BITS #(.width(32), .high(11), .low(10)) bits_702 (
        .y(_T_904),
        .in(io_in)
    );
    wire [1:0] _T_905;
    BITS #(.width(32), .high(4), .low(3)) bits_703 (
        .y(_T_905),
        .in(io_in)
    );
    wire [3:0] _T_907;
    CAT #(.width_a(2), .width_b(2)) cat_704 (
        .y(_T_907),
        .a(_T_904),
        .b(_T_905)
    );
    wire [4:0] _T_908;
    CAT #(.width_a(4), .width_b(1)) cat_705 (
        .y(_T_908),
        .a(_T_907),
        .b(1'h0)
    );
    wire [6:0] _T_909;
    CAT #(.width_a(5), .width_b(2)) cat_706 (
        .y(_T_909),
        .a(_T_901),
        .b(_T_902)
    );
    wire [7:0] _T_910;
    CAT #(.width_a(7), .width_b(1)) cat_707 (
        .y(_T_910),
        .a(_T_909),
        .b(_T_903)
    );
    wire [12:0] _T_911;
    CAT #(.width_a(8), .width_b(5)) cat_708 (
        .y(_T_911),
        .a(_T_910),
        .b(_T_908)
    );
    wire [3:0] _T_912;
    BITS #(.width(13), .high(4), .low(1)) bits_709 (
        .y(_T_912),
        .in(_T_911)
    );
    wire _T_913;
    BITS #(.width(32), .high(12), .low(12)) bits_710 (
        .y(_T_913),
        .in(io_in)
    );
    wire _T_914;
    BITS #(.width(1), .high(0), .low(0)) bits_711 (
        .y(_T_914),
        .in(_T_913)
    );
    wire [4:0] _T_917;
    MUX_UNSIGNED #(.width(5)) u_mux_712 (
        .y(_T_917),
        .sel(_T_914),
        .a(5'h1F),
        .b(5'h0)
    );
    wire [1:0] _T_918;
    BITS #(.width(32), .high(6), .low(5)) bits_713 (
        .y(_T_918),
        .in(io_in)
    );
    wire _T_919;
    BITS #(.width(32), .high(2), .low(2)) bits_714 (
        .y(_T_919),
        .in(io_in)
    );
    wire [1:0] _T_920;
    BITS #(.width(32), .high(11), .low(10)) bits_715 (
        .y(_T_920),
        .in(io_in)
    );
    wire [1:0] _T_921;
    BITS #(.width(32), .high(4), .low(3)) bits_716 (
        .y(_T_921),
        .in(io_in)
    );
    wire [3:0] _T_923;
    CAT #(.width_a(2), .width_b(2)) cat_717 (
        .y(_T_923),
        .a(_T_920),
        .b(_T_921)
    );
    wire [4:0] _T_924;
    CAT #(.width_a(4), .width_b(1)) cat_718 (
        .y(_T_924),
        .a(_T_923),
        .b(1'h0)
    );
    wire [6:0] _T_925;
    CAT #(.width_a(5), .width_b(2)) cat_719 (
        .y(_T_925),
        .a(_T_917),
        .b(_T_918)
    );
    wire [7:0] _T_926;
    CAT #(.width_a(7), .width_b(1)) cat_720 (
        .y(_T_926),
        .a(_T_925),
        .b(_T_919)
    );
    wire [12:0] _T_927;
    CAT #(.width_a(8), .width_b(5)) cat_721 (
        .y(_T_927),
        .a(_T_926),
        .b(_T_924)
    );
    wire _T_928;
    BITS #(.width(13), .high(11), .low(11)) bits_722 (
        .y(_T_928),
        .in(_T_927)
    );
    wire [7:0] _T_930;
    CAT #(.width_a(1), .width_b(7)) cat_723 (
        .y(_T_930),
        .a(_T_928),
        .b(7'h63)
    );
    wire [6:0] _T_931;
    CAT #(.width_a(3), .width_b(4)) cat_724 (
        .y(_T_931),
        .a(3'h0),
        .b(_T_912)
    );
    wire [14:0] _T_932;
    CAT #(.width_a(7), .width_b(8)) cat_725 (
        .y(_T_932),
        .a(_T_931),
        .b(_T_930)
    );
    wire [9:0] _T_933;
    CAT #(.width_a(5), .width_b(5)) cat_726 (
        .y(_T_933),
        .a(5'h0),
        .b(_T_895)
    );
    wire [6:0] _T_934;
    CAT #(.width_a(1), .width_b(6)) cat_727 (
        .y(_T_934),
        .a(_T_875),
        .b(_T_891)
    );
    wire [16:0] _T_935;
    CAT #(.width_a(7), .width_b(10)) cat_728 (
        .y(_T_935),
        .a(_T_934),
        .b(_T_933)
    );
    wire [31:0] _T_936;
    CAT #(.width_a(17), .width_b(15)) cat_729 (
        .y(_T_936),
        .a(_T_935),
        .b(_T_932)
    );
    wire [2:0] _T_938;
    BITS #(.width(32), .high(9), .low(7)) bits_730 (
        .y(_T_938),
        .in(io_in)
    );
    wire [4:0] _T_939;
    CAT #(.width_a(2), .width_b(3)) cat_731 (
        .y(_T_939),
        .a(2'h1),
        .b(_T_938)
    );
    wire [2:0] _T_941;
    BITS #(.width(32), .high(9), .low(7)) bits_732 (
        .y(_T_941),
        .in(io_in)
    );
    wire [4:0] _T_942;
    CAT #(.width_a(2), .width_b(3)) cat_733 (
        .y(_T_942),
        .a(2'h1),
        .b(_T_941)
    );
    wire [4:0] _T_944;
    BITS #(.width(32), .high(31), .low(27)) bits_734 (
        .y(_T_944),
        .in(io_in)
    );
    wire [31:0] _T_951_bits;
    wire [4:0] _T_951_rd;
    wire [4:0] _T_951_rs1;
    wire [4:0] _T_951_rs2;
    wire [4:0] _T_951_rs3;
    wire _T_957;
    BITS #(.width(32), .high(12), .low(12)) bits_735 (
        .y(_T_957),
        .in(io_in)
    );
    wire _T_958;
    BITS #(.width(1), .high(0), .low(0)) bits_736 (
        .y(_T_958),
        .in(_T_957)
    );
    wire [4:0] _T_961;
    MUX_UNSIGNED #(.width(5)) u_mux_737 (
        .y(_T_961),
        .sel(_T_958),
        .a(5'h1F),
        .b(5'h0)
    );
    wire [1:0] _T_962;
    BITS #(.width(32), .high(6), .low(5)) bits_738 (
        .y(_T_962),
        .in(io_in)
    );
    wire _T_963;
    BITS #(.width(32), .high(2), .low(2)) bits_739 (
        .y(_T_963),
        .in(io_in)
    );
    wire [1:0] _T_964;
    BITS #(.width(32), .high(11), .low(10)) bits_740 (
        .y(_T_964),
        .in(io_in)
    );
    wire [1:0] _T_965;
    BITS #(.width(32), .high(4), .low(3)) bits_741 (
        .y(_T_965),
        .in(io_in)
    );
    wire [3:0] _T_967;
    CAT #(.width_a(2), .width_b(2)) cat_742 (
        .y(_T_967),
        .a(_T_964),
        .b(_T_965)
    );
    wire [4:0] _T_968;
    CAT #(.width_a(4), .width_b(1)) cat_743 (
        .y(_T_968),
        .a(_T_967),
        .b(1'h0)
    );
    wire [6:0] _T_969;
    CAT #(.width_a(5), .width_b(2)) cat_744 (
        .y(_T_969),
        .a(_T_961),
        .b(_T_962)
    );
    wire [7:0] _T_970;
    CAT #(.width_a(7), .width_b(1)) cat_745 (
        .y(_T_970),
        .a(_T_969),
        .b(_T_963)
    );
    wire [12:0] _T_971;
    CAT #(.width_a(8), .width_b(5)) cat_746 (
        .y(_T_971),
        .a(_T_970),
        .b(_T_968)
    );
    wire _T_972;
    BITS #(.width(13), .high(12), .low(12)) bits_747 (
        .y(_T_972),
        .in(_T_971)
    );
    wire _T_973;
    BITS #(.width(32), .high(12), .low(12)) bits_748 (
        .y(_T_973),
        .in(io_in)
    );
    wire _T_974;
    BITS #(.width(1), .high(0), .low(0)) bits_749 (
        .y(_T_974),
        .in(_T_973)
    );
    wire [4:0] _T_977;
    MUX_UNSIGNED #(.width(5)) u_mux_750 (
        .y(_T_977),
        .sel(_T_974),
        .a(5'h1F),
        .b(5'h0)
    );
    wire [1:0] _T_978;
    BITS #(.width(32), .high(6), .low(5)) bits_751 (
        .y(_T_978),
        .in(io_in)
    );
    wire _T_979;
    BITS #(.width(32), .high(2), .low(2)) bits_752 (
        .y(_T_979),
        .in(io_in)
    );
    wire [1:0] _T_980;
    BITS #(.width(32), .high(11), .low(10)) bits_753 (
        .y(_T_980),
        .in(io_in)
    );
    wire [1:0] _T_981;
    BITS #(.width(32), .high(4), .low(3)) bits_754 (
        .y(_T_981),
        .in(io_in)
    );
    wire [3:0] _T_983;
    CAT #(.width_a(2), .width_b(2)) cat_755 (
        .y(_T_983),
        .a(_T_980),
        .b(_T_981)
    );
    wire [4:0] _T_984;
    CAT #(.width_a(4), .width_b(1)) cat_756 (
        .y(_T_984),
        .a(_T_983),
        .b(1'h0)
    );
    wire [6:0] _T_985;
    CAT #(.width_a(5), .width_b(2)) cat_757 (
        .y(_T_985),
        .a(_T_977),
        .b(_T_978)
    );
    wire [7:0] _T_986;
    CAT #(.width_a(7), .width_b(1)) cat_758 (
        .y(_T_986),
        .a(_T_985),
        .b(_T_979)
    );
    wire [12:0] _T_987;
    CAT #(.width_a(8), .width_b(5)) cat_759 (
        .y(_T_987),
        .a(_T_986),
        .b(_T_984)
    );
    wire [5:0] _T_988;
    BITS #(.width(13), .high(10), .low(5)) bits_760 (
        .y(_T_988),
        .in(_T_987)
    );
    wire [2:0] _T_991;
    BITS #(.width(32), .high(9), .low(7)) bits_761 (
        .y(_T_991),
        .in(io_in)
    );
    wire [4:0] _T_992;
    CAT #(.width_a(2), .width_b(3)) cat_762 (
        .y(_T_992),
        .a(2'h1),
        .b(_T_991)
    );
    wire _T_994;
    BITS #(.width(32), .high(12), .low(12)) bits_763 (
        .y(_T_994),
        .in(io_in)
    );
    wire _T_995;
    BITS #(.width(1), .high(0), .low(0)) bits_764 (
        .y(_T_995),
        .in(_T_994)
    );
    wire [4:0] _T_998;
    MUX_UNSIGNED #(.width(5)) u_mux_765 (
        .y(_T_998),
        .sel(_T_995),
        .a(5'h1F),
        .b(5'h0)
    );
    wire [1:0] _T_999;
    BITS #(.width(32), .high(6), .low(5)) bits_766 (
        .y(_T_999),
        .in(io_in)
    );
    wire _T_1000;
    BITS #(.width(32), .high(2), .low(2)) bits_767 (
        .y(_T_1000),
        .in(io_in)
    );
    wire [1:0] _T_1001;
    BITS #(.width(32), .high(11), .low(10)) bits_768 (
        .y(_T_1001),
        .in(io_in)
    );
    wire [1:0] _T_1002;
    BITS #(.width(32), .high(4), .low(3)) bits_769 (
        .y(_T_1002),
        .in(io_in)
    );
    wire [3:0] _T_1004;
    CAT #(.width_a(2), .width_b(2)) cat_770 (
        .y(_T_1004),
        .a(_T_1001),
        .b(_T_1002)
    );
    wire [4:0] _T_1005;
    CAT #(.width_a(4), .width_b(1)) cat_771 (
        .y(_T_1005),
        .a(_T_1004),
        .b(1'h0)
    );
    wire [6:0] _T_1006;
    CAT #(.width_a(5), .width_b(2)) cat_772 (
        .y(_T_1006),
        .a(_T_998),
        .b(_T_999)
    );
    wire [7:0] _T_1007;
    CAT #(.width_a(7), .width_b(1)) cat_773 (
        .y(_T_1007),
        .a(_T_1006),
        .b(_T_1000)
    );
    wire [12:0] _T_1008;
    CAT #(.width_a(8), .width_b(5)) cat_774 (
        .y(_T_1008),
        .a(_T_1007),
        .b(_T_1005)
    );
    wire [3:0] _T_1009;
    BITS #(.width(13), .high(4), .low(1)) bits_775 (
        .y(_T_1009),
        .in(_T_1008)
    );
    wire _T_1010;
    BITS #(.width(32), .high(12), .low(12)) bits_776 (
        .y(_T_1010),
        .in(io_in)
    );
    wire _T_1011;
    BITS #(.width(1), .high(0), .low(0)) bits_777 (
        .y(_T_1011),
        .in(_T_1010)
    );
    wire [4:0] _T_1014;
    MUX_UNSIGNED #(.width(5)) u_mux_778 (
        .y(_T_1014),
        .sel(_T_1011),
        .a(5'h1F),
        .b(5'h0)
    );
    wire [1:0] _T_1015;
    BITS #(.width(32), .high(6), .low(5)) bits_779 (
        .y(_T_1015),
        .in(io_in)
    );
    wire _T_1016;
    BITS #(.width(32), .high(2), .low(2)) bits_780 (
        .y(_T_1016),
        .in(io_in)
    );
    wire [1:0] _T_1017;
    BITS #(.width(32), .high(11), .low(10)) bits_781 (
        .y(_T_1017),
        .in(io_in)
    );
    wire [1:0] _T_1018;
    BITS #(.width(32), .high(4), .low(3)) bits_782 (
        .y(_T_1018),
        .in(io_in)
    );
    wire [3:0] _T_1020;
    CAT #(.width_a(2), .width_b(2)) cat_783 (
        .y(_T_1020),
        .a(_T_1017),
        .b(_T_1018)
    );
    wire [4:0] _T_1021;
    CAT #(.width_a(4), .width_b(1)) cat_784 (
        .y(_T_1021),
        .a(_T_1020),
        .b(1'h0)
    );
    wire [6:0] _T_1022;
    CAT #(.width_a(5), .width_b(2)) cat_785 (
        .y(_T_1022),
        .a(_T_1014),
        .b(_T_1015)
    );
    wire [7:0] _T_1023;
    CAT #(.width_a(7), .width_b(1)) cat_786 (
        .y(_T_1023),
        .a(_T_1022),
        .b(_T_1016)
    );
    wire [12:0] _T_1024;
    CAT #(.width_a(8), .width_b(5)) cat_787 (
        .y(_T_1024),
        .a(_T_1023),
        .b(_T_1021)
    );
    wire _T_1025;
    BITS #(.width(13), .high(11), .low(11)) bits_788 (
        .y(_T_1025),
        .in(_T_1024)
    );
    wire [7:0] _T_1027;
    CAT #(.width_a(1), .width_b(7)) cat_789 (
        .y(_T_1027),
        .a(_T_1025),
        .b(7'h63)
    );
    wire [6:0] _T_1028;
    CAT #(.width_a(3), .width_b(4)) cat_790 (
        .y(_T_1028),
        .a(3'h1),
        .b(_T_1009)
    );
    wire [14:0] _T_1029;
    CAT #(.width_a(7), .width_b(8)) cat_791 (
        .y(_T_1029),
        .a(_T_1028),
        .b(_T_1027)
    );
    wire [9:0] _T_1030;
    CAT #(.width_a(5), .width_b(5)) cat_792 (
        .y(_T_1030),
        .a(5'h0),
        .b(_T_992)
    );
    wire [6:0] _T_1031;
    CAT #(.width_a(1), .width_b(6)) cat_793 (
        .y(_T_1031),
        .a(_T_972),
        .b(_T_988)
    );
    wire [16:0] _T_1032;
    CAT #(.width_a(7), .width_b(10)) cat_794 (
        .y(_T_1032),
        .a(_T_1031),
        .b(_T_1030)
    );
    wire [31:0] _T_1033;
    CAT #(.width_a(17), .width_b(15)) cat_795 (
        .y(_T_1033),
        .a(_T_1032),
        .b(_T_1029)
    );
    wire [2:0] _T_1036;
    BITS #(.width(32), .high(9), .low(7)) bits_796 (
        .y(_T_1036),
        .in(io_in)
    );
    wire [4:0] _T_1037;
    CAT #(.width_a(2), .width_b(3)) cat_797 (
        .y(_T_1037),
        .a(2'h1),
        .b(_T_1036)
    );
    wire [4:0] _T_1039;
    BITS #(.width(32), .high(31), .low(27)) bits_798 (
        .y(_T_1039),
        .in(io_in)
    );
    wire [31:0] _T_1046_bits;
    wire [4:0] _T_1046_rd;
    wire [4:0] _T_1046_rs1;
    wire [4:0] _T_1046_rs2;
    wire [4:0] _T_1046_rs3;
    wire _T_1052;
    BITS #(.width(32), .high(12), .low(12)) bits_799 (
        .y(_T_1052),
        .in(io_in)
    );
    wire [4:0] _T_1053;
    BITS #(.width(32), .high(6), .low(2)) bits_800 (
        .y(_T_1053),
        .in(io_in)
    );
    wire [5:0] _T_1054;
    CAT #(.width_a(1), .width_b(5)) cat_801 (
        .y(_T_1054),
        .a(_T_1052),
        .b(_T_1053)
    );
    wire [4:0] _T_1055;
    BITS #(.width(32), .high(11), .low(7)) bits_802 (
        .y(_T_1055),
        .in(io_in)
    );
    wire [4:0] _T_1057;
    BITS #(.width(32), .high(11), .low(7)) bits_803 (
        .y(_T_1057),
        .in(io_in)
    );
    wire [11:0] _T_1059;
    CAT #(.width_a(5), .width_b(7)) cat_804 (
        .y(_T_1059),
        .a(_T_1057),
        .b(7'h13)
    );
    wire [10:0] _T_1060;
    CAT #(.width_a(6), .width_b(5)) cat_805 (
        .y(_T_1060),
        .a(_T_1054),
        .b(_T_1055)
    );
    wire [13:0] _T_1061;
    CAT #(.width_a(11), .width_b(3)) cat_806 (
        .y(_T_1061),
        .a(_T_1060),
        .b(3'h1)
    );
    wire [25:0] _T_1062;
    CAT #(.width_a(14), .width_b(12)) cat_807 (
        .y(_T_1062),
        .a(_T_1061),
        .b(_T_1059)
    );
    wire [4:0] _T_1063;
    BITS #(.width(32), .high(11), .low(7)) bits_808 (
        .y(_T_1063),
        .in(io_in)
    );
    wire [4:0] _T_1064;
    BITS #(.width(32), .high(11), .low(7)) bits_809 (
        .y(_T_1064),
        .in(io_in)
    );
    wire [4:0] _T_1065;
    BITS #(.width(32), .high(6), .low(2)) bits_810 (
        .y(_T_1065),
        .in(io_in)
    );
    wire [4:0] _T_1066;
    BITS #(.width(32), .high(31), .low(27)) bits_811 (
        .y(_T_1066),
        .in(io_in)
    );
    wire [31:0] _T_1073_bits;
    wire [4:0] _T_1073_rd;
    wire [4:0] _T_1073_rs1;
    wire [4:0] _T_1073_rs2;
    wire [4:0] _T_1073_rs3;
    wire [2:0] _T_1079;
    BITS #(.width(32), .high(4), .low(2)) bits_812 (
        .y(_T_1079),
        .in(io_in)
    );
    wire _T_1080;
    BITS #(.width(32), .high(12), .low(12)) bits_813 (
        .y(_T_1080),
        .in(io_in)
    );
    wire [1:0] _T_1081;
    BITS #(.width(32), .high(6), .low(5)) bits_814 (
        .y(_T_1081),
        .in(io_in)
    );
    wire [4:0] _T_1083;
    CAT #(.width_a(2), .width_b(3)) cat_815 (
        .y(_T_1083),
        .a(_T_1081),
        .b(3'h0)
    );
    wire [3:0] _T_1084;
    CAT #(.width_a(3), .width_b(1)) cat_816 (
        .y(_T_1084),
        .a(_T_1079),
        .b(_T_1080)
    );
    wire [8:0] _T_1085;
    CAT #(.width_a(4), .width_b(5)) cat_817 (
        .y(_T_1085),
        .a(_T_1084),
        .b(_T_1083)
    );
    wire [4:0] _T_1088;
    BITS #(.width(32), .high(11), .low(7)) bits_818 (
        .y(_T_1088),
        .in(io_in)
    );
    wire [11:0] _T_1090;
    CAT #(.width_a(5), .width_b(7)) cat_819 (
        .y(_T_1090),
        .a(_T_1088),
        .b(7'h7)
    );
    wire [13:0] _T_1091;
    CAT #(.width_a(9), .width_b(5)) cat_820 (
        .y(_T_1091),
        .a(_T_1085),
        .b(5'h2)
    );
    wire [16:0] _T_1092;
    CAT #(.width_a(14), .width_b(3)) cat_821 (
        .y(_T_1092),
        .a(_T_1091),
        .b(3'h3)
    );
    wire [28:0] _T_1093;
    CAT #(.width_a(17), .width_b(12)) cat_822 (
        .y(_T_1093),
        .a(_T_1092),
        .b(_T_1090)
    );
    wire [4:0] _T_1094;
    BITS #(.width(32), .high(11), .low(7)) bits_823 (
        .y(_T_1094),
        .in(io_in)
    );
    wire [4:0] _T_1096;
    BITS #(.width(32), .high(6), .low(2)) bits_824 (
        .y(_T_1096),
        .in(io_in)
    );
    wire [4:0] _T_1097;
    BITS #(.width(32), .high(31), .low(27)) bits_825 (
        .y(_T_1097),
        .in(io_in)
    );
    wire [31:0] _T_1104_bits;
    wire [4:0] _T_1104_rd;
    wire [4:0] _T_1104_rs1;
    wire [4:0] _T_1104_rs2;
    wire [4:0] _T_1104_rs3;
    wire [1:0] _T_1110;
    BITS #(.width(32), .high(3), .low(2)) bits_826 (
        .y(_T_1110),
        .in(io_in)
    );
    wire _T_1111;
    BITS #(.width(32), .high(12), .low(12)) bits_827 (
        .y(_T_1111),
        .in(io_in)
    );
    wire [2:0] _T_1112;
    BITS #(.width(32), .high(6), .low(4)) bits_828 (
        .y(_T_1112),
        .in(io_in)
    );
    wire [4:0] _T_1114;
    CAT #(.width_a(3), .width_b(2)) cat_829 (
        .y(_T_1114),
        .a(_T_1112),
        .b(2'h0)
    );
    wire [2:0] _T_1115;
    CAT #(.width_a(2), .width_b(1)) cat_830 (
        .y(_T_1115),
        .a(_T_1110),
        .b(_T_1111)
    );
    wire [7:0] _T_1116;
    CAT #(.width_a(3), .width_b(5)) cat_831 (
        .y(_T_1116),
        .a(_T_1115),
        .b(_T_1114)
    );
    wire [4:0] _T_1119;
    BITS #(.width(32), .high(11), .low(7)) bits_832 (
        .y(_T_1119),
        .in(io_in)
    );
    wire [11:0] _T_1121;
    CAT #(.width_a(5), .width_b(7)) cat_833 (
        .y(_T_1121),
        .a(_T_1119),
        .b(7'h3)
    );
    wire [12:0] _T_1122;
    CAT #(.width_a(8), .width_b(5)) cat_834 (
        .y(_T_1122),
        .a(_T_1116),
        .b(5'h2)
    );
    wire [15:0] _T_1123;
    CAT #(.width_a(13), .width_b(3)) cat_835 (
        .y(_T_1123),
        .a(_T_1122),
        .b(3'h2)
    );
    wire [27:0] _T_1124;
    CAT #(.width_a(16), .width_b(12)) cat_836 (
        .y(_T_1124),
        .a(_T_1123),
        .b(_T_1121)
    );
    wire [4:0] _T_1125;
    BITS #(.width(32), .high(11), .low(7)) bits_837 (
        .y(_T_1125),
        .in(io_in)
    );
    wire [4:0] _T_1127;
    BITS #(.width(32), .high(6), .low(2)) bits_838 (
        .y(_T_1127),
        .in(io_in)
    );
    wire [4:0] _T_1128;
    BITS #(.width(32), .high(31), .low(27)) bits_839 (
        .y(_T_1128),
        .in(io_in)
    );
    wire [31:0] _T_1135_bits;
    wire [4:0] _T_1135_rd;
    wire [4:0] _T_1135_rs1;
    wire [4:0] _T_1135_rs2;
    wire [4:0] _T_1135_rs3;
    wire [2:0] _T_1141;
    BITS #(.width(32), .high(4), .low(2)) bits_840 (
        .y(_T_1141),
        .in(io_in)
    );
    wire _T_1142;
    BITS #(.width(32), .high(12), .low(12)) bits_841 (
        .y(_T_1142),
        .in(io_in)
    );
    wire [1:0] _T_1143;
    BITS #(.width(32), .high(6), .low(5)) bits_842 (
        .y(_T_1143),
        .in(io_in)
    );
    wire [4:0] _T_1145;
    CAT #(.width_a(2), .width_b(3)) cat_843 (
        .y(_T_1145),
        .a(_T_1143),
        .b(3'h0)
    );
    wire [3:0] _T_1146;
    CAT #(.width_a(3), .width_b(1)) cat_844 (
        .y(_T_1146),
        .a(_T_1141),
        .b(_T_1142)
    );
    wire [8:0] _T_1147;
    CAT #(.width_a(4), .width_b(5)) cat_845 (
        .y(_T_1147),
        .a(_T_1146),
        .b(_T_1145)
    );
    wire [4:0] _T_1150;
    BITS #(.width(32), .high(11), .low(7)) bits_846 (
        .y(_T_1150),
        .in(io_in)
    );
    wire [11:0] _T_1152;
    CAT #(.width_a(5), .width_b(7)) cat_847 (
        .y(_T_1152),
        .a(_T_1150),
        .b(7'h3)
    );
    wire [13:0] _T_1153;
    CAT #(.width_a(9), .width_b(5)) cat_848 (
        .y(_T_1153),
        .a(_T_1147),
        .b(5'h2)
    );
    wire [16:0] _T_1154;
    CAT #(.width_a(14), .width_b(3)) cat_849 (
        .y(_T_1154),
        .a(_T_1153),
        .b(3'h3)
    );
    wire [28:0] _T_1155;
    CAT #(.width_a(17), .width_b(12)) cat_850 (
        .y(_T_1155),
        .a(_T_1154),
        .b(_T_1152)
    );
    wire [4:0] _T_1156;
    BITS #(.width(32), .high(11), .low(7)) bits_851 (
        .y(_T_1156),
        .in(io_in)
    );
    wire [4:0] _T_1158;
    BITS #(.width(32), .high(6), .low(2)) bits_852 (
        .y(_T_1158),
        .in(io_in)
    );
    wire [4:0] _T_1159;
    BITS #(.width(32), .high(31), .low(27)) bits_853 (
        .y(_T_1159),
        .in(io_in)
    );
    wire [31:0] _T_1166_bits;
    wire [4:0] _T_1166_rd;
    wire [4:0] _T_1166_rs1;
    wire [4:0] _T_1166_rs2;
    wire [4:0] _T_1166_rs3;
    wire [4:0] _T_1172;
    BITS #(.width(32), .high(6), .low(2)) bits_854 (
        .y(_T_1172),
        .in(io_in)
    );
    wire [4:0] _T_1175;
    BITS #(.width(32), .high(11), .low(7)) bits_855 (
        .y(_T_1175),
        .in(io_in)
    );
    wire [11:0] _T_1177;
    CAT #(.width_a(5), .width_b(7)) cat_856 (
        .y(_T_1177),
        .a(_T_1175),
        .b(7'h33)
    );
    wire [9:0] _T_1178;
    CAT #(.width_a(5), .width_b(5)) cat_857 (
        .y(_T_1178),
        .a(_T_1172),
        .b(5'h0)
    );
    wire [12:0] _T_1179;
    CAT #(.width_a(10), .width_b(3)) cat_858 (
        .y(_T_1179),
        .a(_T_1178),
        .b(3'h0)
    );
    wire [24:0] _T_1180;
    CAT #(.width_a(13), .width_b(12)) cat_859 (
        .y(_T_1180),
        .a(_T_1179),
        .b(_T_1177)
    );
    wire [4:0] _T_1181;
    BITS #(.width(32), .high(11), .low(7)) bits_860 (
        .y(_T_1181),
        .in(io_in)
    );
    wire [4:0] _T_1183;
    BITS #(.width(32), .high(6), .low(2)) bits_861 (
        .y(_T_1183),
        .in(io_in)
    );
    wire [4:0] _T_1184;
    BITS #(.width(32), .high(31), .low(27)) bits_862 (
        .y(_T_1184),
        .in(io_in)
    );
    wire [31:0] _T_1191_bits;
    wire [4:0] _T_1191_rd;
    wire [4:0] _T_1191_rs1;
    wire [4:0] _T_1191_rs2;
    wire [4:0] _T_1191_rs3;
    wire [4:0] _T_1197;
    BITS #(.width(32), .high(6), .low(2)) bits_863 (
        .y(_T_1197),
        .in(io_in)
    );
    wire [4:0] _T_1198;
    BITS #(.width(32), .high(11), .low(7)) bits_864 (
        .y(_T_1198),
        .in(io_in)
    );
    wire [4:0] _T_1200;
    BITS #(.width(32), .high(11), .low(7)) bits_865 (
        .y(_T_1200),
        .in(io_in)
    );
    wire [11:0] _T_1202;
    CAT #(.width_a(5), .width_b(7)) cat_866 (
        .y(_T_1202),
        .a(_T_1200),
        .b(7'h33)
    );
    wire [9:0] _T_1203;
    CAT #(.width_a(5), .width_b(5)) cat_867 (
        .y(_T_1203),
        .a(_T_1197),
        .b(_T_1198)
    );
    wire [12:0] _T_1204;
    CAT #(.width_a(10), .width_b(3)) cat_868 (
        .y(_T_1204),
        .a(_T_1203),
        .b(3'h0)
    );
    wire [24:0] _T_1205;
    CAT #(.width_a(13), .width_b(12)) cat_869 (
        .y(_T_1205),
        .a(_T_1204),
        .b(_T_1202)
    );
    wire [4:0] _T_1206;
    BITS #(.width(32), .high(11), .low(7)) bits_870 (
        .y(_T_1206),
        .in(io_in)
    );
    wire [4:0] _T_1207;
    BITS #(.width(32), .high(11), .low(7)) bits_871 (
        .y(_T_1207),
        .in(io_in)
    );
    wire [4:0] _T_1208;
    BITS #(.width(32), .high(6), .low(2)) bits_872 (
        .y(_T_1208),
        .in(io_in)
    );
    wire [4:0] _T_1209;
    BITS #(.width(32), .high(31), .low(27)) bits_873 (
        .y(_T_1209),
        .in(io_in)
    );
    wire [31:0] _T_1216_bits;
    wire [4:0] _T_1216_rd;
    wire [4:0] _T_1216_rs1;
    wire [4:0] _T_1216_rs2;
    wire [4:0] _T_1216_rs3;
    wire [4:0] _T_1222;
    BITS #(.width(32), .high(6), .low(2)) bits_874 (
        .y(_T_1222),
        .in(io_in)
    );
    wire [4:0] _T_1223;
    BITS #(.width(32), .high(11), .low(7)) bits_875 (
        .y(_T_1223),
        .in(io_in)
    );
    wire [11:0] _T_1227;
    assign _T_1227 = 12'h67;
    wire [9:0] _T_1228;
    CAT #(.width_a(5), .width_b(5)) cat_876 (
        .y(_T_1228),
        .a(_T_1222),
        .b(_T_1223)
    );
    wire [12:0] _T_1229;
    CAT #(.width_a(10), .width_b(3)) cat_877 (
        .y(_T_1229),
        .a(_T_1228),
        .b(3'h0)
    );
    wire [24:0] _T_1230;
    CAT #(.width_a(13), .width_b(12)) cat_878 (
        .y(_T_1230),
        .a(_T_1229),
        .b(_T_1227)
    );
    wire [17:0] _T_1231;
    SHR_UNSIGNED #(.width(25), .n(7)) u_shr_879 (
        .y(_T_1231),
        .in(_T_1230)
    );
    wire [24:0] _T_1233;
    CAT #(.width_a(18), .width_b(7)) cat_880 (
        .y(_T_1233),
        .a(_T_1231),
        .b(7'h1F)
    );
    wire [4:0] _T_1234;
    BITS #(.width(32), .high(11), .low(7)) bits_881 (
        .y(_T_1234),
        .in(io_in)
    );
    wire _T_1236;
    wire [4:0] _WTEMP_56;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_882 (
        .y(_WTEMP_56),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(5)) u_neq_883 (
        .y(_T_1236),
        .a(_T_1234),
        .b(_WTEMP_56)
    );
    wire [24:0] _T_1237;
    MUX_UNSIGNED #(.width(25)) u_mux_884 (
        .y(_T_1237),
        .sel(_T_1236),
        .a(_T_1230),
        .b(_T_1233)
    );
    wire [4:0] _T_1239;
    BITS #(.width(32), .high(11), .low(7)) bits_885 (
        .y(_T_1239),
        .in(io_in)
    );
    wire [4:0] _T_1240;
    BITS #(.width(32), .high(6), .low(2)) bits_886 (
        .y(_T_1240),
        .in(io_in)
    );
    wire [4:0] _T_1241;
    BITS #(.width(32), .high(31), .low(27)) bits_887 (
        .y(_T_1241),
        .in(io_in)
    );
    wire [31:0] _T_1248_bits;
    wire [4:0] _T_1248_rd;
    wire [4:0] _T_1248_rs1;
    wire [4:0] _T_1248_rs2;
    wire [4:0] _T_1248_rs3;
    wire [4:0] _T_1254;
    BITS #(.width(32), .high(6), .low(2)) bits_888 (
        .y(_T_1254),
        .in(io_in)
    );
    wire _T_1256;
    wire [4:0] _WTEMP_57;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_889 (
        .y(_WTEMP_57),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(5)) u_neq_890 (
        .y(_T_1256),
        .a(_T_1254),
        .b(_WTEMP_57)
    );
    wire [31:0] _T_1257_bits;
    MUX_UNSIGNED #(.width(32)) u_mux_891 (
        .y(_T_1257_bits),
        .sel(_T_1256),
        .a(_T_1191_bits),
        .b(_T_1248_bits)
    );
    wire [4:0] _T_1257_rd;
    MUX_UNSIGNED #(.width(5)) u_mux_892 (
        .y(_T_1257_rd),
        .sel(_T_1256),
        .a(_T_1191_rd),
        .b(_T_1248_rd)
    );
    wire [4:0] _T_1257_rs1;
    MUX_UNSIGNED #(.width(5)) u_mux_893 (
        .y(_T_1257_rs1),
        .sel(_T_1256),
        .a(_T_1191_rs1),
        .b(_T_1248_rs1)
    );
    wire [4:0] _T_1257_rs2;
    MUX_UNSIGNED #(.width(5)) u_mux_894 (
        .y(_T_1257_rs2),
        .sel(_T_1256),
        .a(_T_1191_rs2),
        .b(_T_1248_rs2)
    );
    wire [4:0] _T_1257_rs3;
    MUX_UNSIGNED #(.width(5)) u_mux_895 (
        .y(_T_1257_rs3),
        .sel(_T_1256),
        .a(_T_1191_rs3),
        .b(_T_1248_rs3)
    );
    wire [4:0] _T_1263;
    BITS #(.width(32), .high(6), .low(2)) bits_896 (
        .y(_T_1263),
        .in(io_in)
    );
    wire [4:0] _T_1264;
    BITS #(.width(32), .high(11), .low(7)) bits_897 (
        .y(_T_1264),
        .in(io_in)
    );
    wire [11:0] _T_1268;
    assign _T_1268 = 12'hE7;
    wire [9:0] _T_1269;
    CAT #(.width_a(5), .width_b(5)) cat_898 (
        .y(_T_1269),
        .a(_T_1263),
        .b(_T_1264)
    );
    wire [12:0] _T_1270;
    CAT #(.width_a(10), .width_b(3)) cat_899 (
        .y(_T_1270),
        .a(_T_1269),
        .b(3'h0)
    );
    wire [24:0] _T_1271;
    CAT #(.width_a(13), .width_b(12)) cat_900 (
        .y(_T_1271),
        .a(_T_1270),
        .b(_T_1268)
    );
    wire [17:0] _T_1272;
    SHR_UNSIGNED #(.width(25), .n(7)) u_shr_901 (
        .y(_T_1272),
        .in(_T_1230)
    );
    wire [24:0] _T_1274;
    CAT #(.width_a(18), .width_b(7)) cat_902 (
        .y(_T_1274),
        .a(_T_1272),
        .b(7'h73)
    );
    wire [24:0] _T_1276;
    wire [24:0] _WTEMP_58;
    PAD_UNSIGNED #(.width(21), .n(25)) u_pad_903 (
        .y(_WTEMP_58),
        .in(21'h100000)
    );
    BITWISEOR #(.width(25)) bitwiseor_904 (
        .y(_T_1276),
        .a(_T_1274),
        .b(_WTEMP_58)
    );
    wire [4:0] _T_1277;
    BITS #(.width(32), .high(11), .low(7)) bits_905 (
        .y(_T_1277),
        .in(io_in)
    );
    wire _T_1279;
    wire [4:0] _WTEMP_59;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_906 (
        .y(_WTEMP_59),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(5)) u_neq_907 (
        .y(_T_1279),
        .a(_T_1277),
        .b(_WTEMP_59)
    );
    wire [24:0] _T_1280;
    MUX_UNSIGNED #(.width(25)) u_mux_908 (
        .y(_T_1280),
        .sel(_T_1279),
        .a(_T_1271),
        .b(_T_1276)
    );
    wire [4:0] _T_1282;
    BITS #(.width(32), .high(11), .low(7)) bits_909 (
        .y(_T_1282),
        .in(io_in)
    );
    wire [4:0] _T_1283;
    BITS #(.width(32), .high(6), .low(2)) bits_910 (
        .y(_T_1283),
        .in(io_in)
    );
    wire [4:0] _T_1284;
    BITS #(.width(32), .high(31), .low(27)) bits_911 (
        .y(_T_1284),
        .in(io_in)
    );
    wire [31:0] _T_1291_bits;
    wire [4:0] _T_1291_rd;
    wire [4:0] _T_1291_rs1;
    wire [4:0] _T_1291_rs2;
    wire [4:0] _T_1291_rs3;
    wire [4:0] _T_1297;
    BITS #(.width(32), .high(6), .low(2)) bits_912 (
        .y(_T_1297),
        .in(io_in)
    );
    wire _T_1299;
    wire [4:0] _WTEMP_60;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_913 (
        .y(_WTEMP_60),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(5)) u_neq_914 (
        .y(_T_1299),
        .a(_T_1297),
        .b(_WTEMP_60)
    );
    wire [31:0] _T_1300_bits;
    MUX_UNSIGNED #(.width(32)) u_mux_915 (
        .y(_T_1300_bits),
        .sel(_T_1299),
        .a(_T_1216_bits),
        .b(_T_1291_bits)
    );
    wire [4:0] _T_1300_rd;
    MUX_UNSIGNED #(.width(5)) u_mux_916 (
        .y(_T_1300_rd),
        .sel(_T_1299),
        .a(_T_1216_rd),
        .b(_T_1291_rd)
    );
    wire [4:0] _T_1300_rs1;
    MUX_UNSIGNED #(.width(5)) u_mux_917 (
        .y(_T_1300_rs1),
        .sel(_T_1299),
        .a(_T_1216_rs1),
        .b(_T_1291_rs1)
    );
    wire [4:0] _T_1300_rs2;
    MUX_UNSIGNED #(.width(5)) u_mux_918 (
        .y(_T_1300_rs2),
        .sel(_T_1299),
        .a(_T_1216_rs2),
        .b(_T_1291_rs2)
    );
    wire [4:0] _T_1300_rs3;
    MUX_UNSIGNED #(.width(5)) u_mux_919 (
        .y(_T_1300_rs3),
        .sel(_T_1299),
        .a(_T_1216_rs3),
        .b(_T_1291_rs3)
    );
    wire _T_1306;
    BITS #(.width(32), .high(12), .low(12)) bits_920 (
        .y(_T_1306),
        .in(io_in)
    );
    wire [31:0] _T_1307_bits;
    MUX_UNSIGNED #(.width(32)) u_mux_921 (
        .y(_T_1307_bits),
        .sel(_T_1306),
        .a(_T_1300_bits),
        .b(_T_1257_bits)
    );
    wire [4:0] _T_1307_rd;
    MUX_UNSIGNED #(.width(5)) u_mux_922 (
        .y(_T_1307_rd),
        .sel(_T_1306),
        .a(_T_1300_rd),
        .b(_T_1257_rd)
    );
    wire [4:0] _T_1307_rs1;
    MUX_UNSIGNED #(.width(5)) u_mux_923 (
        .y(_T_1307_rs1),
        .sel(_T_1306),
        .a(_T_1300_rs1),
        .b(_T_1257_rs1)
    );
    wire [4:0] _T_1307_rs2;
    MUX_UNSIGNED #(.width(5)) u_mux_924 (
        .y(_T_1307_rs2),
        .sel(_T_1306),
        .a(_T_1300_rs2),
        .b(_T_1257_rs2)
    );
    wire [4:0] _T_1307_rs3;
    MUX_UNSIGNED #(.width(5)) u_mux_925 (
        .y(_T_1307_rs3),
        .sel(_T_1306),
        .a(_T_1300_rs3),
        .b(_T_1257_rs3)
    );
    wire [2:0] _T_1313;
    BITS #(.width(32), .high(9), .low(7)) bits_926 (
        .y(_T_1313),
        .in(io_in)
    );
    wire [2:0] _T_1314;
    BITS #(.width(32), .high(12), .low(10)) bits_927 (
        .y(_T_1314),
        .in(io_in)
    );
    wire [5:0] _T_1316;
    CAT #(.width_a(3), .width_b(3)) cat_928 (
        .y(_T_1316),
        .a(_T_1313),
        .b(_T_1314)
    );
    wire [8:0] _T_1317;
    CAT #(.width_a(6), .width_b(3)) cat_929 (
        .y(_T_1317),
        .a(_T_1316),
        .b(3'h0)
    );
    wire [3:0] _T_1318;
    SHR_UNSIGNED #(.width(9), .n(5)) u_shr_930 (
        .y(_T_1318),
        .in(_T_1317)
    );
    wire [4:0] _T_1319;
    BITS #(.width(32), .high(6), .low(2)) bits_931 (
        .y(_T_1319),
        .in(io_in)
    );
    wire [2:0] _T_1322;
    BITS #(.width(32), .high(9), .low(7)) bits_932 (
        .y(_T_1322),
        .in(io_in)
    );
    wire [2:0] _T_1323;
    BITS #(.width(32), .high(12), .low(10)) bits_933 (
        .y(_T_1323),
        .in(io_in)
    );
    wire [5:0] _T_1325;
    CAT #(.width_a(3), .width_b(3)) cat_934 (
        .y(_T_1325),
        .a(_T_1322),
        .b(_T_1323)
    );
    wire [8:0] _T_1326;
    CAT #(.width_a(6), .width_b(3)) cat_935 (
        .y(_T_1326),
        .a(_T_1325),
        .b(3'h0)
    );
    wire [4:0] _T_1327;
    BITS #(.width(9), .high(4), .low(0)) bits_936 (
        .y(_T_1327),
        .in(_T_1326)
    );
    wire [7:0] _T_1329;
    CAT #(.width_a(3), .width_b(5)) cat_937 (
        .y(_T_1329),
        .a(3'h3),
        .b(_T_1327)
    );
    wire [14:0] _T_1330;
    CAT #(.width_a(8), .width_b(7)) cat_938 (
        .y(_T_1330),
        .a(_T_1329),
        .b(7'h27)
    );
    wire [8:0] _T_1331;
    CAT #(.width_a(4), .width_b(5)) cat_939 (
        .y(_T_1331),
        .a(_T_1318),
        .b(_T_1319)
    );
    wire [13:0] _T_1332;
    CAT #(.width_a(9), .width_b(5)) cat_940 (
        .y(_T_1332),
        .a(_T_1331),
        .b(5'h2)
    );
    wire [28:0] _T_1333;
    CAT #(.width_a(14), .width_b(15)) cat_941 (
        .y(_T_1333),
        .a(_T_1332),
        .b(_T_1330)
    );
    wire [4:0] _T_1334;
    BITS #(.width(32), .high(11), .low(7)) bits_942 (
        .y(_T_1334),
        .in(io_in)
    );
    wire [4:0] _T_1336;
    BITS #(.width(32), .high(6), .low(2)) bits_943 (
        .y(_T_1336),
        .in(io_in)
    );
    wire [4:0] _T_1337;
    BITS #(.width(32), .high(31), .low(27)) bits_944 (
        .y(_T_1337),
        .in(io_in)
    );
    wire [31:0] _T_1344_bits;
    wire [4:0] _T_1344_rd;
    wire [4:0] _T_1344_rs1;
    wire [4:0] _T_1344_rs2;
    wire [4:0] _T_1344_rs3;
    wire [1:0] _T_1350;
    BITS #(.width(32), .high(8), .low(7)) bits_945 (
        .y(_T_1350),
        .in(io_in)
    );
    wire [3:0] _T_1351;
    BITS #(.width(32), .high(12), .low(9)) bits_946 (
        .y(_T_1351),
        .in(io_in)
    );
    wire [5:0] _T_1353;
    CAT #(.width_a(2), .width_b(4)) cat_947 (
        .y(_T_1353),
        .a(_T_1350),
        .b(_T_1351)
    );
    wire [7:0] _T_1354;
    CAT #(.width_a(6), .width_b(2)) cat_948 (
        .y(_T_1354),
        .a(_T_1353),
        .b(2'h0)
    );
    wire [2:0] _T_1355;
    SHR_UNSIGNED #(.width(8), .n(5)) u_shr_949 (
        .y(_T_1355),
        .in(_T_1354)
    );
    wire [4:0] _T_1356;
    BITS #(.width(32), .high(6), .low(2)) bits_950 (
        .y(_T_1356),
        .in(io_in)
    );
    wire [1:0] _T_1359;
    BITS #(.width(32), .high(8), .low(7)) bits_951 (
        .y(_T_1359),
        .in(io_in)
    );
    wire [3:0] _T_1360;
    BITS #(.width(32), .high(12), .low(9)) bits_952 (
        .y(_T_1360),
        .in(io_in)
    );
    wire [5:0] _T_1362;
    CAT #(.width_a(2), .width_b(4)) cat_953 (
        .y(_T_1362),
        .a(_T_1359),
        .b(_T_1360)
    );
    wire [7:0] _T_1363;
    CAT #(.width_a(6), .width_b(2)) cat_954 (
        .y(_T_1363),
        .a(_T_1362),
        .b(2'h0)
    );
    wire [4:0] _T_1364;
    BITS #(.width(8), .high(4), .low(0)) bits_955 (
        .y(_T_1364),
        .in(_T_1363)
    );
    wire [7:0] _T_1366;
    CAT #(.width_a(3), .width_b(5)) cat_956 (
        .y(_T_1366),
        .a(3'h2),
        .b(_T_1364)
    );
    wire [14:0] _T_1367;
    CAT #(.width_a(8), .width_b(7)) cat_957 (
        .y(_T_1367),
        .a(_T_1366),
        .b(7'h23)
    );
    wire [7:0] _T_1368;
    CAT #(.width_a(3), .width_b(5)) cat_958 (
        .y(_T_1368),
        .a(_T_1355),
        .b(_T_1356)
    );
    wire [12:0] _T_1369;
    CAT #(.width_a(8), .width_b(5)) cat_959 (
        .y(_T_1369),
        .a(_T_1368),
        .b(5'h2)
    );
    wire [27:0] _T_1370;
    CAT #(.width_a(13), .width_b(15)) cat_960 (
        .y(_T_1370),
        .a(_T_1369),
        .b(_T_1367)
    );
    wire [4:0] _T_1371;
    BITS #(.width(32), .high(11), .low(7)) bits_961 (
        .y(_T_1371),
        .in(io_in)
    );
    wire [4:0] _T_1373;
    BITS #(.width(32), .high(6), .low(2)) bits_962 (
        .y(_T_1373),
        .in(io_in)
    );
    wire [4:0] _T_1374;
    BITS #(.width(32), .high(31), .low(27)) bits_963 (
        .y(_T_1374),
        .in(io_in)
    );
    wire [31:0] _T_1381_bits;
    wire [4:0] _T_1381_rd;
    wire [4:0] _T_1381_rs1;
    wire [4:0] _T_1381_rs2;
    wire [4:0] _T_1381_rs3;
    wire [2:0] _T_1387;
    BITS #(.width(32), .high(9), .low(7)) bits_964 (
        .y(_T_1387),
        .in(io_in)
    );
    wire [2:0] _T_1388;
    BITS #(.width(32), .high(12), .low(10)) bits_965 (
        .y(_T_1388),
        .in(io_in)
    );
    wire [5:0] _T_1390;
    CAT #(.width_a(3), .width_b(3)) cat_966 (
        .y(_T_1390),
        .a(_T_1387),
        .b(_T_1388)
    );
    wire [8:0] _T_1391;
    CAT #(.width_a(6), .width_b(3)) cat_967 (
        .y(_T_1391),
        .a(_T_1390),
        .b(3'h0)
    );
    wire [3:0] _T_1392;
    SHR_UNSIGNED #(.width(9), .n(5)) u_shr_968 (
        .y(_T_1392),
        .in(_T_1391)
    );
    wire [4:0] _T_1393;
    BITS #(.width(32), .high(6), .low(2)) bits_969 (
        .y(_T_1393),
        .in(io_in)
    );
    wire [2:0] _T_1396;
    BITS #(.width(32), .high(9), .low(7)) bits_970 (
        .y(_T_1396),
        .in(io_in)
    );
    wire [2:0] _T_1397;
    BITS #(.width(32), .high(12), .low(10)) bits_971 (
        .y(_T_1397),
        .in(io_in)
    );
    wire [5:0] _T_1399;
    CAT #(.width_a(3), .width_b(3)) cat_972 (
        .y(_T_1399),
        .a(_T_1396),
        .b(_T_1397)
    );
    wire [8:0] _T_1400;
    CAT #(.width_a(6), .width_b(3)) cat_973 (
        .y(_T_1400),
        .a(_T_1399),
        .b(3'h0)
    );
    wire [4:0] _T_1401;
    BITS #(.width(9), .high(4), .low(0)) bits_974 (
        .y(_T_1401),
        .in(_T_1400)
    );
    wire [7:0] _T_1403;
    CAT #(.width_a(3), .width_b(5)) cat_975 (
        .y(_T_1403),
        .a(3'h3),
        .b(_T_1401)
    );
    wire [14:0] _T_1404;
    CAT #(.width_a(8), .width_b(7)) cat_976 (
        .y(_T_1404),
        .a(_T_1403),
        .b(7'h23)
    );
    wire [8:0] _T_1405;
    CAT #(.width_a(4), .width_b(5)) cat_977 (
        .y(_T_1405),
        .a(_T_1392),
        .b(_T_1393)
    );
    wire [13:0] _T_1406;
    CAT #(.width_a(9), .width_b(5)) cat_978 (
        .y(_T_1406),
        .a(_T_1405),
        .b(5'h2)
    );
    wire [28:0] _T_1407;
    CAT #(.width_a(14), .width_b(15)) cat_979 (
        .y(_T_1407),
        .a(_T_1406),
        .b(_T_1404)
    );
    wire [4:0] _T_1408;
    BITS #(.width(32), .high(11), .low(7)) bits_980 (
        .y(_T_1408),
        .in(io_in)
    );
    wire [4:0] _T_1410;
    BITS #(.width(32), .high(6), .low(2)) bits_981 (
        .y(_T_1410),
        .in(io_in)
    );
    wire [4:0] _T_1411;
    BITS #(.width(32), .high(31), .low(27)) bits_982 (
        .y(_T_1411),
        .in(io_in)
    );
    wire [31:0] _T_1418_bits;
    wire [4:0] _T_1418_rd;
    wire [4:0] _T_1418_rs1;
    wire [4:0] _T_1418_rs2;
    wire [4:0] _T_1418_rs3;
    wire [4:0] _T_1424;
    BITS #(.width(32), .high(11), .low(7)) bits_983 (
        .y(_T_1424),
        .in(io_in)
    );
    wire [4:0] _T_1425;
    BITS #(.width(32), .high(19), .low(15)) bits_984 (
        .y(_T_1425),
        .in(io_in)
    );
    wire [4:0] _T_1426;
    BITS #(.width(32), .high(24), .low(20)) bits_985 (
        .y(_T_1426),
        .in(io_in)
    );
    wire [4:0] _T_1427;
    BITS #(.width(32), .high(31), .low(27)) bits_986 (
        .y(_T_1427),
        .in(io_in)
    );
    wire [31:0] _T_1434_bits;
    wire [4:0] _T_1434_rd;
    wire [4:0] _T_1434_rs1;
    wire [4:0] _T_1434_rs2;
    wire [4:0] _T_1434_rs3;
    wire [4:0] _T_1440;
    BITS #(.width(32), .high(11), .low(7)) bits_987 (
        .y(_T_1440),
        .in(io_in)
    );
    wire [4:0] _T_1441;
    BITS #(.width(32), .high(19), .low(15)) bits_988 (
        .y(_T_1441),
        .in(io_in)
    );
    wire [4:0] _T_1442;
    BITS #(.width(32), .high(24), .low(20)) bits_989 (
        .y(_T_1442),
        .in(io_in)
    );
    wire [4:0] _T_1443;
    BITS #(.width(32), .high(31), .low(27)) bits_990 (
        .y(_T_1443),
        .in(io_in)
    );
    wire [31:0] _T_1450_bits;
    wire [4:0] _T_1450_rd;
    wire [4:0] _T_1450_rs1;
    wire [4:0] _T_1450_rs2;
    wire [4:0] _T_1450_rs3;
    wire [4:0] _T_1456;
    BITS #(.width(32), .high(11), .low(7)) bits_991 (
        .y(_T_1456),
        .in(io_in)
    );
    wire [4:0] _T_1457;
    BITS #(.width(32), .high(19), .low(15)) bits_992 (
        .y(_T_1457),
        .in(io_in)
    );
    wire [4:0] _T_1458;
    BITS #(.width(32), .high(24), .low(20)) bits_993 (
        .y(_T_1458),
        .in(io_in)
    );
    wire [4:0] _T_1459;
    BITS #(.width(32), .high(31), .low(27)) bits_994 (
        .y(_T_1459),
        .in(io_in)
    );
    wire [31:0] _T_1466_bits;
    wire [4:0] _T_1466_rd;
    wire [4:0] _T_1466_rs1;
    wire [4:0] _T_1466_rs2;
    wire [4:0] _T_1466_rs3;
    wire [4:0] _T_1472;
    BITS #(.width(32), .high(11), .low(7)) bits_995 (
        .y(_T_1472),
        .in(io_in)
    );
    wire [4:0] _T_1473;
    BITS #(.width(32), .high(19), .low(15)) bits_996 (
        .y(_T_1473),
        .in(io_in)
    );
    wire [4:0] _T_1474;
    BITS #(.width(32), .high(24), .low(20)) bits_997 (
        .y(_T_1474),
        .in(io_in)
    );
    wire [4:0] _T_1475;
    BITS #(.width(32), .high(31), .low(27)) bits_998 (
        .y(_T_1475),
        .in(io_in)
    );
    wire [31:0] _T_1482_bits;
    wire [4:0] _T_1482_rd;
    wire [4:0] _T_1482_rs1;
    wire [4:0] _T_1482_rs2;
    wire [4:0] _T_1482_rs3;
    wire [4:0] _T_1488;
    BITS #(.width(32), .high(11), .low(7)) bits_999 (
        .y(_T_1488),
        .in(io_in)
    );
    wire [4:0] _T_1489;
    BITS #(.width(32), .high(19), .low(15)) bits_1000 (
        .y(_T_1489),
        .in(io_in)
    );
    wire [4:0] _T_1490;
    BITS #(.width(32), .high(24), .low(20)) bits_1001 (
        .y(_T_1490),
        .in(io_in)
    );
    wire [4:0] _T_1491;
    BITS #(.width(32), .high(31), .low(27)) bits_1002 (
        .y(_T_1491),
        .in(io_in)
    );
    wire [31:0] _T_1498_bits;
    wire [4:0] _T_1498_rd;
    wire [4:0] _T_1498_rs1;
    wire [4:0] _T_1498_rs2;
    wire [4:0] _T_1498_rs3;
    wire [4:0] _T_1504;
    BITS #(.width(32), .high(11), .low(7)) bits_1003 (
        .y(_T_1504),
        .in(io_in)
    );
    wire [4:0] _T_1505;
    BITS #(.width(32), .high(19), .low(15)) bits_1004 (
        .y(_T_1505),
        .in(io_in)
    );
    wire [4:0] _T_1506;
    BITS #(.width(32), .high(24), .low(20)) bits_1005 (
        .y(_T_1506),
        .in(io_in)
    );
    wire [4:0] _T_1507;
    BITS #(.width(32), .high(31), .low(27)) bits_1006 (
        .y(_T_1507),
        .in(io_in)
    );
    wire [31:0] _T_1514_bits;
    wire [4:0] _T_1514_rd;
    wire [4:0] _T_1514_rs1;
    wire [4:0] _T_1514_rs2;
    wire [4:0] _T_1514_rs3;
    wire [4:0] _T_1520;
    BITS #(.width(32), .high(11), .low(7)) bits_1007 (
        .y(_T_1520),
        .in(io_in)
    );
    wire [4:0] _T_1521;
    BITS #(.width(32), .high(19), .low(15)) bits_1008 (
        .y(_T_1521),
        .in(io_in)
    );
    wire [4:0] _T_1522;
    BITS #(.width(32), .high(24), .low(20)) bits_1009 (
        .y(_T_1522),
        .in(io_in)
    );
    wire [4:0] _T_1523;
    BITS #(.width(32), .high(31), .low(27)) bits_1010 (
        .y(_T_1523),
        .in(io_in)
    );
    wire [31:0] _T_1530_bits;
    wire [4:0] _T_1530_rd;
    wire [4:0] _T_1530_rs1;
    wire [4:0] _T_1530_rs2;
    wire [4:0] _T_1530_rs3;
    wire [4:0] _T_1536;
    BITS #(.width(32), .high(11), .low(7)) bits_1011 (
        .y(_T_1536),
        .in(io_in)
    );
    wire [4:0] _T_1537;
    BITS #(.width(32), .high(19), .low(15)) bits_1012 (
        .y(_T_1537),
        .in(io_in)
    );
    wire [4:0] _T_1538;
    BITS #(.width(32), .high(24), .low(20)) bits_1013 (
        .y(_T_1538),
        .in(io_in)
    );
    wire [4:0] _T_1539;
    BITS #(.width(32), .high(31), .low(27)) bits_1014 (
        .y(_T_1539),
        .in(io_in)
    );
    wire [31:0] _T_1546_bits;
    wire [4:0] _T_1546_rd;
    wire [4:0] _T_1546_rs1;
    wire [4:0] _T_1546_rs2;
    wire [4:0] _T_1546_rs3;
    wire [1:0] _T_1552;
    BITS #(.width(32), .high(1), .low(0)) bits_1015 (
        .y(_T_1552),
        .in(io_in)
    );
    wire [2:0] _T_1553;
    BITS #(.width(32), .high(15), .low(13)) bits_1016 (
        .y(_T_1553),
        .in(io_in)
    );
    wire [4:0] _T_1554;
    CAT #(.width_a(2), .width_b(3)) cat_1017 (
        .y(_T_1554),
        .a(_T_1552),
        .b(_T_1553)
    );
    wire [4:0] _T_1556;
    wire [4:0] _WTEMP_61;
    PAD_UNSIGNED #(.width(4), .n(5)) u_pad_1018 (
        .y(_WTEMP_61),
        .in(4'hF)
    );
    BITWISEAND #(.width(5)) bitwiseand_1019 (
        .y(_T_1556),
        .a(_T_1554),
        .b(_WTEMP_61)
    );
    wire _T_1558;
    GEQ_UNSIGNED #(.width(5)) u_geq_1020 (
        .y(_T_1558),
        .a(_T_1554),
        .b(5'h10)
    );
    wire [4:0] _T_1560;
    wire [4:0] _WTEMP_62;
    PAD_UNSIGNED #(.width(3), .n(5)) u_pad_1021 (
        .y(_WTEMP_62),
        .in(3'h7)
    );
    BITWISEAND #(.width(5)) bitwiseand_1022 (
        .y(_T_1560),
        .a(_T_1556),
        .b(_WTEMP_62)
    );
    wire _T_1562;
    wire [4:0] _WTEMP_63;
    PAD_UNSIGNED #(.width(4), .n(5)) u_pad_1023 (
        .y(_WTEMP_63),
        .in(4'h8)
    );
    GEQ_UNSIGNED #(.width(5)) u_geq_1024 (
        .y(_T_1562),
        .a(_T_1556),
        .b(_WTEMP_63)
    );
    wire [4:0] _T_1564;
    wire [4:0] _WTEMP_64;
    PAD_UNSIGNED #(.width(2), .n(5)) u_pad_1025 (
        .y(_WTEMP_64),
        .in(2'h3)
    );
    BITWISEAND #(.width(5)) bitwiseand_1026 (
        .y(_T_1564),
        .a(_T_1560),
        .b(_WTEMP_64)
    );
    wire _T_1566;
    wire [4:0] _WTEMP_65;
    PAD_UNSIGNED #(.width(3), .n(5)) u_pad_1027 (
        .y(_WTEMP_65),
        .in(3'h4)
    );
    GEQ_UNSIGNED #(.width(5)) u_geq_1028 (
        .y(_T_1566),
        .a(_T_1560),
        .b(_WTEMP_65)
    );
    wire [4:0] _T_1568;
    wire [4:0] _WTEMP_66;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_1029 (
        .y(_WTEMP_66),
        .in(1'h1)
    );
    BITWISEAND #(.width(5)) bitwiseand_1030 (
        .y(_T_1568),
        .a(_T_1564),
        .b(_WTEMP_66)
    );
    wire _T_1570;
    wire [4:0] _WTEMP_67;
    PAD_UNSIGNED #(.width(2), .n(5)) u_pad_1031 (
        .y(_WTEMP_67),
        .in(2'h2)
    );
    GEQ_UNSIGNED #(.width(5)) u_geq_1032 (
        .y(_T_1570),
        .a(_T_1564),
        .b(_WTEMP_67)
    );
    wire [4:0] _T_1572;
    assign _T_1572 = 5'h0;
    wire _T_1574;
    wire [4:0] _WTEMP_68;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_1033 (
        .y(_WTEMP_68),
        .in(1'h1)
    );
    GEQ_UNSIGNED #(.width(5)) u_geq_1034 (
        .y(_T_1574),
        .a(_T_1568),
        .b(_WTEMP_68)
    );
    wire [31:0] _T_1575_bits;
    MUX_UNSIGNED #(.width(32)) u_mux_1035 (
        .y(_T_1575_bits),
        .sel(_T_1574),
        .a(_T_1546_bits),
        .b(_T_1530_bits)
    );
    wire [4:0] _T_1575_rd;
    MUX_UNSIGNED #(.width(5)) u_mux_1036 (
        .y(_T_1575_rd),
        .sel(_T_1574),
        .a(_T_1546_rd),
        .b(_T_1530_rd)
    );
    wire [4:0] _T_1575_rs1;
    MUX_UNSIGNED #(.width(5)) u_mux_1037 (
        .y(_T_1575_rs1),
        .sel(_T_1574),
        .a(_T_1546_rs1),
        .b(_T_1530_rs1)
    );
    wire [4:0] _T_1575_rs2;
    MUX_UNSIGNED #(.width(5)) u_mux_1038 (
        .y(_T_1575_rs2),
        .sel(_T_1574),
        .a(_T_1546_rs2),
        .b(_T_1530_rs2)
    );
    wire [4:0] _T_1575_rs3;
    MUX_UNSIGNED #(.width(5)) u_mux_1039 (
        .y(_T_1575_rs3),
        .sel(_T_1574),
        .a(_T_1546_rs3),
        .b(_T_1530_rs3)
    );
    wire [4:0] _T_1582;
    assign _T_1582 = 5'h0;
    wire _T_1584;
    wire [4:0] _WTEMP_69;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_1040 (
        .y(_WTEMP_69),
        .in(1'h1)
    );
    GEQ_UNSIGNED #(.width(5)) u_geq_1041 (
        .y(_T_1584),
        .a(_T_1568),
        .b(_WTEMP_69)
    );
    wire [31:0] _T_1585_bits;
    MUX_UNSIGNED #(.width(32)) u_mux_1042 (
        .y(_T_1585_bits),
        .sel(_T_1584),
        .a(_T_1514_bits),
        .b(_T_1498_bits)
    );
    wire [4:0] _T_1585_rd;
    MUX_UNSIGNED #(.width(5)) u_mux_1043 (
        .y(_T_1585_rd),
        .sel(_T_1584),
        .a(_T_1514_rd),
        .b(_T_1498_rd)
    );
    wire [4:0] _T_1585_rs1;
    MUX_UNSIGNED #(.width(5)) u_mux_1044 (
        .y(_T_1585_rs1),
        .sel(_T_1584),
        .a(_T_1514_rs1),
        .b(_T_1498_rs1)
    );
    wire [4:0] _T_1585_rs2;
    MUX_UNSIGNED #(.width(5)) u_mux_1045 (
        .y(_T_1585_rs2),
        .sel(_T_1584),
        .a(_T_1514_rs2),
        .b(_T_1498_rs2)
    );
    wire [4:0] _T_1585_rs3;
    MUX_UNSIGNED #(.width(5)) u_mux_1046 (
        .y(_T_1585_rs3),
        .sel(_T_1584),
        .a(_T_1514_rs3),
        .b(_T_1498_rs3)
    );
    wire [31:0] _T_1591_bits;
    MUX_UNSIGNED #(.width(32)) u_mux_1047 (
        .y(_T_1591_bits),
        .sel(_T_1570),
        .a(_T_1575_bits),
        .b(_T_1585_bits)
    );
    wire [4:0] _T_1591_rd;
    MUX_UNSIGNED #(.width(5)) u_mux_1048 (
        .y(_T_1591_rd),
        .sel(_T_1570),
        .a(_T_1575_rd),
        .b(_T_1585_rd)
    );
    wire [4:0] _T_1591_rs1;
    MUX_UNSIGNED #(.width(5)) u_mux_1049 (
        .y(_T_1591_rs1),
        .sel(_T_1570),
        .a(_T_1575_rs1),
        .b(_T_1585_rs1)
    );
    wire [4:0] _T_1591_rs2;
    MUX_UNSIGNED #(.width(5)) u_mux_1050 (
        .y(_T_1591_rs2),
        .sel(_T_1570),
        .a(_T_1575_rs2),
        .b(_T_1585_rs2)
    );
    wire [4:0] _T_1591_rs3;
    MUX_UNSIGNED #(.width(5)) u_mux_1051 (
        .y(_T_1591_rs3),
        .sel(_T_1570),
        .a(_T_1575_rs3),
        .b(_T_1585_rs3)
    );
    wire [4:0] _T_1598;
    wire [4:0] _WTEMP_70;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_1052 (
        .y(_WTEMP_70),
        .in(1'h1)
    );
    BITWISEAND #(.width(5)) bitwiseand_1053 (
        .y(_T_1598),
        .a(_T_1564),
        .b(_WTEMP_70)
    );
    wire _T_1600;
    wire [4:0] _WTEMP_71;
    PAD_UNSIGNED #(.width(2), .n(5)) u_pad_1054 (
        .y(_WTEMP_71),
        .in(2'h2)
    );
    GEQ_UNSIGNED #(.width(5)) u_geq_1055 (
        .y(_T_1600),
        .a(_T_1564),
        .b(_WTEMP_71)
    );
    wire [4:0] _T_1602;
    assign _T_1602 = 5'h0;
    wire _T_1604;
    wire [4:0] _WTEMP_72;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_1056 (
        .y(_WTEMP_72),
        .in(1'h1)
    );
    GEQ_UNSIGNED #(.width(5)) u_geq_1057 (
        .y(_T_1604),
        .a(_T_1598),
        .b(_WTEMP_72)
    );
    wire [31:0] _T_1605_bits;
    MUX_UNSIGNED #(.width(32)) u_mux_1058 (
        .y(_T_1605_bits),
        .sel(_T_1604),
        .a(_T_1482_bits),
        .b(_T_1466_bits)
    );
    wire [4:0] _T_1605_rd;
    MUX_UNSIGNED #(.width(5)) u_mux_1059 (
        .y(_T_1605_rd),
        .sel(_T_1604),
        .a(_T_1482_rd),
        .b(_T_1466_rd)
    );
    wire [4:0] _T_1605_rs1;
    MUX_UNSIGNED #(.width(5)) u_mux_1060 (
        .y(_T_1605_rs1),
        .sel(_T_1604),
        .a(_T_1482_rs1),
        .b(_T_1466_rs1)
    );
    wire [4:0] _T_1605_rs2;
    MUX_UNSIGNED #(.width(5)) u_mux_1061 (
        .y(_T_1605_rs2),
        .sel(_T_1604),
        .a(_T_1482_rs2),
        .b(_T_1466_rs2)
    );
    wire [4:0] _T_1605_rs3;
    MUX_UNSIGNED #(.width(5)) u_mux_1062 (
        .y(_T_1605_rs3),
        .sel(_T_1604),
        .a(_T_1482_rs3),
        .b(_T_1466_rs3)
    );
    wire [4:0] _T_1612;
    assign _T_1612 = 5'h0;
    wire _T_1614;
    wire [4:0] _WTEMP_73;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_1063 (
        .y(_WTEMP_73),
        .in(1'h1)
    );
    GEQ_UNSIGNED #(.width(5)) u_geq_1064 (
        .y(_T_1614),
        .a(_T_1598),
        .b(_WTEMP_73)
    );
    wire [31:0] _T_1615_bits;
    MUX_UNSIGNED #(.width(32)) u_mux_1065 (
        .y(_T_1615_bits),
        .sel(_T_1614),
        .a(_T_1450_bits),
        .b(_T_1434_bits)
    );
    wire [4:0] _T_1615_rd;
    MUX_UNSIGNED #(.width(5)) u_mux_1066 (
        .y(_T_1615_rd),
        .sel(_T_1614),
        .a(_T_1450_rd),
        .b(_T_1434_rd)
    );
    wire [4:0] _T_1615_rs1;
    MUX_UNSIGNED #(.width(5)) u_mux_1067 (
        .y(_T_1615_rs1),
        .sel(_T_1614),
        .a(_T_1450_rs1),
        .b(_T_1434_rs1)
    );
    wire [4:0] _T_1615_rs2;
    MUX_UNSIGNED #(.width(5)) u_mux_1068 (
        .y(_T_1615_rs2),
        .sel(_T_1614),
        .a(_T_1450_rs2),
        .b(_T_1434_rs2)
    );
    wire [4:0] _T_1615_rs3;
    MUX_UNSIGNED #(.width(5)) u_mux_1069 (
        .y(_T_1615_rs3),
        .sel(_T_1614),
        .a(_T_1450_rs3),
        .b(_T_1434_rs3)
    );
    wire [31:0] _T_1621_bits;
    MUX_UNSIGNED #(.width(32)) u_mux_1070 (
        .y(_T_1621_bits),
        .sel(_T_1600),
        .a(_T_1605_bits),
        .b(_T_1615_bits)
    );
    wire [4:0] _T_1621_rd;
    MUX_UNSIGNED #(.width(5)) u_mux_1071 (
        .y(_T_1621_rd),
        .sel(_T_1600),
        .a(_T_1605_rd),
        .b(_T_1615_rd)
    );
    wire [4:0] _T_1621_rs1;
    MUX_UNSIGNED #(.width(5)) u_mux_1072 (
        .y(_T_1621_rs1),
        .sel(_T_1600),
        .a(_T_1605_rs1),
        .b(_T_1615_rs1)
    );
    wire [4:0] _T_1621_rs2;
    MUX_UNSIGNED #(.width(5)) u_mux_1073 (
        .y(_T_1621_rs2),
        .sel(_T_1600),
        .a(_T_1605_rs2),
        .b(_T_1615_rs2)
    );
    wire [4:0] _T_1621_rs3;
    MUX_UNSIGNED #(.width(5)) u_mux_1074 (
        .y(_T_1621_rs3),
        .sel(_T_1600),
        .a(_T_1605_rs3),
        .b(_T_1615_rs3)
    );
    wire [31:0] _T_1627_bits;
    MUX_UNSIGNED #(.width(32)) u_mux_1075 (
        .y(_T_1627_bits),
        .sel(_T_1566),
        .a(_T_1591_bits),
        .b(_T_1621_bits)
    );
    wire [4:0] _T_1627_rd;
    MUX_UNSIGNED #(.width(5)) u_mux_1076 (
        .y(_T_1627_rd),
        .sel(_T_1566),
        .a(_T_1591_rd),
        .b(_T_1621_rd)
    );
    wire [4:0] _T_1627_rs1;
    MUX_UNSIGNED #(.width(5)) u_mux_1077 (
        .y(_T_1627_rs1),
        .sel(_T_1566),
        .a(_T_1591_rs1),
        .b(_T_1621_rs1)
    );
    wire [4:0] _T_1627_rs2;
    MUX_UNSIGNED #(.width(5)) u_mux_1078 (
        .y(_T_1627_rs2),
        .sel(_T_1566),
        .a(_T_1591_rs2),
        .b(_T_1621_rs2)
    );
    wire [4:0] _T_1627_rs3;
    MUX_UNSIGNED #(.width(5)) u_mux_1079 (
        .y(_T_1627_rs3),
        .sel(_T_1566),
        .a(_T_1591_rs3),
        .b(_T_1621_rs3)
    );
    wire [4:0] _T_1634;
    wire [4:0] _WTEMP_74;
    PAD_UNSIGNED #(.width(2), .n(5)) u_pad_1080 (
        .y(_WTEMP_74),
        .in(2'h3)
    );
    BITWISEAND #(.width(5)) bitwiseand_1081 (
        .y(_T_1634),
        .a(_T_1560),
        .b(_WTEMP_74)
    );
    wire _T_1636;
    wire [4:0] _WTEMP_75;
    PAD_UNSIGNED #(.width(3), .n(5)) u_pad_1082 (
        .y(_WTEMP_75),
        .in(3'h4)
    );
    GEQ_UNSIGNED #(.width(5)) u_geq_1083 (
        .y(_T_1636),
        .a(_T_1560),
        .b(_WTEMP_75)
    );
    wire [4:0] _T_1638;
    wire [4:0] _WTEMP_76;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_1084 (
        .y(_WTEMP_76),
        .in(1'h1)
    );
    BITWISEAND #(.width(5)) bitwiseand_1085 (
        .y(_T_1638),
        .a(_T_1634),
        .b(_WTEMP_76)
    );
    wire _T_1640;
    wire [4:0] _WTEMP_77;
    PAD_UNSIGNED #(.width(2), .n(5)) u_pad_1086 (
        .y(_WTEMP_77),
        .in(2'h2)
    );
    GEQ_UNSIGNED #(.width(5)) u_geq_1087 (
        .y(_T_1640),
        .a(_T_1634),
        .b(_WTEMP_77)
    );
    wire [4:0] _T_1642;
    assign _T_1642 = 5'h0;
    wire _T_1644;
    wire [4:0] _WTEMP_78;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_1088 (
        .y(_WTEMP_78),
        .in(1'h1)
    );
    GEQ_UNSIGNED #(.width(5)) u_geq_1089 (
        .y(_T_1644),
        .a(_T_1638),
        .b(_WTEMP_78)
    );
    wire [31:0] _T_1645_bits;
    MUX_UNSIGNED #(.width(32)) u_mux_1090 (
        .y(_T_1645_bits),
        .sel(_T_1644),
        .a(_T_1418_bits),
        .b(_T_1381_bits)
    );
    wire [4:0] _T_1645_rd;
    MUX_UNSIGNED #(.width(5)) u_mux_1091 (
        .y(_T_1645_rd),
        .sel(_T_1644),
        .a(_T_1418_rd),
        .b(_T_1381_rd)
    );
    wire [4:0] _T_1645_rs1;
    MUX_UNSIGNED #(.width(5)) u_mux_1092 (
        .y(_T_1645_rs1),
        .sel(_T_1644),
        .a(_T_1418_rs1),
        .b(_T_1381_rs1)
    );
    wire [4:0] _T_1645_rs2;
    MUX_UNSIGNED #(.width(5)) u_mux_1093 (
        .y(_T_1645_rs2),
        .sel(_T_1644),
        .a(_T_1418_rs2),
        .b(_T_1381_rs2)
    );
    wire [4:0] _T_1645_rs3;
    MUX_UNSIGNED #(.width(5)) u_mux_1094 (
        .y(_T_1645_rs3),
        .sel(_T_1644),
        .a(_T_1418_rs3),
        .b(_T_1381_rs3)
    );
    wire [4:0] _T_1652;
    assign _T_1652 = 5'h0;
    wire _T_1654;
    wire [4:0] _WTEMP_79;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_1095 (
        .y(_WTEMP_79),
        .in(1'h1)
    );
    GEQ_UNSIGNED #(.width(5)) u_geq_1096 (
        .y(_T_1654),
        .a(_T_1638),
        .b(_WTEMP_79)
    );
    wire [31:0] _T_1655_bits;
    MUX_UNSIGNED #(.width(32)) u_mux_1097 (
        .y(_T_1655_bits),
        .sel(_T_1654),
        .a(_T_1344_bits),
        .b(_T_1307_bits)
    );
    wire [4:0] _T_1655_rd;
    MUX_UNSIGNED #(.width(5)) u_mux_1098 (
        .y(_T_1655_rd),
        .sel(_T_1654),
        .a(_T_1344_rd),
        .b(_T_1307_rd)
    );
    wire [4:0] _T_1655_rs1;
    MUX_UNSIGNED #(.width(5)) u_mux_1099 (
        .y(_T_1655_rs1),
        .sel(_T_1654),
        .a(_T_1344_rs1),
        .b(_T_1307_rs1)
    );
    wire [4:0] _T_1655_rs2;
    MUX_UNSIGNED #(.width(5)) u_mux_1100 (
        .y(_T_1655_rs2),
        .sel(_T_1654),
        .a(_T_1344_rs2),
        .b(_T_1307_rs2)
    );
    wire [4:0] _T_1655_rs3;
    MUX_UNSIGNED #(.width(5)) u_mux_1101 (
        .y(_T_1655_rs3),
        .sel(_T_1654),
        .a(_T_1344_rs3),
        .b(_T_1307_rs3)
    );
    wire [31:0] _T_1661_bits;
    MUX_UNSIGNED #(.width(32)) u_mux_1102 (
        .y(_T_1661_bits),
        .sel(_T_1640),
        .a(_T_1645_bits),
        .b(_T_1655_bits)
    );
    wire [4:0] _T_1661_rd;
    MUX_UNSIGNED #(.width(5)) u_mux_1103 (
        .y(_T_1661_rd),
        .sel(_T_1640),
        .a(_T_1645_rd),
        .b(_T_1655_rd)
    );
    wire [4:0] _T_1661_rs1;
    MUX_UNSIGNED #(.width(5)) u_mux_1104 (
        .y(_T_1661_rs1),
        .sel(_T_1640),
        .a(_T_1645_rs1),
        .b(_T_1655_rs1)
    );
    wire [4:0] _T_1661_rs2;
    MUX_UNSIGNED #(.width(5)) u_mux_1105 (
        .y(_T_1661_rs2),
        .sel(_T_1640),
        .a(_T_1645_rs2),
        .b(_T_1655_rs2)
    );
    wire [4:0] _T_1661_rs3;
    MUX_UNSIGNED #(.width(5)) u_mux_1106 (
        .y(_T_1661_rs3),
        .sel(_T_1640),
        .a(_T_1645_rs3),
        .b(_T_1655_rs3)
    );
    wire [4:0] _T_1668;
    wire [4:0] _WTEMP_80;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_1107 (
        .y(_WTEMP_80),
        .in(1'h1)
    );
    BITWISEAND #(.width(5)) bitwiseand_1108 (
        .y(_T_1668),
        .a(_T_1634),
        .b(_WTEMP_80)
    );
    wire _T_1670;
    wire [4:0] _WTEMP_81;
    PAD_UNSIGNED #(.width(2), .n(5)) u_pad_1109 (
        .y(_WTEMP_81),
        .in(2'h2)
    );
    GEQ_UNSIGNED #(.width(5)) u_geq_1110 (
        .y(_T_1670),
        .a(_T_1634),
        .b(_WTEMP_81)
    );
    wire [4:0] _T_1672;
    assign _T_1672 = 5'h0;
    wire _T_1674;
    wire [4:0] _WTEMP_82;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_1111 (
        .y(_WTEMP_82),
        .in(1'h1)
    );
    GEQ_UNSIGNED #(.width(5)) u_geq_1112 (
        .y(_T_1674),
        .a(_T_1668),
        .b(_WTEMP_82)
    );
    wire [31:0] _T_1675_bits;
    MUX_UNSIGNED #(.width(32)) u_mux_1113 (
        .y(_T_1675_bits),
        .sel(_T_1674),
        .a(_T_1166_bits),
        .b(_T_1135_bits)
    );
    wire [4:0] _T_1675_rd;
    MUX_UNSIGNED #(.width(5)) u_mux_1114 (
        .y(_T_1675_rd),
        .sel(_T_1674),
        .a(_T_1166_rd),
        .b(_T_1135_rd)
    );
    wire [4:0] _T_1675_rs1;
    MUX_UNSIGNED #(.width(5)) u_mux_1115 (
        .y(_T_1675_rs1),
        .sel(_T_1674),
        .a(_T_1166_rs1),
        .b(_T_1135_rs1)
    );
    wire [4:0] _T_1675_rs2;
    MUX_UNSIGNED #(.width(5)) u_mux_1116 (
        .y(_T_1675_rs2),
        .sel(_T_1674),
        .a(_T_1166_rs2),
        .b(_T_1135_rs2)
    );
    wire [4:0] _T_1675_rs3;
    MUX_UNSIGNED #(.width(5)) u_mux_1117 (
        .y(_T_1675_rs3),
        .sel(_T_1674),
        .a(_T_1166_rs3),
        .b(_T_1135_rs3)
    );
    wire [4:0] _T_1682;
    assign _T_1682 = 5'h0;
    wire _T_1684;
    wire [4:0] _WTEMP_83;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_1118 (
        .y(_WTEMP_83),
        .in(1'h1)
    );
    GEQ_UNSIGNED #(.width(5)) u_geq_1119 (
        .y(_T_1684),
        .a(_T_1668),
        .b(_WTEMP_83)
    );
    wire [31:0] _T_1685_bits;
    MUX_UNSIGNED #(.width(32)) u_mux_1120 (
        .y(_T_1685_bits),
        .sel(_T_1684),
        .a(_T_1104_bits),
        .b(_T_1073_bits)
    );
    wire [4:0] _T_1685_rd;
    MUX_UNSIGNED #(.width(5)) u_mux_1121 (
        .y(_T_1685_rd),
        .sel(_T_1684),
        .a(_T_1104_rd),
        .b(_T_1073_rd)
    );
    wire [4:0] _T_1685_rs1;
    MUX_UNSIGNED #(.width(5)) u_mux_1122 (
        .y(_T_1685_rs1),
        .sel(_T_1684),
        .a(_T_1104_rs1),
        .b(_T_1073_rs1)
    );
    wire [4:0] _T_1685_rs2;
    MUX_UNSIGNED #(.width(5)) u_mux_1123 (
        .y(_T_1685_rs2),
        .sel(_T_1684),
        .a(_T_1104_rs2),
        .b(_T_1073_rs2)
    );
    wire [4:0] _T_1685_rs3;
    MUX_UNSIGNED #(.width(5)) u_mux_1124 (
        .y(_T_1685_rs3),
        .sel(_T_1684),
        .a(_T_1104_rs3),
        .b(_T_1073_rs3)
    );
    wire [31:0] _T_1691_bits;
    MUX_UNSIGNED #(.width(32)) u_mux_1125 (
        .y(_T_1691_bits),
        .sel(_T_1670),
        .a(_T_1675_bits),
        .b(_T_1685_bits)
    );
    wire [4:0] _T_1691_rd;
    MUX_UNSIGNED #(.width(5)) u_mux_1126 (
        .y(_T_1691_rd),
        .sel(_T_1670),
        .a(_T_1675_rd),
        .b(_T_1685_rd)
    );
    wire [4:0] _T_1691_rs1;
    MUX_UNSIGNED #(.width(5)) u_mux_1127 (
        .y(_T_1691_rs1),
        .sel(_T_1670),
        .a(_T_1675_rs1),
        .b(_T_1685_rs1)
    );
    wire [4:0] _T_1691_rs2;
    MUX_UNSIGNED #(.width(5)) u_mux_1128 (
        .y(_T_1691_rs2),
        .sel(_T_1670),
        .a(_T_1675_rs2),
        .b(_T_1685_rs2)
    );
    wire [4:0] _T_1691_rs3;
    MUX_UNSIGNED #(.width(5)) u_mux_1129 (
        .y(_T_1691_rs3),
        .sel(_T_1670),
        .a(_T_1675_rs3),
        .b(_T_1685_rs3)
    );
    wire [31:0] _T_1697_bits;
    MUX_UNSIGNED #(.width(32)) u_mux_1130 (
        .y(_T_1697_bits),
        .sel(_T_1636),
        .a(_T_1661_bits),
        .b(_T_1691_bits)
    );
    wire [4:0] _T_1697_rd;
    MUX_UNSIGNED #(.width(5)) u_mux_1131 (
        .y(_T_1697_rd),
        .sel(_T_1636),
        .a(_T_1661_rd),
        .b(_T_1691_rd)
    );
    wire [4:0] _T_1697_rs1;
    MUX_UNSIGNED #(.width(5)) u_mux_1132 (
        .y(_T_1697_rs1),
        .sel(_T_1636),
        .a(_T_1661_rs1),
        .b(_T_1691_rs1)
    );
    wire [4:0] _T_1697_rs2;
    MUX_UNSIGNED #(.width(5)) u_mux_1133 (
        .y(_T_1697_rs2),
        .sel(_T_1636),
        .a(_T_1661_rs2),
        .b(_T_1691_rs2)
    );
    wire [4:0] _T_1697_rs3;
    MUX_UNSIGNED #(.width(5)) u_mux_1134 (
        .y(_T_1697_rs3),
        .sel(_T_1636),
        .a(_T_1661_rs3),
        .b(_T_1691_rs3)
    );
    wire [31:0] _T_1703_bits;
    MUX_UNSIGNED #(.width(32)) u_mux_1135 (
        .y(_T_1703_bits),
        .sel(_T_1562),
        .a(_T_1627_bits),
        .b(_T_1697_bits)
    );
    wire [4:0] _T_1703_rd;
    MUX_UNSIGNED #(.width(5)) u_mux_1136 (
        .y(_T_1703_rd),
        .sel(_T_1562),
        .a(_T_1627_rd),
        .b(_T_1697_rd)
    );
    wire [4:0] _T_1703_rs1;
    MUX_UNSIGNED #(.width(5)) u_mux_1137 (
        .y(_T_1703_rs1),
        .sel(_T_1562),
        .a(_T_1627_rs1),
        .b(_T_1697_rs1)
    );
    wire [4:0] _T_1703_rs2;
    MUX_UNSIGNED #(.width(5)) u_mux_1138 (
        .y(_T_1703_rs2),
        .sel(_T_1562),
        .a(_T_1627_rs2),
        .b(_T_1697_rs2)
    );
    wire [4:0] _T_1703_rs3;
    MUX_UNSIGNED #(.width(5)) u_mux_1139 (
        .y(_T_1703_rs3),
        .sel(_T_1562),
        .a(_T_1627_rs3),
        .b(_T_1697_rs3)
    );
    wire [4:0] _T_1710;
    wire [4:0] _WTEMP_84;
    PAD_UNSIGNED #(.width(3), .n(5)) u_pad_1140 (
        .y(_WTEMP_84),
        .in(3'h7)
    );
    BITWISEAND #(.width(5)) bitwiseand_1141 (
        .y(_T_1710),
        .a(_T_1556),
        .b(_WTEMP_84)
    );
    wire _T_1712;
    wire [4:0] _WTEMP_85;
    PAD_UNSIGNED #(.width(4), .n(5)) u_pad_1142 (
        .y(_WTEMP_85),
        .in(4'h8)
    );
    GEQ_UNSIGNED #(.width(5)) u_geq_1143 (
        .y(_T_1712),
        .a(_T_1556),
        .b(_WTEMP_85)
    );
    wire [4:0] _T_1714;
    wire [4:0] _WTEMP_86;
    PAD_UNSIGNED #(.width(2), .n(5)) u_pad_1144 (
        .y(_WTEMP_86),
        .in(2'h3)
    );
    BITWISEAND #(.width(5)) bitwiseand_1145 (
        .y(_T_1714),
        .a(_T_1710),
        .b(_WTEMP_86)
    );
    wire _T_1716;
    wire [4:0] _WTEMP_87;
    PAD_UNSIGNED #(.width(3), .n(5)) u_pad_1146 (
        .y(_WTEMP_87),
        .in(3'h4)
    );
    GEQ_UNSIGNED #(.width(5)) u_geq_1147 (
        .y(_T_1716),
        .a(_T_1710),
        .b(_WTEMP_87)
    );
    wire [4:0] _T_1718;
    wire [4:0] _WTEMP_88;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_1148 (
        .y(_WTEMP_88),
        .in(1'h1)
    );
    BITWISEAND #(.width(5)) bitwiseand_1149 (
        .y(_T_1718),
        .a(_T_1714),
        .b(_WTEMP_88)
    );
    wire _T_1720;
    wire [4:0] _WTEMP_89;
    PAD_UNSIGNED #(.width(2), .n(5)) u_pad_1150 (
        .y(_WTEMP_89),
        .in(2'h2)
    );
    GEQ_UNSIGNED #(.width(5)) u_geq_1151 (
        .y(_T_1720),
        .a(_T_1714),
        .b(_WTEMP_89)
    );
    wire [4:0] _T_1722;
    assign _T_1722 = 5'h0;
    wire _T_1724;
    wire [4:0] _WTEMP_90;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_1152 (
        .y(_WTEMP_90),
        .in(1'h1)
    );
    GEQ_UNSIGNED #(.width(5)) u_geq_1153 (
        .y(_T_1724),
        .a(_T_1718),
        .b(_WTEMP_90)
    );
    wire [31:0] _T_1725_bits;
    MUX_UNSIGNED #(.width(32)) u_mux_1154 (
        .y(_T_1725_bits),
        .sel(_T_1724),
        .a(_T_1046_bits),
        .b(_T_951_bits)
    );
    wire [4:0] _T_1725_rd;
    MUX_UNSIGNED #(.width(5)) u_mux_1155 (
        .y(_T_1725_rd),
        .sel(_T_1724),
        .a(_T_1046_rd),
        .b(_T_951_rd)
    );
    wire [4:0] _T_1725_rs1;
    MUX_UNSIGNED #(.width(5)) u_mux_1156 (
        .y(_T_1725_rs1),
        .sel(_T_1724),
        .a(_T_1046_rs1),
        .b(_T_951_rs1)
    );
    wire [4:0] _T_1725_rs2;
    MUX_UNSIGNED #(.width(5)) u_mux_1157 (
        .y(_T_1725_rs2),
        .sel(_T_1724),
        .a(_T_1046_rs2),
        .b(_T_951_rs2)
    );
    wire [4:0] _T_1725_rs3;
    MUX_UNSIGNED #(.width(5)) u_mux_1158 (
        .y(_T_1725_rs3),
        .sel(_T_1724),
        .a(_T_1046_rs3),
        .b(_T_951_rs3)
    );
    wire [4:0] _T_1732;
    assign _T_1732 = 5'h0;
    wire _T_1734;
    wire [4:0] _WTEMP_91;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_1159 (
        .y(_WTEMP_91),
        .in(1'h1)
    );
    GEQ_UNSIGNED #(.width(5)) u_geq_1160 (
        .y(_T_1734),
        .a(_T_1718),
        .b(_WTEMP_91)
    );
    wire [31:0] _T_1735_bits;
    MUX_UNSIGNED #(.width(32)) u_mux_1161 (
        .y(_T_1735_bits),
        .sel(_T_1734),
        .a(_T_854_bits),
        .b(_T_739_bits)
    );
    wire [4:0] _T_1735_rd;
    MUX_UNSIGNED #(.width(5)) u_mux_1162 (
        .y(_T_1735_rd),
        .sel(_T_1734),
        .a(_T_854_rd),
        .b(_T_739_rd)
    );
    wire [4:0] _T_1735_rs1;
    MUX_UNSIGNED #(.width(5)) u_mux_1163 (
        .y(_T_1735_rs1),
        .sel(_T_1734),
        .a(_T_854_rs1),
        .b(_T_739_rs1)
    );
    wire [4:0] _T_1735_rs2;
    MUX_UNSIGNED #(.width(5)) u_mux_1164 (
        .y(_T_1735_rs2),
        .sel(_T_1734),
        .a(_T_854_rs2),
        .b(_T_739_rs2)
    );
    wire [4:0] _T_1735_rs3;
    MUX_UNSIGNED #(.width(5)) u_mux_1165 (
        .y(_T_1735_rs3),
        .sel(_T_1734),
        .a(_T_854_rs3),
        .b(_T_739_rs3)
    );
    wire [31:0] _T_1741_bits;
    MUX_UNSIGNED #(.width(32)) u_mux_1166 (
        .y(_T_1741_bits),
        .sel(_T_1720),
        .a(_T_1725_bits),
        .b(_T_1735_bits)
    );
    wire [4:0] _T_1741_rd;
    MUX_UNSIGNED #(.width(5)) u_mux_1167 (
        .y(_T_1741_rd),
        .sel(_T_1720),
        .a(_T_1725_rd),
        .b(_T_1735_rd)
    );
    wire [4:0] _T_1741_rs1;
    MUX_UNSIGNED #(.width(5)) u_mux_1168 (
        .y(_T_1741_rs1),
        .sel(_T_1720),
        .a(_T_1725_rs1),
        .b(_T_1735_rs1)
    );
    wire [4:0] _T_1741_rs2;
    MUX_UNSIGNED #(.width(5)) u_mux_1169 (
        .y(_T_1741_rs2),
        .sel(_T_1720),
        .a(_T_1725_rs2),
        .b(_T_1735_rs2)
    );
    wire [4:0] _T_1741_rs3;
    MUX_UNSIGNED #(.width(5)) u_mux_1170 (
        .y(_T_1741_rs3),
        .sel(_T_1720),
        .a(_T_1725_rs3),
        .b(_T_1735_rs3)
    );
    wire [4:0] _T_1748;
    wire [4:0] _WTEMP_92;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_1171 (
        .y(_WTEMP_92),
        .in(1'h1)
    );
    BITWISEAND #(.width(5)) bitwiseand_1172 (
        .y(_T_1748),
        .a(_T_1714),
        .b(_WTEMP_92)
    );
    wire _T_1750;
    wire [4:0] _WTEMP_93;
    PAD_UNSIGNED #(.width(2), .n(5)) u_pad_1173 (
        .y(_WTEMP_93),
        .in(2'h2)
    );
    GEQ_UNSIGNED #(.width(5)) u_geq_1174 (
        .y(_T_1750),
        .a(_T_1714),
        .b(_WTEMP_93)
    );
    wire [4:0] _T_1752;
    assign _T_1752 = 5'h0;
    wire _T_1754;
    wire [4:0] _WTEMP_94;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_1175 (
        .y(_WTEMP_94),
        .in(1'h1)
    );
    GEQ_UNSIGNED #(.width(5)) u_geq_1176 (
        .y(_T_1754),
        .a(_T_1748),
        .b(_WTEMP_94)
    );
    wire [31:0] _T_1755_bits;
    MUX_UNSIGNED #(.width(32)) u_mux_1177 (
        .y(_T_1755_bits),
        .sel(_T_1754),
        .a(_T_580_bits),
        .b(_T_472_bits)
    );
    wire [4:0] _T_1755_rd;
    MUX_UNSIGNED #(.width(5)) u_mux_1178 (
        .y(_T_1755_rd),
        .sel(_T_1754),
        .a(_T_580_rd),
        .b(_T_472_rd)
    );
    wire [4:0] _T_1755_rs1;
    MUX_UNSIGNED #(.width(5)) u_mux_1179 (
        .y(_T_1755_rs1),
        .sel(_T_1754),
        .a(_T_580_rs1),
        .b(_T_472_rs1)
    );
    wire [4:0] _T_1755_rs2;
    MUX_UNSIGNED #(.width(5)) u_mux_1180 (
        .y(_T_1755_rs2),
        .sel(_T_1754),
        .a(_T_580_rs2),
        .b(_T_472_rs2)
    );
    wire [4:0] _T_1755_rs3;
    MUX_UNSIGNED #(.width(5)) u_mux_1181 (
        .y(_T_1755_rs3),
        .sel(_T_1754),
        .a(_T_580_rs3),
        .b(_T_472_rs3)
    );
    wire [4:0] _T_1762;
    assign _T_1762 = 5'h0;
    wire _T_1764;
    wire [4:0] _WTEMP_95;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_1182 (
        .y(_WTEMP_95),
        .in(1'h1)
    );
    GEQ_UNSIGNED #(.width(5)) u_geq_1183 (
        .y(_T_1764),
        .a(_T_1748),
        .b(_WTEMP_95)
    );
    wire [31:0] _T_1765_bits;
    MUX_UNSIGNED #(.width(32)) u_mux_1184 (
        .y(_T_1765_bits),
        .sel(_T_1764),
        .a(_T_439_bits),
        .b(_T_401_bits)
    );
    wire [4:0] _T_1765_rd;
    MUX_UNSIGNED #(.width(5)) u_mux_1185 (
        .y(_T_1765_rd),
        .sel(_T_1764),
        .a(_T_439_rd),
        .b(_T_401_rd)
    );
    wire [4:0] _T_1765_rs1;
    MUX_UNSIGNED #(.width(5)) u_mux_1186 (
        .y(_T_1765_rs1),
        .sel(_T_1764),
        .a(_T_439_rs1),
        .b(_T_401_rs1)
    );
    wire [4:0] _T_1765_rs2;
    MUX_UNSIGNED #(.width(5)) u_mux_1187 (
        .y(_T_1765_rs2),
        .sel(_T_1764),
        .a(_T_439_rs2),
        .b(_T_401_rs2)
    );
    wire [4:0] _T_1765_rs3;
    MUX_UNSIGNED #(.width(5)) u_mux_1188 (
        .y(_T_1765_rs3),
        .sel(_T_1764),
        .a(_T_439_rs3),
        .b(_T_401_rs3)
    );
    wire [31:0] _T_1771_bits;
    MUX_UNSIGNED #(.width(32)) u_mux_1189 (
        .y(_T_1771_bits),
        .sel(_T_1750),
        .a(_T_1755_bits),
        .b(_T_1765_bits)
    );
    wire [4:0] _T_1771_rd;
    MUX_UNSIGNED #(.width(5)) u_mux_1190 (
        .y(_T_1771_rd),
        .sel(_T_1750),
        .a(_T_1755_rd),
        .b(_T_1765_rd)
    );
    wire [4:0] _T_1771_rs1;
    MUX_UNSIGNED #(.width(5)) u_mux_1191 (
        .y(_T_1771_rs1),
        .sel(_T_1750),
        .a(_T_1755_rs1),
        .b(_T_1765_rs1)
    );
    wire [4:0] _T_1771_rs2;
    MUX_UNSIGNED #(.width(5)) u_mux_1192 (
        .y(_T_1771_rs2),
        .sel(_T_1750),
        .a(_T_1755_rs2),
        .b(_T_1765_rs2)
    );
    wire [4:0] _T_1771_rs3;
    MUX_UNSIGNED #(.width(5)) u_mux_1193 (
        .y(_T_1771_rs3),
        .sel(_T_1750),
        .a(_T_1755_rs3),
        .b(_T_1765_rs3)
    );
    wire [31:0] _T_1777_bits;
    MUX_UNSIGNED #(.width(32)) u_mux_1194 (
        .y(_T_1777_bits),
        .sel(_T_1716),
        .a(_T_1741_bits),
        .b(_T_1771_bits)
    );
    wire [4:0] _T_1777_rd;
    MUX_UNSIGNED #(.width(5)) u_mux_1195 (
        .y(_T_1777_rd),
        .sel(_T_1716),
        .a(_T_1741_rd),
        .b(_T_1771_rd)
    );
    wire [4:0] _T_1777_rs1;
    MUX_UNSIGNED #(.width(5)) u_mux_1196 (
        .y(_T_1777_rs1),
        .sel(_T_1716),
        .a(_T_1741_rs1),
        .b(_T_1771_rs1)
    );
    wire [4:0] _T_1777_rs2;
    MUX_UNSIGNED #(.width(5)) u_mux_1197 (
        .y(_T_1777_rs2),
        .sel(_T_1716),
        .a(_T_1741_rs2),
        .b(_T_1771_rs2)
    );
    wire [4:0] _T_1777_rs3;
    MUX_UNSIGNED #(.width(5)) u_mux_1198 (
        .y(_T_1777_rs3),
        .sel(_T_1716),
        .a(_T_1741_rs3),
        .b(_T_1771_rs3)
    );
    wire [4:0] _T_1784;
    wire [4:0] _WTEMP_96;
    PAD_UNSIGNED #(.width(2), .n(5)) u_pad_1199 (
        .y(_WTEMP_96),
        .in(2'h3)
    );
    BITWISEAND #(.width(5)) bitwiseand_1200 (
        .y(_T_1784),
        .a(_T_1710),
        .b(_WTEMP_96)
    );
    wire _T_1786;
    wire [4:0] _WTEMP_97;
    PAD_UNSIGNED #(.width(3), .n(5)) u_pad_1201 (
        .y(_WTEMP_97),
        .in(3'h4)
    );
    GEQ_UNSIGNED #(.width(5)) u_geq_1202 (
        .y(_T_1786),
        .a(_T_1710),
        .b(_WTEMP_97)
    );
    wire [4:0] _T_1788;
    wire [4:0] _WTEMP_98;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_1203 (
        .y(_WTEMP_98),
        .in(1'h1)
    );
    BITWISEAND #(.width(5)) bitwiseand_1204 (
        .y(_T_1788),
        .a(_T_1784),
        .b(_WTEMP_98)
    );
    wire _T_1790;
    wire [4:0] _WTEMP_99;
    PAD_UNSIGNED #(.width(2), .n(5)) u_pad_1205 (
        .y(_WTEMP_99),
        .in(2'h2)
    );
    GEQ_UNSIGNED #(.width(5)) u_geq_1206 (
        .y(_T_1790),
        .a(_T_1784),
        .b(_WTEMP_99)
    );
    wire [4:0] _T_1792;
    assign _T_1792 = 5'h0;
    wire _T_1794;
    wire [4:0] _WTEMP_100;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_1207 (
        .y(_WTEMP_100),
        .in(1'h1)
    );
    GEQ_UNSIGNED #(.width(5)) u_geq_1208 (
        .y(_T_1794),
        .a(_T_1788),
        .b(_WTEMP_100)
    );
    wire [31:0] _T_1795_bits;
    MUX_UNSIGNED #(.width(32)) u_mux_1209 (
        .y(_T_1795_bits),
        .sel(_T_1794),
        .a(_T_368_bits),
        .b(_T_321_bits)
    );
    wire [4:0] _T_1795_rd;
    MUX_UNSIGNED #(.width(5)) u_mux_1210 (
        .y(_T_1795_rd),
        .sel(_T_1794),
        .a(_T_368_rd),
        .b(_T_321_rd)
    );
    wire [4:0] _T_1795_rs1;
    MUX_UNSIGNED #(.width(5)) u_mux_1211 (
        .y(_T_1795_rs1),
        .sel(_T_1794),
        .a(_T_368_rs1),
        .b(_T_321_rs1)
    );
    wire [4:0] _T_1795_rs2;
    MUX_UNSIGNED #(.width(5)) u_mux_1212 (
        .y(_T_1795_rs2),
        .sel(_T_1794),
        .a(_T_368_rs2),
        .b(_T_321_rs2)
    );
    wire [4:0] _T_1795_rs3;
    MUX_UNSIGNED #(.width(5)) u_mux_1213 (
        .y(_T_1795_rs3),
        .sel(_T_1794),
        .a(_T_368_rs3),
        .b(_T_321_rs3)
    );
    wire [4:0] _T_1802;
    assign _T_1802 = 5'h0;
    wire _T_1804;
    wire [4:0] _WTEMP_101;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_1214 (
        .y(_WTEMP_101),
        .in(1'h1)
    );
    GEQ_UNSIGNED #(.width(5)) u_geq_1215 (
        .y(_T_1804),
        .a(_T_1788),
        .b(_WTEMP_101)
    );
    wire [31:0] _T_1805_bits;
    MUX_UNSIGNED #(.width(32)) u_mux_1216 (
        .y(_T_1805_bits),
        .sel(_T_1804),
        .a(_T_270_bits),
        .b(_T_223_bits)
    );
    wire [4:0] _T_1805_rd;
    MUX_UNSIGNED #(.width(5)) u_mux_1217 (
        .y(_T_1805_rd),
        .sel(_T_1804),
        .a(_T_270_rd),
        .b(_T_223_rd)
    );
    wire [4:0] _T_1805_rs1;
    MUX_UNSIGNED #(.width(5)) u_mux_1218 (
        .y(_T_1805_rs1),
        .sel(_T_1804),
        .a(_T_270_rs1),
        .b(_T_223_rs1)
    );
    wire [4:0] _T_1805_rs2;
    MUX_UNSIGNED #(.width(5)) u_mux_1219 (
        .y(_T_1805_rs2),
        .sel(_T_1804),
        .a(_T_270_rs2),
        .b(_T_223_rs2)
    );
    wire [4:0] _T_1805_rs3;
    MUX_UNSIGNED #(.width(5)) u_mux_1220 (
        .y(_T_1805_rs3),
        .sel(_T_1804),
        .a(_T_270_rs3),
        .b(_T_223_rs3)
    );
    wire [31:0] _T_1811_bits;
    MUX_UNSIGNED #(.width(32)) u_mux_1221 (
        .y(_T_1811_bits),
        .sel(_T_1790),
        .a(_T_1795_bits),
        .b(_T_1805_bits)
    );
    wire [4:0] _T_1811_rd;
    MUX_UNSIGNED #(.width(5)) u_mux_1222 (
        .y(_T_1811_rd),
        .sel(_T_1790),
        .a(_T_1795_rd),
        .b(_T_1805_rd)
    );
    wire [4:0] _T_1811_rs1;
    MUX_UNSIGNED #(.width(5)) u_mux_1223 (
        .y(_T_1811_rs1),
        .sel(_T_1790),
        .a(_T_1795_rs1),
        .b(_T_1805_rs1)
    );
    wire [4:0] _T_1811_rs2;
    MUX_UNSIGNED #(.width(5)) u_mux_1224 (
        .y(_T_1811_rs2),
        .sel(_T_1790),
        .a(_T_1795_rs2),
        .b(_T_1805_rs2)
    );
    wire [4:0] _T_1811_rs3;
    MUX_UNSIGNED #(.width(5)) u_mux_1225 (
        .y(_T_1811_rs3),
        .sel(_T_1790),
        .a(_T_1795_rs3),
        .b(_T_1805_rs3)
    );
    wire [4:0] _T_1818;
    wire [4:0] _WTEMP_102;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_1226 (
        .y(_WTEMP_102),
        .in(1'h1)
    );
    BITWISEAND #(.width(5)) bitwiseand_1227 (
        .y(_T_1818),
        .a(_T_1784),
        .b(_WTEMP_102)
    );
    wire _T_1820;
    wire [4:0] _WTEMP_103;
    PAD_UNSIGNED #(.width(2), .n(5)) u_pad_1228 (
        .y(_WTEMP_103),
        .in(2'h2)
    );
    GEQ_UNSIGNED #(.width(5)) u_geq_1229 (
        .y(_T_1820),
        .a(_T_1784),
        .b(_WTEMP_103)
    );
    wire [4:0] _T_1822;
    assign _T_1822 = 5'h0;
    wire _T_1824;
    wire [4:0] _WTEMP_104;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_1230 (
        .y(_WTEMP_104),
        .in(1'h1)
    );
    GEQ_UNSIGNED #(.width(5)) u_geq_1231 (
        .y(_T_1824),
        .a(_T_1818),
        .b(_WTEMP_104)
    );
    wire [31:0] _T_1825_bits;
    MUX_UNSIGNED #(.width(32)) u_mux_1232 (
        .y(_T_1825_bits),
        .sel(_T_1824),
        .a(_T_172_bits),
        .b(_T_133_bits)
    );
    wire [4:0] _T_1825_rd;
    MUX_UNSIGNED #(.width(5)) u_mux_1233 (
        .y(_T_1825_rd),
        .sel(_T_1824),
        .a(_T_172_rd),
        .b(_T_133_rd)
    );
    wire [4:0] _T_1825_rs1;
    MUX_UNSIGNED #(.width(5)) u_mux_1234 (
        .y(_T_1825_rs1),
        .sel(_T_1824),
        .a(_T_172_rs1),
        .b(_T_133_rs1)
    );
    wire [4:0] _T_1825_rs2;
    MUX_UNSIGNED #(.width(5)) u_mux_1235 (
        .y(_T_1825_rs2),
        .sel(_T_1824),
        .a(_T_172_rs2),
        .b(_T_133_rs2)
    );
    wire [4:0] _T_1825_rs3;
    MUX_UNSIGNED #(.width(5)) u_mux_1236 (
        .y(_T_1825_rs3),
        .sel(_T_1824),
        .a(_T_172_rs3),
        .b(_T_133_rs3)
    );
    wire [4:0] _T_1832;
    assign _T_1832 = 5'h0;
    wire _T_1834;
    wire [4:0] _WTEMP_105;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_1237 (
        .y(_WTEMP_105),
        .in(1'h1)
    );
    GEQ_UNSIGNED #(.width(5)) u_geq_1238 (
        .y(_T_1834),
        .a(_T_1818),
        .b(_WTEMP_105)
    );
    wire [31:0] _T_1835_bits;
    MUX_UNSIGNED #(.width(32)) u_mux_1239 (
        .y(_T_1835_bits),
        .sel(_T_1834),
        .a(_T_92_bits),
        .b(_T_53_bits)
    );
    wire [4:0] _T_1835_rd;
    MUX_UNSIGNED #(.width(5)) u_mux_1240 (
        .y(_T_1835_rd),
        .sel(_T_1834),
        .a(_T_92_rd),
        .b(_T_53_rd)
    );
    wire [4:0] _T_1835_rs1;
    MUX_UNSIGNED #(.width(5)) u_mux_1241 (
        .y(_T_1835_rs1),
        .sel(_T_1834),
        .a(_T_92_rs1),
        .b(_T_53_rs1)
    );
    wire [4:0] _T_1835_rs2;
    MUX_UNSIGNED #(.width(5)) u_mux_1242 (
        .y(_T_1835_rs2),
        .sel(_T_1834),
        .a(_T_92_rs2),
        .b(_T_53_rs2)
    );
    wire [4:0] _T_1835_rs3;
    MUX_UNSIGNED #(.width(5)) u_mux_1243 (
        .y(_T_1835_rs3),
        .sel(_T_1834),
        .a(_T_92_rs3),
        .b(_T_53_rs3)
    );
    wire [31:0] _T_1841_bits;
    MUX_UNSIGNED #(.width(32)) u_mux_1244 (
        .y(_T_1841_bits),
        .sel(_T_1820),
        .a(_T_1825_bits),
        .b(_T_1835_bits)
    );
    wire [4:0] _T_1841_rd;
    MUX_UNSIGNED #(.width(5)) u_mux_1245 (
        .y(_T_1841_rd),
        .sel(_T_1820),
        .a(_T_1825_rd),
        .b(_T_1835_rd)
    );
    wire [4:0] _T_1841_rs1;
    MUX_UNSIGNED #(.width(5)) u_mux_1246 (
        .y(_T_1841_rs1),
        .sel(_T_1820),
        .a(_T_1825_rs1),
        .b(_T_1835_rs1)
    );
    wire [4:0] _T_1841_rs2;
    MUX_UNSIGNED #(.width(5)) u_mux_1247 (
        .y(_T_1841_rs2),
        .sel(_T_1820),
        .a(_T_1825_rs2),
        .b(_T_1835_rs2)
    );
    wire [4:0] _T_1841_rs3;
    MUX_UNSIGNED #(.width(5)) u_mux_1248 (
        .y(_T_1841_rs3),
        .sel(_T_1820),
        .a(_T_1825_rs3),
        .b(_T_1835_rs3)
    );
    wire [31:0] _T_1847_bits;
    MUX_UNSIGNED #(.width(32)) u_mux_1249 (
        .y(_T_1847_bits),
        .sel(_T_1786),
        .a(_T_1811_bits),
        .b(_T_1841_bits)
    );
    wire [4:0] _T_1847_rd;
    MUX_UNSIGNED #(.width(5)) u_mux_1250 (
        .y(_T_1847_rd),
        .sel(_T_1786),
        .a(_T_1811_rd),
        .b(_T_1841_rd)
    );
    wire [4:0] _T_1847_rs1;
    MUX_UNSIGNED #(.width(5)) u_mux_1251 (
        .y(_T_1847_rs1),
        .sel(_T_1786),
        .a(_T_1811_rs1),
        .b(_T_1841_rs1)
    );
    wire [4:0] _T_1847_rs2;
    MUX_UNSIGNED #(.width(5)) u_mux_1252 (
        .y(_T_1847_rs2),
        .sel(_T_1786),
        .a(_T_1811_rs2),
        .b(_T_1841_rs2)
    );
    wire [4:0] _T_1847_rs3;
    MUX_UNSIGNED #(.width(5)) u_mux_1253 (
        .y(_T_1847_rs3),
        .sel(_T_1786),
        .a(_T_1811_rs3),
        .b(_T_1841_rs3)
    );
    wire [31:0] _T_1853_bits;
    MUX_UNSIGNED #(.width(32)) u_mux_1254 (
        .y(_T_1853_bits),
        .sel(_T_1712),
        .a(_T_1777_bits),
        .b(_T_1847_bits)
    );
    wire [4:0] _T_1853_rd;
    MUX_UNSIGNED #(.width(5)) u_mux_1255 (
        .y(_T_1853_rd),
        .sel(_T_1712),
        .a(_T_1777_rd),
        .b(_T_1847_rd)
    );
    wire [4:0] _T_1853_rs1;
    MUX_UNSIGNED #(.width(5)) u_mux_1256 (
        .y(_T_1853_rs1),
        .sel(_T_1712),
        .a(_T_1777_rs1),
        .b(_T_1847_rs1)
    );
    wire [4:0] _T_1853_rs2;
    MUX_UNSIGNED #(.width(5)) u_mux_1257 (
        .y(_T_1853_rs2),
        .sel(_T_1712),
        .a(_T_1777_rs2),
        .b(_T_1847_rs2)
    );
    wire [4:0] _T_1853_rs3;
    MUX_UNSIGNED #(.width(5)) u_mux_1258 (
        .y(_T_1853_rs3),
        .sel(_T_1712),
        .a(_T_1777_rs3),
        .b(_T_1847_rs3)
    );
    wire [31:0] _T_1859_bits;
    MUX_UNSIGNED #(.width(32)) u_mux_1259 (
        .y(_T_1859_bits),
        .sel(_T_1558),
        .a(_T_1703_bits),
        .b(_T_1853_bits)
    );
    wire [4:0] _T_1859_rd;
    MUX_UNSIGNED #(.width(5)) u_mux_1260 (
        .y(_T_1859_rd),
        .sel(_T_1558),
        .a(_T_1703_rd),
        .b(_T_1853_rd)
    );
    wire [4:0] _T_1859_rs1;
    MUX_UNSIGNED #(.width(5)) u_mux_1261 (
        .y(_T_1859_rs1),
        .sel(_T_1558),
        .a(_T_1703_rs1),
        .b(_T_1853_rs1)
    );
    wire [4:0] _T_1859_rs2;
    MUX_UNSIGNED #(.width(5)) u_mux_1262 (
        .y(_T_1859_rs2),
        .sel(_T_1558),
        .a(_T_1703_rs2),
        .b(_T_1853_rs2)
    );
    wire [4:0] _T_1859_rs3;
    MUX_UNSIGNED #(.width(5)) u_mux_1263 (
        .y(_T_1859_rs3),
        .sel(_T_1558),
        .a(_T_1703_rs3),
        .b(_T_1853_rs3)
    );
    assign _T_1046_bits = _T_1033;
    assign _T_1046_rd = 5'h0;
    assign _T_1046_rs1 = _T_1037;
    assign _T_1046_rs2 = 5'h0;
    assign _T_1046_rs3 = _T_1039;
    PAD_UNSIGNED #(.width(26), .n(32)) u_pad_1264 (
        .y(_T_1073_bits),
        .in(_T_1062)
    );
    assign _T_1073_rd = _T_1063;
    assign _T_1073_rs1 = _T_1064;
    assign _T_1073_rs2 = _T_1065;
    assign _T_1073_rs3 = _T_1066;
    PAD_UNSIGNED #(.width(29), .n(32)) u_pad_1265 (
        .y(_T_1104_bits),
        .in(_T_1093)
    );
    assign _T_1104_rd = _T_1094;
    assign _T_1104_rs1 = 5'h2;
    assign _T_1104_rs2 = _T_1096;
    assign _T_1104_rs3 = _T_1097;
    PAD_UNSIGNED #(.width(28), .n(32)) u_pad_1266 (
        .y(_T_1135_bits),
        .in(_T_1124)
    );
    assign _T_1135_rd = _T_1125;
    assign _T_1135_rs1 = 5'h2;
    assign _T_1135_rs2 = _T_1127;
    assign _T_1135_rs3 = _T_1128;
    PAD_UNSIGNED #(.width(29), .n(32)) u_pad_1267 (
        .y(_T_1166_bits),
        .in(_T_1155)
    );
    assign _T_1166_rd = _T_1156;
    assign _T_1166_rs1 = 5'h2;
    assign _T_1166_rs2 = _T_1158;
    assign _T_1166_rs3 = _T_1159;
    PAD_UNSIGNED #(.width(25), .n(32)) u_pad_1268 (
        .y(_T_1191_bits),
        .in(_T_1180)
    );
    assign _T_1191_rd = _T_1181;
    assign _T_1191_rs1 = 5'h0;
    assign _T_1191_rs2 = _T_1183;
    assign _T_1191_rs3 = _T_1184;
    PAD_UNSIGNED #(.width(25), .n(32)) u_pad_1269 (
        .y(_T_1216_bits),
        .in(_T_1205)
    );
    assign _T_1216_rd = _T_1206;
    assign _T_1216_rs1 = _T_1207;
    assign _T_1216_rs2 = _T_1208;
    assign _T_1216_rs3 = _T_1209;
    PAD_UNSIGNED #(.width(25), .n(32)) u_pad_1270 (
        .y(_T_1248_bits),
        .in(_T_1237)
    );
    assign _T_1248_rd = 5'h0;
    assign _T_1248_rs1 = _T_1239;
    assign _T_1248_rs2 = _T_1240;
    assign _T_1248_rs3 = _T_1241;
    PAD_UNSIGNED #(.width(25), .n(32)) u_pad_1271 (
        .y(_T_1291_bits),
        .in(_T_1280)
    );
    assign _T_1291_rd = 5'h1;
    assign _T_1291_rs1 = _T_1282;
    assign _T_1291_rs2 = _T_1283;
    assign _T_1291_rs3 = _T_1284;
    PAD_UNSIGNED #(.width(27), .n(32)) u_pad_1272 (
        .y(_T_133_bits),
        .in(_T_116)
    );
    assign _T_133_rd = _T_119;
    assign _T_133_rs1 = _T_122;
    assign _T_133_rs2 = _T_125;
    assign _T_133_rs3 = _T_126;
    PAD_UNSIGNED #(.width(29), .n(32)) u_pad_1273 (
        .y(_T_1344_bits),
        .in(_T_1333)
    );
    assign _T_1344_rd = _T_1334;
    assign _T_1344_rs1 = 5'h2;
    assign _T_1344_rs2 = _T_1336;
    assign _T_1344_rs3 = _T_1337;
    PAD_UNSIGNED #(.width(28), .n(32)) u_pad_1274 (
        .y(_T_1381_bits),
        .in(_T_1370)
    );
    assign _T_1381_rd = _T_1371;
    assign _T_1381_rs1 = 5'h2;
    assign _T_1381_rs2 = _T_1373;
    assign _T_1381_rs3 = _T_1374;
    PAD_UNSIGNED #(.width(29), .n(32)) u_pad_1275 (
        .y(_T_1418_bits),
        .in(_T_1407)
    );
    assign _T_1418_rd = _T_1408;
    assign _T_1418_rs1 = 5'h2;
    assign _T_1418_rs2 = _T_1410;
    assign _T_1418_rs3 = _T_1411;
    assign _T_1434_bits = io_in;
    assign _T_1434_rd = _T_1424;
    assign _T_1434_rs1 = _T_1425;
    assign _T_1434_rs2 = _T_1426;
    assign _T_1434_rs3 = _T_1427;
    assign _T_1450_bits = io_in;
    assign _T_1450_rd = _T_1440;
    assign _T_1450_rs1 = _T_1441;
    assign _T_1450_rs2 = _T_1442;
    assign _T_1450_rs3 = _T_1443;
    assign _T_1466_bits = io_in;
    assign _T_1466_rd = _T_1456;
    assign _T_1466_rs1 = _T_1457;
    assign _T_1466_rs2 = _T_1458;
    assign _T_1466_rs3 = _T_1459;
    assign _T_1482_bits = io_in;
    assign _T_1482_rd = _T_1472;
    assign _T_1482_rs1 = _T_1473;
    assign _T_1482_rs2 = _T_1474;
    assign _T_1482_rs3 = _T_1475;
    assign _T_1498_bits = io_in;
    assign _T_1498_rd = _T_1488;
    assign _T_1498_rs1 = _T_1489;
    assign _T_1498_rs2 = _T_1490;
    assign _T_1498_rs3 = _T_1491;
    assign _T_1514_bits = io_in;
    assign _T_1514_rd = _T_1504;
    assign _T_1514_rs1 = _T_1505;
    assign _T_1514_rs2 = _T_1506;
    assign _T_1514_rs3 = _T_1507;
    assign _T_1530_bits = io_in;
    assign _T_1530_rd = _T_1520;
    assign _T_1530_rs1 = _T_1521;
    assign _T_1530_rs2 = _T_1522;
    assign _T_1530_rs3 = _T_1523;
    assign _T_1546_bits = io_in;
    assign _T_1546_rd = _T_1536;
    assign _T_1546_rs1 = _T_1537;
    assign _T_1546_rs2 = _T_1538;
    assign _T_1546_rs3 = _T_1539;
    PAD_UNSIGNED #(.width(28), .n(32)) u_pad_1276 (
        .y(_T_172_bits),
        .in(_T_155)
    );
    assign _T_172_rd = _T_158;
    assign _T_172_rs1 = _T_161;
    assign _T_172_rs2 = _T_164;
    assign _T_172_rs3 = _T_165;
    PAD_UNSIGNED #(.width(27), .n(32)) u_pad_1277 (
        .y(_T_223_bits),
        .in(_T_206)
    );
    assign _T_223_rd = _T_209;
    assign _T_223_rs1 = _T_212;
    assign _T_223_rs2 = _T_215;
    assign _T_223_rs3 = _T_216;
    PAD_UNSIGNED #(.width(28), .n(32)) u_pad_1278 (
        .y(_T_270_bits),
        .in(_T_253)
    );
    assign _T_270_rd = _T_256;
    assign _T_270_rs1 = _T_259;
    assign _T_270_rs2 = _T_262;
    assign _T_270_rs3 = _T_263;
    PAD_UNSIGNED #(.width(27), .n(32)) u_pad_1279 (
        .y(_T_321_bits),
        .in(_T_304)
    );
    assign _T_321_rd = _T_307;
    assign _T_321_rs1 = _T_310;
    assign _T_321_rs2 = _T_313;
    assign _T_321_rs3 = _T_314;
    PAD_UNSIGNED #(.width(28), .n(32)) u_pad_1280 (
        .y(_T_368_bits),
        .in(_T_351)
    );
    assign _T_368_rd = _T_354;
    assign _T_368_rs1 = _T_357;
    assign _T_368_rs2 = _T_360;
    assign _T_368_rs3 = _T_361;
    assign _T_401_bits = _T_388;
    assign _T_401_rd = _T_389;
    assign _T_401_rs1 = _T_390;
    assign _T_401_rs2 = _T_393;
    assign _T_401_rs3 = _T_394;
    assign _T_439_bits = _T_426;
    assign _T_439_rd = _T_427;
    assign _T_439_rs1 = _T_428;
    assign _T_439_rs2 = _T_431;
    assign _T_439_rs3 = _T_432;
    assign _T_472_bits = _T_459;
    assign _T_472_rd = _T_460;
    assign _T_472_rs1 = 5'h0;
    assign _T_472_rs2 = _T_464;
    assign _T_472_rs3 = _T_465;
    assign _T_515_bits = _T_502;
    assign _T_515_rd = _T_503;
    assign _T_515_rs1 = _T_504;
    assign _T_515_rs2 = _T_507;
    assign _T_515_rs3 = _T_508;
    PAD_UNSIGNED #(.width(30), .n(32)) u_pad_1281 (
        .y(_T_53_bits),
        .in(_T_38)
    );
    assign _T_53_rd = _T_41;
    assign _T_53_rs1 = 5'h2;
    assign _T_53_rs2 = _T_45;
    assign _T_53_rs3 = _T_46;
    assign _T_574_bits = _T_561;
    assign _T_574_rd = _T_562;
    assign _T_574_rs1 = _T_563;
    assign _T_574_rs2 = _T_566;
    assign _T_574_rs3 = _T_567;
    assign _T_739_bits = _T_722;
    assign _T_739_rd = _T_725;
    assign _T_739_rs1 = _T_728;
    assign _T_739_rs2 = _T_731;
    assign _T_739_rs3 = _T_732;
    assign _T_854_bits = _T_839;
    assign _T_854_rd = 5'h0;
    assign _T_854_rs1 = _T_843;
    assign _T_854_rs2 = _T_846;
    assign _T_854_rs3 = _T_847;
    PAD_UNSIGNED #(.width(28), .n(32)) u_pad_1282 (
        .y(_T_92_bits),
        .in(_T_75)
    );
    assign _T_92_rd = _T_78;
    assign _T_92_rs1 = _T_81;
    assign _T_92_rs2 = _T_84;
    assign _T_92_rs3 = _T_85;
    assign _T_951_bits = _T_936;
    assign _T_951_rd = _T_939;
    assign _T_951_rs1 = _T_942;
    assign _T_951_rs2 = 5'h0;
    assign _T_951_rs3 = _T_944;
    assign io_out_bits = _T_1859_bits;
    assign io_out_rd = _T_1859_rd;
    assign io_out_rs1 = _T_1859_rs1;
    assign io_out_rs2 = _T_1859_rs2;
    assign io_out_rs3 = _T_1859_rs3;
    assign io_rvc = _T_14;
endmodule //RVCExpander
module MRMWMEM(read_datas, read_clks, read_ens, read_addrs, write_clks, write_ens, write_masks, write_addrs, write_datas);
    parameter depth = 16;
    parameter addrbits = 4;
    parameter width = 32;
    parameter readernum = 2;
    parameter writernum = 2;
    parameter isSyncRead = 0;
    output [(width*readernum-1):0] read_datas;
    input [(1*readernum-1):0] read_clks;
    input [(1*readernum-1):0] read_ens;
    input [(addrbits*readernum-1):0] read_addrs;
    input [1*writernum-1:0] write_clks;
    input [1*writernum-1:0] write_ens;
    input [1*writernum-1:0] write_masks;
    input [(addrbits*writernum-1):0] write_addrs;
    input [(width*writernum-1):0] write_datas;
    reg [width-1:0] memcore [0:depth-1];
    wire [(addrbits*readernum-1):0] final_read_addrs;
    genvar gv_n;
    generate
        for (gv_n = 0; gv_n < readernum; gv_n = gv_n + 1) begin: get_final_raddrs
            if (isSyncRead) begin: raddr_processor
                reg [addrbits-1:0] read_addr_pipe_0;
                always @(posedge read_clks[gv_n]) begin
                    if (read_ens[gv_n]) begin
                        read_addr_pipe_0 <= read_addrs[gv_n*addrbits +: addrbits];
                    end
                end
                assign final_read_addrs[gv_n*addrbits +: addrbits] = read_addr_pipe_0;
            end else begin: raddr_processor
                assign final_read_addrs[gv_n*addrbits +: addrbits] = read_addrs[gv_n*addrbits +: addrbits];
            end
        end
    endgenerate
    genvar gv_k;
    generate
        for (gv_k = 0; gv_k < readernum; gv_k = gv_k + 1) begin: form_read_datas
            assign read_datas[gv_k*width +: width] = memcore[final_read_addrs[gv_k*addrbits +: addrbits]];
        end
    endgenerate
    integer i;
    always @(posedge write_clks[0]) begin
        for (i = 0; i < writernum; i = i + 1) begin
            if (write_ens[i] & write_masks[i]) begin
                memcore[write_addrs[i*addrbits +: addrbits]] <= write_datas[i*width +: width];
            end
        end
    end
endmodule // MRMWMEM
module ASSINT(y, in);
    parameter width = 4;
    output [width-1:0] y;
    input [width-1:0] in;
    assign y = $signed(in);
endmodule // ASSINT
module PAD_SIGNED(y, in);
    parameter width = 4;
    parameter n = 4;
    output [(n > width ? n : width)-1:0] y;
    input [width-1:0] in;
    assign y = n > width ? {{(n - width){in[width-1]}}, in} : in;
endmodule // PAD_SIGNED
module ADD_SIGNED(y, a, b);
    parameter width = 4;
    output [width:0] y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = $signed(a) + $signed(b);
endmodule // ADD_SIGNED
module CSRFile(
    input clock,
    input reset,
    input io_interrupts_debug,
    input io_interrupts_mtip,
    input io_interrupts_msip,
    input io_interrupts_meip,
    input io_interrupts_seip,
    input [63:0] io_hartid,
    input [11:0] io_rw_addr,
    input [2:0] io_rw_cmd,
    output [63:0] io_rw_rdata,
    input [63:0] io_rw_wdata,
    input [11:0] io_decode_csr,
    output io_decode_fp_illegal,
    output io_decode_rocc_illegal,
    output io_decode_read_illegal,
    output io_decode_write_illegal,
    output io_decode_write_flush,
    output io_decode_system_illegal,
    output io_csr_stall,
    output io_eret,
    output io_singleStep,
    output io_status_debug,
    output [31:0] io_status_isa,
    output [1:0] io_status_prv,
    output io_status_sd,
    output [26:0] io_status_zero2,
    output [1:0] io_status_sxl,
    output [1:0] io_status_uxl,
    output io_status_sd_rv32,
    output [7:0] io_status_zero1,
    output io_status_tsr,
    output io_status_tw,
    output io_status_tvm,
    output io_status_mxr,
    output io_status_pum,
    output io_status_mprv,
    output [1:0] io_status_xs,
    output [1:0] io_status_fs,
    output [1:0] io_status_mpp,
    output [1:0] io_status_hpp,
    output io_status_spp,
    output io_status_mpie,
    output io_status_hpie,
    output io_status_spie,
    output io_status_upie,
    output io_status_mie,
    output io_status_hie,
    output io_status_sie,
    output io_status_uie,
    output [3:0] io_ptbr_mode,
    output [15:0] io_ptbr_asid,
    output [43:0] io_ptbr_ppn,
    output [39:0] io_evec,
    input io_exception,
    input io_retire,
    input [63:0] io_cause,
    input [39:0] io_pc,
    input [39:0] io_badaddr,
    output io_fatc,
    output [63:0] io_time,
    output [2:0] io_fcsr_rm,
    input io_fcsr_flags_valid,
    input [4:0] io_fcsr_flags_bits,
    input io_rocc_interrupt,
    output io_interrupt,
    output [63:0] io_interrupt_cause,
    output [3:0] io_bp_0_control_ttype,
    output io_bp_0_control_dmode,
    output [5:0] io_bp_0_control_maskmax,
    output [39:0] io_bp_0_control_reserved,
    output io_bp_0_control_action,
    output io_bp_0_control_chain,
    output [1:0] io_bp_0_control_zero,
    output [1:0] io_bp_0_control_tmatch,
    output io_bp_0_control_m,
    output io_bp_0_control_h,
    output io_bp_0_control_s,
    output io_bp_0_control_u,
    output io_bp_0_control_x,
    output io_bp_0_control_w,
    output io_bp_0_control_r,
    output [38:0] io_bp_0_address
);
    wire _T_347_debug;
    wire [31:0] _T_347_isa;
    wire [1:0] _T_347_prv;
    wire _T_347_sd;
    wire [26:0] _T_347_zero2;
    wire [1:0] _T_347_sxl;
    wire [1:0] _T_347_uxl;
    wire _T_347_sd_rv32;
    wire [7:0] _T_347_zero1;
    wire _T_347_tsr;
    wire _T_347_tw;
    wire _T_347_tvm;
    wire _T_347_mxr;
    wire _T_347_pum;
    wire _T_347_mprv;
    wire [1:0] _T_347_xs;
    wire [1:0] _T_347_fs;
    wire [1:0] _T_347_mpp;
    wire [1:0] _T_347_hpp;
    wire _T_347_spp;
    wire _T_347_mpie;
    wire _T_347_hpie;
    wire _T_347_spie;
    wire _T_347_upie;
    wire _T_347_mie;
    wire _T_347_hie;
    wire _T_347_sie;
    wire _T_347_uie;
    wire [98:0] _T_377;
    wire _T_378;
    BITS #(.width(99), .high(0), .low(0)) bits_1825 (
        .y(_T_378),
        .in(_T_377)
    );
    wire _T_379;
    BITS #(.width(99), .high(1), .low(1)) bits_1826 (
        .y(_T_379),
        .in(_T_377)
    );
    wire _T_380;
    BITS #(.width(99), .high(2), .low(2)) bits_1827 (
        .y(_T_380),
        .in(_T_377)
    );
    wire _T_381;
    BITS #(.width(99), .high(3), .low(3)) bits_1828 (
        .y(_T_381),
        .in(_T_377)
    );
    wire _T_382;
    BITS #(.width(99), .high(4), .low(4)) bits_1829 (
        .y(_T_382),
        .in(_T_377)
    );
    wire _T_383;
    BITS #(.width(99), .high(5), .low(5)) bits_1830 (
        .y(_T_383),
        .in(_T_377)
    );
    wire _T_384;
    BITS #(.width(99), .high(6), .low(6)) bits_1831 (
        .y(_T_384),
        .in(_T_377)
    );
    wire _T_385;
    BITS #(.width(99), .high(7), .low(7)) bits_1832 (
        .y(_T_385),
        .in(_T_377)
    );
    wire _T_386;
    BITS #(.width(99), .high(8), .low(8)) bits_1833 (
        .y(_T_386),
        .in(_T_377)
    );
    wire [1:0] _T_387;
    BITS #(.width(99), .high(10), .low(9)) bits_1834 (
        .y(_T_387),
        .in(_T_377)
    );
    wire [1:0] _T_388;
    BITS #(.width(99), .high(12), .low(11)) bits_1835 (
        .y(_T_388),
        .in(_T_377)
    );
    wire [1:0] _T_389;
    BITS #(.width(99), .high(14), .low(13)) bits_1836 (
        .y(_T_389),
        .in(_T_377)
    );
    wire [1:0] _T_390;
    BITS #(.width(99), .high(16), .low(15)) bits_1837 (
        .y(_T_390),
        .in(_T_377)
    );
    wire _T_391;
    BITS #(.width(99), .high(17), .low(17)) bits_1838 (
        .y(_T_391),
        .in(_T_377)
    );
    wire _T_392;
    BITS #(.width(99), .high(18), .low(18)) bits_1839 (
        .y(_T_392),
        .in(_T_377)
    );
    wire _T_393;
    BITS #(.width(99), .high(19), .low(19)) bits_1840 (
        .y(_T_393),
        .in(_T_377)
    );
    wire _T_394;
    BITS #(.width(99), .high(20), .low(20)) bits_1841 (
        .y(_T_394),
        .in(_T_377)
    );
    wire _T_395;
    BITS #(.width(99), .high(21), .low(21)) bits_1842 (
        .y(_T_395),
        .in(_T_377)
    );
    wire _T_396;
    BITS #(.width(99), .high(22), .low(22)) bits_1843 (
        .y(_T_396),
        .in(_T_377)
    );
    wire [7:0] _T_397;
    BITS #(.width(99), .high(30), .low(23)) bits_1844 (
        .y(_T_397),
        .in(_T_377)
    );
    wire _T_398;
    BITS #(.width(99), .high(31), .low(31)) bits_1845 (
        .y(_T_398),
        .in(_T_377)
    );
    wire [1:0] _T_399;
    BITS #(.width(99), .high(33), .low(32)) bits_1846 (
        .y(_T_399),
        .in(_T_377)
    );
    wire [1:0] _T_400;
    BITS #(.width(99), .high(35), .low(34)) bits_1847 (
        .y(_T_400),
        .in(_T_377)
    );
    wire [26:0] _T_401;
    BITS #(.width(99), .high(62), .low(36)) bits_1848 (
        .y(_T_401),
        .in(_T_377)
    );
    wire _T_402;
    BITS #(.width(99), .high(63), .low(63)) bits_1849 (
        .y(_T_402),
        .in(_T_377)
    );
    wire [1:0] _T_403;
    BITS #(.width(99), .high(65), .low(64)) bits_1850 (
        .y(_T_403),
        .in(_T_377)
    );
    wire [31:0] _T_404;
    BITS #(.width(99), .high(97), .low(66)) bits_1851 (
        .y(_T_404),
        .in(_T_377)
    );
    wire _T_405;
    BITS #(.width(99), .high(98), .low(98)) bits_1852 (
        .y(_T_405),
        .in(_T_377)
    );
    wire [1:0] reset_mstatus_prv;
    wire reset_mstatus_tsr;
    wire reset_mstatus_tw;
    wire reset_mstatus_tvm;
    wire reset_mstatus_mxr;
    wire reset_mstatus_pum;
    wire reset_mstatus_mprv;
    wire [1:0] reset_mstatus_fs;
    wire [1:0] reset_mstatus_mpp;
    wire reset_mstatus_spp;
    wire reset_mstatus_mpie;
    wire reset_mstatus_spie;
    wire reset_mstatus_mie;
    wire reset_mstatus_sie;
    wire [1:0] _reg_mstatus_prv__q;
    wire [1:0] _reg_mstatus_prv__d;
    DFF_POSCLK #(.width(2)) reg_mstatus_prv (
        .q(_reg_mstatus_prv__q),
        .d(_reg_mstatus_prv__d),
        .clk(clock)
    );
    wire [1:0] _WTEMP_118;
    MUX_UNSIGNED #(.width(2)) u_mux_1853 (
        .y(_reg_mstatus_prv__d),
        .sel(reset),
        .a(reset_mstatus_prv),
        .b(_WTEMP_118)
    );
    wire _reg_mstatus_tsr__q;
    wire _reg_mstatus_tsr__d;
    DFF_POSCLK #(.width(1)) reg_mstatus_tsr (
        .q(_reg_mstatus_tsr__q),
        .d(_reg_mstatus_tsr__d),
        .clk(clock)
    );
    wire _WTEMP_119;
    MUX_UNSIGNED #(.width(1)) u_mux_1854 (
        .y(_reg_mstatus_tsr__d),
        .sel(reset),
        .a(reset_mstatus_tsr),
        .b(_WTEMP_119)
    );
    wire _reg_mstatus_tw__q;
    wire _reg_mstatus_tw__d;
    DFF_POSCLK #(.width(1)) reg_mstatus_tw (
        .q(_reg_mstatus_tw__q),
        .d(_reg_mstatus_tw__d),
        .clk(clock)
    );
    wire _WTEMP_120;
    MUX_UNSIGNED #(.width(1)) u_mux_1855 (
        .y(_reg_mstatus_tw__d),
        .sel(reset),
        .a(reset_mstatus_tw),
        .b(_WTEMP_120)
    );
    wire _reg_mstatus_tvm__q;
    wire _reg_mstatus_tvm__d;
    DFF_POSCLK #(.width(1)) reg_mstatus_tvm (
        .q(_reg_mstatus_tvm__q),
        .d(_reg_mstatus_tvm__d),
        .clk(clock)
    );
    wire _WTEMP_121;
    MUX_UNSIGNED #(.width(1)) u_mux_1856 (
        .y(_reg_mstatus_tvm__d),
        .sel(reset),
        .a(reset_mstatus_tvm),
        .b(_WTEMP_121)
    );
    wire _reg_mstatus_mxr__q;
    wire _reg_mstatus_mxr__d;
    DFF_POSCLK #(.width(1)) reg_mstatus_mxr (
        .q(_reg_mstatus_mxr__q),
        .d(_reg_mstatus_mxr__d),
        .clk(clock)
    );
    wire _WTEMP_122;
    MUX_UNSIGNED #(.width(1)) u_mux_1857 (
        .y(_reg_mstatus_mxr__d),
        .sel(reset),
        .a(reset_mstatus_mxr),
        .b(_WTEMP_122)
    );
    wire _reg_mstatus_pum__q;
    wire _reg_mstatus_pum__d;
    DFF_POSCLK #(.width(1)) reg_mstatus_pum (
        .q(_reg_mstatus_pum__q),
        .d(_reg_mstatus_pum__d),
        .clk(clock)
    );
    wire _WTEMP_123;
    MUX_UNSIGNED #(.width(1)) u_mux_1858 (
        .y(_reg_mstatus_pum__d),
        .sel(reset),
        .a(reset_mstatus_pum),
        .b(_WTEMP_123)
    );
    wire _reg_mstatus_mprv__q;
    wire _reg_mstatus_mprv__d;
    DFF_POSCLK #(.width(1)) reg_mstatus_mprv (
        .q(_reg_mstatus_mprv__q),
        .d(_reg_mstatus_mprv__d),
        .clk(clock)
    );
    wire _WTEMP_124;
    MUX_UNSIGNED #(.width(1)) u_mux_1859 (
        .y(_reg_mstatus_mprv__d),
        .sel(reset),
        .a(reset_mstatus_mprv),
        .b(_WTEMP_124)
    );
    wire [1:0] _reg_mstatus_fs__q;
    wire [1:0] _reg_mstatus_fs__d;
    DFF_POSCLK #(.width(2)) reg_mstatus_fs (
        .q(_reg_mstatus_fs__q),
        .d(_reg_mstatus_fs__d),
        .clk(clock)
    );
    wire [1:0] _WTEMP_125;
    MUX_UNSIGNED #(.width(2)) u_mux_1860 (
        .y(_reg_mstatus_fs__d),
        .sel(reset),
        .a(reset_mstatus_fs),
        .b(_WTEMP_125)
    );
    wire [1:0] _reg_mstatus_mpp__q;
    wire [1:0] _reg_mstatus_mpp__d;
    DFF_POSCLK #(.width(2)) reg_mstatus_mpp (
        .q(_reg_mstatus_mpp__q),
        .d(_reg_mstatus_mpp__d),
        .clk(clock)
    );
    wire [1:0] _WTEMP_126;
    MUX_UNSIGNED #(.width(2)) u_mux_1861 (
        .y(_reg_mstatus_mpp__d),
        .sel(reset),
        .a(reset_mstatus_mpp),
        .b(_WTEMP_126)
    );
    wire _reg_mstatus_spp__q;
    wire _reg_mstatus_spp__d;
    DFF_POSCLK #(.width(1)) reg_mstatus_spp (
        .q(_reg_mstatus_spp__q),
        .d(_reg_mstatus_spp__d),
        .clk(clock)
    );
    wire _WTEMP_127;
    MUX_UNSIGNED #(.width(1)) u_mux_1862 (
        .y(_reg_mstatus_spp__d),
        .sel(reset),
        .a(reset_mstatus_spp),
        .b(_WTEMP_127)
    );
    wire _reg_mstatus_mpie__q;
    wire _reg_mstatus_mpie__d;
    DFF_POSCLK #(.width(1)) reg_mstatus_mpie (
        .q(_reg_mstatus_mpie__q),
        .d(_reg_mstatus_mpie__d),
        .clk(clock)
    );
    wire _WTEMP_128;
    MUX_UNSIGNED #(.width(1)) u_mux_1863 (
        .y(_reg_mstatus_mpie__d),
        .sel(reset),
        .a(reset_mstatus_mpie),
        .b(_WTEMP_128)
    );
    wire _reg_mstatus_spie__q;
    wire _reg_mstatus_spie__d;
    DFF_POSCLK #(.width(1)) reg_mstatus_spie (
        .q(_reg_mstatus_spie__q),
        .d(_reg_mstatus_spie__d),
        .clk(clock)
    );
    wire _WTEMP_129;
    MUX_UNSIGNED #(.width(1)) u_mux_1864 (
        .y(_reg_mstatus_spie__d),
        .sel(reset),
        .a(reset_mstatus_spie),
        .b(_WTEMP_129)
    );
    wire _reg_mstatus_mie__q;
    wire _reg_mstatus_mie__d;
    DFF_POSCLK #(.width(1)) reg_mstatus_mie (
        .q(_reg_mstatus_mie__q),
        .d(_reg_mstatus_mie__d),
        .clk(clock)
    );
    wire _WTEMP_130;
    MUX_UNSIGNED #(.width(1)) u_mux_1865 (
        .y(_reg_mstatus_mie__d),
        .sel(reset),
        .a(reset_mstatus_mie),
        .b(_WTEMP_130)
    );
    wire _reg_mstatus_sie__q;
    wire _reg_mstatus_sie__d;
    DFF_POSCLK #(.width(1)) reg_mstatus_sie (
        .q(_reg_mstatus_sie__q),
        .d(_reg_mstatus_sie__d),
        .clk(clock)
    );
    wire _WTEMP_131;
    MUX_UNSIGNED #(.width(1)) u_mux_1866 (
        .y(_reg_mstatus_sie__d),
        .sel(reset),
        .a(reset_mstatus_sie),
        .b(_WTEMP_131)
    );
    wire [1:0] new_prv;
    wire _T_465;
    EQ_UNSIGNED #(.width(2)) u_eq_1867 (
        .y(_T_465),
        .a(new_prv),
        .b(2'h2)
    );
    wire [1:0] _T_467;
    wire [1:0] _WTEMP_132;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_1868 (
        .y(_WTEMP_132),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_1869 (
        .y(_T_467),
        .sel(_T_465),
        .a(_WTEMP_132),
        .b(new_prv)
    );
    wire [1:0] _T_505_xdebugver;
    wire _T_505_ndreset;
    wire _T_505_fullreset;
    wire [11:0] _T_505_zero3;
    wire _T_505_ebreakm;
    wire _T_505_ebreakh;
    wire _T_505_ebreaks;
    wire _T_505_ebreaku;
    wire _T_505_zero2;
    wire _T_505_stopcycle;
    wire _T_505_stoptime;
    wire [2:0] _T_505_cause;
    wire _T_505_debugint;
    wire _T_505_zero1;
    wire _T_505_halt;
    wire _T_505_step;
    wire [1:0] _T_505_prv;
    wire [31:0] _T_524;
    wire [1:0] _T_525;
    BITS #(.width(32), .high(1), .low(0)) bits_1870 (
        .y(_T_525),
        .in(_T_524)
    );
    wire _T_526;
    BITS #(.width(32), .high(2), .low(2)) bits_1871 (
        .y(_T_526),
        .in(_T_524)
    );
    wire _T_527;
    BITS #(.width(32), .high(3), .low(3)) bits_1872 (
        .y(_T_527),
        .in(_T_524)
    );
    wire _T_528;
    BITS #(.width(32), .high(4), .low(4)) bits_1873 (
        .y(_T_528),
        .in(_T_524)
    );
    wire _T_529;
    BITS #(.width(32), .high(5), .low(5)) bits_1874 (
        .y(_T_529),
        .in(_T_524)
    );
    wire [2:0] _T_530;
    BITS #(.width(32), .high(8), .low(6)) bits_1875 (
        .y(_T_530),
        .in(_T_524)
    );
    wire _T_531;
    BITS #(.width(32), .high(9), .low(9)) bits_1876 (
        .y(_T_531),
        .in(_T_524)
    );
    wire _T_532;
    BITS #(.width(32), .high(10), .low(10)) bits_1877 (
        .y(_T_532),
        .in(_T_524)
    );
    wire _T_533;
    BITS #(.width(32), .high(11), .low(11)) bits_1878 (
        .y(_T_533),
        .in(_T_524)
    );
    wire _T_534;
    BITS #(.width(32), .high(12), .low(12)) bits_1879 (
        .y(_T_534),
        .in(_T_524)
    );
    wire _T_535;
    BITS #(.width(32), .high(13), .low(13)) bits_1880 (
        .y(_T_535),
        .in(_T_524)
    );
    wire _T_536;
    BITS #(.width(32), .high(14), .low(14)) bits_1881 (
        .y(_T_536),
        .in(_T_524)
    );
    wire _T_537;
    BITS #(.width(32), .high(15), .low(15)) bits_1882 (
        .y(_T_537),
        .in(_T_524)
    );
    wire [11:0] _T_538;
    BITS #(.width(32), .high(27), .low(16)) bits_1883 (
        .y(_T_538),
        .in(_T_524)
    );
    wire _T_539;
    BITS #(.width(32), .high(28), .low(28)) bits_1884 (
        .y(_T_539),
        .in(_T_524)
    );
    wire _T_540;
    BITS #(.width(32), .high(29), .low(29)) bits_1885 (
        .y(_T_540),
        .in(_T_524)
    );
    wire [1:0] _T_541;
    BITS #(.width(32), .high(31), .low(30)) bits_1886 (
        .y(_T_541),
        .in(_T_524)
    );
    wire reset_dcsr_ebreakm;
    wire reset_dcsr_ebreaks;
    wire reset_dcsr_ebreaku;
    wire [2:0] reset_dcsr_cause;
    wire reset_dcsr_debugint;
    wire reset_dcsr_halt;
    wire reset_dcsr_step;
    wire [1:0] reset_dcsr_prv;
    wire _reg_dcsr_ebreakm__q;
    wire _reg_dcsr_ebreakm__d;
    DFF_POSCLK #(.width(1)) reg_dcsr_ebreakm (
        .q(_reg_dcsr_ebreakm__q),
        .d(_reg_dcsr_ebreakm__d),
        .clk(clock)
    );
    wire _WTEMP_133;
    MUX_UNSIGNED #(.width(1)) u_mux_1887 (
        .y(_reg_dcsr_ebreakm__d),
        .sel(reset),
        .a(reset_dcsr_ebreakm),
        .b(_WTEMP_133)
    );
    wire _reg_dcsr_ebreaks__q;
    wire _reg_dcsr_ebreaks__d;
    DFF_POSCLK #(.width(1)) reg_dcsr_ebreaks (
        .q(_reg_dcsr_ebreaks__q),
        .d(_reg_dcsr_ebreaks__d),
        .clk(clock)
    );
    wire _WTEMP_134;
    MUX_UNSIGNED #(.width(1)) u_mux_1888 (
        .y(_reg_dcsr_ebreaks__d),
        .sel(reset),
        .a(reset_dcsr_ebreaks),
        .b(_WTEMP_134)
    );
    wire _reg_dcsr_ebreaku__q;
    wire _reg_dcsr_ebreaku__d;
    DFF_POSCLK #(.width(1)) reg_dcsr_ebreaku (
        .q(_reg_dcsr_ebreaku__q),
        .d(_reg_dcsr_ebreaku__d),
        .clk(clock)
    );
    wire _WTEMP_135;
    MUX_UNSIGNED #(.width(1)) u_mux_1889 (
        .y(_reg_dcsr_ebreaku__d),
        .sel(reset),
        .a(reset_dcsr_ebreaku),
        .b(_WTEMP_135)
    );
    wire [2:0] _reg_dcsr_cause__q;
    wire [2:0] _reg_dcsr_cause__d;
    DFF_POSCLK #(.width(3)) reg_dcsr_cause (
        .q(_reg_dcsr_cause__q),
        .d(_reg_dcsr_cause__d),
        .clk(clock)
    );
    wire [2:0] _WTEMP_136;
    MUX_UNSIGNED #(.width(3)) u_mux_1890 (
        .y(_reg_dcsr_cause__d),
        .sel(reset),
        .a(reset_dcsr_cause),
        .b(_WTEMP_136)
    );
    wire _reg_dcsr_debugint__q;
    wire _reg_dcsr_debugint__d;
    DFF_POSCLK #(.width(1)) reg_dcsr_debugint (
        .q(_reg_dcsr_debugint__q),
        .d(_reg_dcsr_debugint__d),
        .clk(clock)
    );
    wire _WTEMP_137;
    MUX_UNSIGNED #(.width(1)) u_mux_1891 (
        .y(_reg_dcsr_debugint__d),
        .sel(reset),
        .a(reset_dcsr_debugint),
        .b(_WTEMP_137)
    );
    wire _reg_dcsr_halt__q;
    wire _reg_dcsr_halt__d;
    DFF_POSCLK #(.width(1)) reg_dcsr_halt (
        .q(_reg_dcsr_halt__q),
        .d(_reg_dcsr_halt__d),
        .clk(clock)
    );
    wire _WTEMP_138;
    MUX_UNSIGNED #(.width(1)) u_mux_1892 (
        .y(_reg_dcsr_halt__d),
        .sel(reset),
        .a(reset_dcsr_halt),
        .b(_WTEMP_138)
    );
    wire _reg_dcsr_step__q;
    wire _reg_dcsr_step__d;
    DFF_POSCLK #(.width(1)) reg_dcsr_step (
        .q(_reg_dcsr_step__q),
        .d(_reg_dcsr_step__d),
        .clk(clock)
    );
    wire _WTEMP_139;
    MUX_UNSIGNED #(.width(1)) u_mux_1893 (
        .y(_reg_dcsr_step__d),
        .sel(reset),
        .a(reset_dcsr_step),
        .b(_WTEMP_139)
    );
    wire [1:0] _reg_dcsr_prv__q;
    wire [1:0] _reg_dcsr_prv__d;
    DFF_POSCLK #(.width(2)) reg_dcsr_prv (
        .q(_reg_dcsr_prv__q),
        .d(_reg_dcsr_prv__d),
        .clk(clock)
    );
    wire [1:0] _WTEMP_140;
    MUX_UNSIGNED #(.width(2)) u_mux_1894 (
        .y(_reg_dcsr_prv__d),
        .sel(reset),
        .a(reset_dcsr_prv),
        .b(_WTEMP_140)
    );
    wire _T_607_rocc;
    wire _T_607_meip;
    wire _T_607_heip;
    wire _T_607_seip;
    wire _T_607_ueip;
    wire _T_607_mtip;
    wire _T_607_htip;
    wire _T_607_stip;
    wire _T_607_utip;
    wire _T_607_msip;
    wire _T_607_hsip;
    wire _T_607_ssip;
    wire _T_607_usip;
    wire [12:0] _T_622;
    wire _T_623;
    BITS #(.width(13), .high(0), .low(0)) bits_1895 (
        .y(_T_623),
        .in(_T_622)
    );
    wire _T_624;
    BITS #(.width(13), .high(1), .low(1)) bits_1896 (
        .y(_T_624),
        .in(_T_622)
    );
    wire _T_625;
    BITS #(.width(13), .high(2), .low(2)) bits_1897 (
        .y(_T_625),
        .in(_T_622)
    );
    wire _T_626;
    BITS #(.width(13), .high(3), .low(3)) bits_1898 (
        .y(_T_626),
        .in(_T_622)
    );
    wire _T_627;
    BITS #(.width(13), .high(4), .low(4)) bits_1899 (
        .y(_T_627),
        .in(_T_622)
    );
    wire _T_628;
    BITS #(.width(13), .high(5), .low(5)) bits_1900 (
        .y(_T_628),
        .in(_T_622)
    );
    wire _T_629;
    BITS #(.width(13), .high(6), .low(6)) bits_1901 (
        .y(_T_629),
        .in(_T_622)
    );
    wire _T_630;
    BITS #(.width(13), .high(7), .low(7)) bits_1902 (
        .y(_T_630),
        .in(_T_622)
    );
    wire _T_631;
    BITS #(.width(13), .high(8), .low(8)) bits_1903 (
        .y(_T_631),
        .in(_T_622)
    );
    wire _T_632;
    BITS #(.width(13), .high(9), .low(9)) bits_1904 (
        .y(_T_632),
        .in(_T_622)
    );
    wire _T_633;
    BITS #(.width(13), .high(10), .low(10)) bits_1905 (
        .y(_T_633),
        .in(_T_622)
    );
    wire _T_634;
    BITS #(.width(13), .high(11), .low(11)) bits_1906 (
        .y(_T_634),
        .in(_T_622)
    );
    wire _T_635;
    BITS #(.width(13), .high(12), .low(12)) bits_1907 (
        .y(_T_635),
        .in(_T_622)
    );
    wire _T_636_rocc;
    wire _T_636_meip;
    wire _T_636_heip;
    wire _T_636_seip;
    wire _T_636_ueip;
    wire _T_636_mtip;
    wire _T_636_htip;
    wire _T_636_stip;
    wire _T_636_utip;
    wire _T_636_msip;
    wire _T_636_hsip;
    wire _T_636_ssip;
    wire _T_636_usip;
    wire _T_657_rocc;
    wire _T_657_meip;
    wire _T_657_heip;
    wire _T_657_seip;
    wire _T_657_ueip;
    wire _T_657_mtip;
    wire _T_657_htip;
    wire _T_657_stip;
    wire _T_657_utip;
    wire _T_657_msip;
    wire _T_657_hsip;
    wire _T_657_ssip;
    wire _T_657_usip;
    wire [1:0] _T_674;
    CAT #(.width_a(1), .width_b(1)) cat_1908 (
        .y(_T_674),
        .a(_T_636_hsip),
        .b(_T_636_ssip)
    );
    wire [2:0] _T_675;
    CAT #(.width_a(2), .width_b(1)) cat_1909 (
        .y(_T_675),
        .a(_T_674),
        .b(_T_636_usip)
    );
    wire [1:0] _T_676;
    CAT #(.width_a(1), .width_b(1)) cat_1910 (
        .y(_T_676),
        .a(_T_636_stip),
        .b(_T_636_utip)
    );
    wire [2:0] _T_677;
    CAT #(.width_a(2), .width_b(1)) cat_1911 (
        .y(_T_677),
        .a(_T_676),
        .b(_T_636_msip)
    );
    wire [5:0] _T_678;
    CAT #(.width_a(3), .width_b(3)) cat_1912 (
        .y(_T_678),
        .a(_T_677),
        .b(_T_675)
    );
    wire [1:0] _T_679;
    CAT #(.width_a(1), .width_b(1)) cat_1913 (
        .y(_T_679),
        .a(_T_636_ueip),
        .b(_T_636_mtip)
    );
    wire [2:0] _T_680;
    CAT #(.width_a(2), .width_b(1)) cat_1914 (
        .y(_T_680),
        .a(_T_679),
        .b(_T_636_htip)
    );
    wire [1:0] _T_681;
    CAT #(.width_a(1), .width_b(1)) cat_1915 (
        .y(_T_681),
        .a(_T_636_heip),
        .b(_T_636_seip)
    );
    wire [1:0] _T_682;
    CAT #(.width_a(1), .width_b(1)) cat_1916 (
        .y(_T_682),
        .a(_T_636_rocc),
        .b(_T_636_meip)
    );
    wire [3:0] _T_683;
    CAT #(.width_a(2), .width_b(2)) cat_1917 (
        .y(_T_683),
        .a(_T_682),
        .b(_T_681)
    );
    wire [6:0] _T_684;
    CAT #(.width_a(4), .width_b(3)) cat_1918 (
        .y(_T_684),
        .a(_T_683),
        .b(_T_680)
    );
    wire [12:0] supported_interrupts;
    CAT #(.width_a(7), .width_b(6)) cat_1919 (
        .y(supported_interrupts),
        .a(_T_684),
        .b(_T_678)
    );
    wire [1:0] _T_685;
    CAT #(.width_a(1), .width_b(1)) cat_1920 (
        .y(_T_685),
        .a(_T_657_hsip),
        .b(_T_657_ssip)
    );
    wire [2:0] _T_686;
    CAT #(.width_a(2), .width_b(1)) cat_1921 (
        .y(_T_686),
        .a(_T_685),
        .b(_T_657_usip)
    );
    wire [1:0] _T_687;
    CAT #(.width_a(1), .width_b(1)) cat_1922 (
        .y(_T_687),
        .a(_T_657_stip),
        .b(_T_657_utip)
    );
    wire [2:0] _T_688;
    CAT #(.width_a(2), .width_b(1)) cat_1923 (
        .y(_T_688),
        .a(_T_687),
        .b(_T_657_msip)
    );
    wire [5:0] _T_689;
    CAT #(.width_a(3), .width_b(3)) cat_1924 (
        .y(_T_689),
        .a(_T_688),
        .b(_T_686)
    );
    wire [1:0] _T_690;
    CAT #(.width_a(1), .width_b(1)) cat_1925 (
        .y(_T_690),
        .a(_T_657_ueip),
        .b(_T_657_mtip)
    );
    wire [2:0] _T_691;
    CAT #(.width_a(2), .width_b(1)) cat_1926 (
        .y(_T_691),
        .a(_T_690),
        .b(_T_657_htip)
    );
    wire [1:0] _T_692;
    CAT #(.width_a(1), .width_b(1)) cat_1927 (
        .y(_T_692),
        .a(_T_657_heip),
        .b(_T_657_seip)
    );
    wire [1:0] _T_693;
    CAT #(.width_a(1), .width_b(1)) cat_1928 (
        .y(_T_693),
        .a(_T_657_rocc),
        .b(_T_657_meip)
    );
    wire [3:0] _T_694;
    CAT #(.width_a(2), .width_b(2)) cat_1929 (
        .y(_T_694),
        .a(_T_693),
        .b(_T_692)
    );
    wire [6:0] _T_695;
    CAT #(.width_a(4), .width_b(3)) cat_1930 (
        .y(_T_695),
        .a(_T_694),
        .b(_T_691)
    );
    wire [12:0] delegable_interrupts;
    CAT #(.width_a(7), .width_b(6)) cat_1931 (
        .y(delegable_interrupts),
        .a(_T_695),
        .b(_T_689)
    );
    wire _reg_debug__q;
    wire _reg_debug__d;
    DFF_POSCLK #(.width(1)) reg_debug (
        .q(_reg_debug__q),
        .d(_reg_debug__d),
        .clk(clock)
    );
    wire _WTEMP_141;
    MUX_UNSIGNED #(.width(1)) u_mux_1932 (
        .y(_reg_debug__d),
        .sel(reset),
        .a(1'h0),
        .b(_WTEMP_141)
    );
    wire [2:0] effective_prv;
    CAT #(.width_a(1), .width_b(2)) cat_1933 (
        .y(effective_prv),
        .a(_reg_debug__q),
        .b(_reg_mstatus_prv__q)
    );
    wire [39:0] _reg_dpc__q;
    wire [39:0] _reg_dpc__d;
    DFF_POSCLK #(.width(40)) reg_dpc (
        .q(_reg_dpc__q),
        .d(_reg_dpc__d),
        .clk(clock)
    );
    wire [63:0] _reg_dscratch__q;
    wire [63:0] _reg_dscratch__d;
    DFF_POSCLK #(.width(64)) reg_dscratch (
        .q(_reg_dscratch__q),
        .d(_reg_dscratch__d),
        .clk(clock)
    );
    wire _reg_singleStepped__q;
    wire _reg_singleStepped__d;
    DFF_POSCLK #(.width(1)) reg_singleStepped (
        .q(_reg_singleStepped__q),
        .d(_reg_singleStepped__d),
        .clk(clock)
    );
    wire _reg_bp_0_control_dmode__q;
    wire _reg_bp_0_control_dmode__d;
    DFF_POSCLK #(.width(1)) reg_bp_0_control_dmode (
        .q(_reg_bp_0_control_dmode__q),
        .d(_reg_bp_0_control_dmode__d),
        .clk(clock)
    );
    wire _reg_bp_0_control_action__q;
    wire _reg_bp_0_control_action__d;
    DFF_POSCLK #(.width(1)) reg_bp_0_control_action (
        .q(_reg_bp_0_control_action__q),
        .d(_reg_bp_0_control_action__d),
        .clk(clock)
    );
    wire [1:0] _reg_bp_0_control_tmatch__q;
    wire [1:0] _reg_bp_0_control_tmatch__d;
    DFF_POSCLK #(.width(2)) reg_bp_0_control_tmatch (
        .q(_reg_bp_0_control_tmatch__q),
        .d(_reg_bp_0_control_tmatch__d),
        .clk(clock)
    );
    wire _reg_bp_0_control_m__q;
    wire _reg_bp_0_control_m__d;
    DFF_POSCLK #(.width(1)) reg_bp_0_control_m (
        .q(_reg_bp_0_control_m__q),
        .d(_reg_bp_0_control_m__d),
        .clk(clock)
    );
    wire _reg_bp_0_control_s__q;
    wire _reg_bp_0_control_s__d;
    DFF_POSCLK #(.width(1)) reg_bp_0_control_s (
        .q(_reg_bp_0_control_s__q),
        .d(_reg_bp_0_control_s__d),
        .clk(clock)
    );
    wire _reg_bp_0_control_u__q;
    wire _reg_bp_0_control_u__d;
    DFF_POSCLK #(.width(1)) reg_bp_0_control_u (
        .q(_reg_bp_0_control_u__q),
        .d(_reg_bp_0_control_u__d),
        .clk(clock)
    );
    wire _reg_bp_0_control_x__q;
    wire _reg_bp_0_control_x__d;
    DFF_POSCLK #(.width(1)) reg_bp_0_control_x (
        .q(_reg_bp_0_control_x__q),
        .d(_reg_bp_0_control_x__d),
        .clk(clock)
    );
    wire _reg_bp_0_control_w__q;
    wire _reg_bp_0_control_w__d;
    DFF_POSCLK #(.width(1)) reg_bp_0_control_w (
        .q(_reg_bp_0_control_w__q),
        .d(_reg_bp_0_control_w__d),
        .clk(clock)
    );
    wire _reg_bp_0_control_r__q;
    wire _reg_bp_0_control_r__d;
    DFF_POSCLK #(.width(1)) reg_bp_0_control_r (
        .q(_reg_bp_0_control_r__q),
        .d(_reg_bp_0_control_r__d),
        .clk(clock)
    );
    wire [38:0] _reg_bp_0_address__q;
    wire [38:0] _reg_bp_0_address__d;
    DFF_POSCLK #(.width(39)) reg_bp_0_address (
        .q(_reg_bp_0_address__q),
        .d(_reg_bp_0_address__d),
        .clk(clock)
    );
    wire _reg_bp_1_control_dmode__q;
    wire _reg_bp_1_control_dmode__d;
    DFF_POSCLK #(.width(1)) reg_bp_1_control_dmode (
        .q(_reg_bp_1_control_dmode__q),
        .d(_reg_bp_1_control_dmode__d),
        .clk(clock)
    );
    wire _reg_bp_1_control_action__q;
    wire _reg_bp_1_control_action__d;
    DFF_POSCLK #(.width(1)) reg_bp_1_control_action (
        .q(_reg_bp_1_control_action__q),
        .d(_reg_bp_1_control_action__d),
        .clk(clock)
    );
    wire [1:0] _reg_bp_1_control_tmatch__q;
    wire [1:0] _reg_bp_1_control_tmatch__d;
    DFF_POSCLK #(.width(2)) reg_bp_1_control_tmatch (
        .q(_reg_bp_1_control_tmatch__q),
        .d(_reg_bp_1_control_tmatch__d),
        .clk(clock)
    );
    wire _reg_bp_1_control_m__q;
    wire _reg_bp_1_control_m__d;
    DFF_POSCLK #(.width(1)) reg_bp_1_control_m (
        .q(_reg_bp_1_control_m__q),
        .d(_reg_bp_1_control_m__d),
        .clk(clock)
    );
    wire _reg_bp_1_control_s__q;
    wire _reg_bp_1_control_s__d;
    DFF_POSCLK #(.width(1)) reg_bp_1_control_s (
        .q(_reg_bp_1_control_s__q),
        .d(_reg_bp_1_control_s__d),
        .clk(clock)
    );
    wire _reg_bp_1_control_u__q;
    wire _reg_bp_1_control_u__d;
    DFF_POSCLK #(.width(1)) reg_bp_1_control_u (
        .q(_reg_bp_1_control_u__q),
        .d(_reg_bp_1_control_u__d),
        .clk(clock)
    );
    wire _reg_bp_1_control_x__q;
    wire _reg_bp_1_control_x__d;
    DFF_POSCLK #(.width(1)) reg_bp_1_control_x (
        .q(_reg_bp_1_control_x__q),
        .d(_reg_bp_1_control_x__d),
        .clk(clock)
    );
    wire _reg_bp_1_control_w__q;
    wire _reg_bp_1_control_w__d;
    DFF_POSCLK #(.width(1)) reg_bp_1_control_w (
        .q(_reg_bp_1_control_w__q),
        .d(_reg_bp_1_control_w__d),
        .clk(clock)
    );
    wire _reg_bp_1_control_r__q;
    wire _reg_bp_1_control_r__d;
    DFF_POSCLK #(.width(1)) reg_bp_1_control_r (
        .q(_reg_bp_1_control_r__q),
        .d(_reg_bp_1_control_r__d),
        .clk(clock)
    );
    wire [38:0] _reg_bp_1_address__q;
    wire [38:0] _reg_bp_1_address__d;
    DFF_POSCLK #(.width(39)) reg_bp_1_address (
        .q(_reg_bp_1_address__q),
        .d(_reg_bp_1_address__d),
        .clk(clock)
    );
    wire [63:0] _reg_mie__q;
    wire [63:0] _reg_mie__d;
    DFF_POSCLK #(.width(64)) reg_mie (
        .q(_reg_mie__q),
        .d(_reg_mie__d),
        .clk(clock)
    );
    wire [63:0] _reg_mideleg__q;
    wire [63:0] _reg_mideleg__d;
    DFF_POSCLK #(.width(64)) reg_mideleg (
        .q(_reg_mideleg__q),
        .d(_reg_mideleg__d),
        .clk(clock)
    );
    wire [63:0] _reg_medeleg__q;
    wire [63:0] _reg_medeleg__d;
    DFF_POSCLK #(.width(64)) reg_medeleg (
        .q(_reg_medeleg__q),
        .d(_reg_medeleg__d),
        .clk(clock)
    );
    wire _reg_mip_rocc__q;
    wire _reg_mip_rocc__d;
    DFF_POSCLK #(.width(1)) reg_mip_rocc (
        .q(_reg_mip_rocc__q),
        .d(_reg_mip_rocc__d),
        .clk(clock)
    );
    wire _reg_mip_meip__q;
    wire _reg_mip_meip__d;
    DFF_POSCLK #(.width(1)) reg_mip_meip (
        .q(_reg_mip_meip__q),
        .d(_reg_mip_meip__d),
        .clk(clock)
    );
    wire _reg_mip_heip__q;
    wire _reg_mip_heip__d;
    DFF_POSCLK #(.width(1)) reg_mip_heip (
        .q(_reg_mip_heip__q),
        .d(_reg_mip_heip__d),
        .clk(clock)
    );
    wire _reg_mip_seip__q;
    wire _reg_mip_seip__d;
    DFF_POSCLK #(.width(1)) reg_mip_seip (
        .q(_reg_mip_seip__q),
        .d(_reg_mip_seip__d),
        .clk(clock)
    );
    wire _reg_mip_ueip__q;
    wire _reg_mip_ueip__d;
    DFF_POSCLK #(.width(1)) reg_mip_ueip (
        .q(_reg_mip_ueip__q),
        .d(_reg_mip_ueip__d),
        .clk(clock)
    );
    wire _reg_mip_mtip__q;
    wire _reg_mip_mtip__d;
    DFF_POSCLK #(.width(1)) reg_mip_mtip (
        .q(_reg_mip_mtip__q),
        .d(_reg_mip_mtip__d),
        .clk(clock)
    );
    wire _reg_mip_htip__q;
    wire _reg_mip_htip__d;
    DFF_POSCLK #(.width(1)) reg_mip_htip (
        .q(_reg_mip_htip__q),
        .d(_reg_mip_htip__d),
        .clk(clock)
    );
    wire _reg_mip_stip__q;
    wire _reg_mip_stip__d;
    DFF_POSCLK #(.width(1)) reg_mip_stip (
        .q(_reg_mip_stip__q),
        .d(_reg_mip_stip__d),
        .clk(clock)
    );
    wire _reg_mip_utip__q;
    wire _reg_mip_utip__d;
    DFF_POSCLK #(.width(1)) reg_mip_utip (
        .q(_reg_mip_utip__q),
        .d(_reg_mip_utip__d),
        .clk(clock)
    );
    wire _reg_mip_msip__q;
    wire _reg_mip_msip__d;
    DFF_POSCLK #(.width(1)) reg_mip_msip (
        .q(_reg_mip_msip__q),
        .d(_reg_mip_msip__d),
        .clk(clock)
    );
    wire _reg_mip_hsip__q;
    wire _reg_mip_hsip__d;
    DFF_POSCLK #(.width(1)) reg_mip_hsip (
        .q(_reg_mip_hsip__q),
        .d(_reg_mip_hsip__d),
        .clk(clock)
    );
    wire _reg_mip_ssip__q;
    wire _reg_mip_ssip__d;
    DFF_POSCLK #(.width(1)) reg_mip_ssip (
        .q(_reg_mip_ssip__q),
        .d(_reg_mip_ssip__d),
        .clk(clock)
    );
    wire _reg_mip_usip__q;
    wire _reg_mip_usip__d;
    DFF_POSCLK #(.width(1)) reg_mip_usip (
        .q(_reg_mip_usip__q),
        .d(_reg_mip_usip__d),
        .clk(clock)
    );
    wire [39:0] _reg_mepc__q;
    wire [39:0] _reg_mepc__d;
    DFF_POSCLK #(.width(40)) reg_mepc (
        .q(_reg_mepc__q),
        .d(_reg_mepc__d),
        .clk(clock)
    );
    wire [63:0] _reg_mcause__q;
    wire [63:0] _reg_mcause__d;
    DFF_POSCLK #(.width(64)) reg_mcause (
        .q(_reg_mcause__q),
        .d(_reg_mcause__d),
        .clk(clock)
    );
    wire [39:0] _reg_mbadaddr__q;
    wire [39:0] _reg_mbadaddr__d;
    DFF_POSCLK #(.width(40)) reg_mbadaddr (
        .q(_reg_mbadaddr__q),
        .d(_reg_mbadaddr__d),
        .clk(clock)
    );
    wire [63:0] _reg_mscratch__q;
    wire [63:0] _reg_mscratch__d;
    DFF_POSCLK #(.width(64)) reg_mscratch (
        .q(_reg_mscratch__q),
        .d(_reg_mscratch__d),
        .clk(clock)
    );
    wire [31:0] _reg_mtvec__q;
    wire [31:0] _reg_mtvec__d;
    DFF_POSCLK #(.width(32)) reg_mtvec (
        .q(_reg_mtvec__q),
        .d(_reg_mtvec__d),
        .clk(clock)
    );
    wire [31:0] _WTEMP_142;
    MUX_UNSIGNED #(.width(32)) u_mux_1934 (
        .y(_reg_mtvec__d),
        .sel(reset),
        .a(32'h0),
        .b(_WTEMP_142)
    );
    wire [31:0] _reg_mcounteren__q;
    wire [31:0] _reg_mcounteren__d;
    DFF_POSCLK #(.width(32)) reg_mcounteren (
        .q(_reg_mcounteren__q),
        .d(_reg_mcounteren__d),
        .clk(clock)
    );
    wire [31:0] _reg_scounteren__q;
    wire [31:0] _reg_scounteren__d;
    DFF_POSCLK #(.width(32)) reg_scounteren (
        .q(_reg_scounteren__q),
        .d(_reg_scounteren__d),
        .clk(clock)
    );
    wire [39:0] _reg_sepc__q;
    wire [39:0] _reg_sepc__d;
    DFF_POSCLK #(.width(40)) reg_sepc (
        .q(_reg_sepc__q),
        .d(_reg_sepc__d),
        .clk(clock)
    );
    wire [63:0] _reg_scause__q;
    wire [63:0] _reg_scause__d;
    DFF_POSCLK #(.width(64)) reg_scause (
        .q(_reg_scause__q),
        .d(_reg_scause__d),
        .clk(clock)
    );
    wire [39:0] _reg_sbadaddr__q;
    wire [39:0] _reg_sbadaddr__d;
    DFF_POSCLK #(.width(40)) reg_sbadaddr (
        .q(_reg_sbadaddr__q),
        .d(_reg_sbadaddr__d),
        .clk(clock)
    );
    wire [63:0] _reg_sscratch__q;
    wire [63:0] _reg_sscratch__d;
    DFF_POSCLK #(.width(64)) reg_sscratch (
        .q(_reg_sscratch__q),
        .d(_reg_sscratch__d),
        .clk(clock)
    );
    wire [38:0] _reg_stvec__q;
    wire [38:0] _reg_stvec__d;
    DFF_POSCLK #(.width(39)) reg_stvec (
        .q(_reg_stvec__q),
        .d(_reg_stvec__d),
        .clk(clock)
    );
    wire [3:0] _reg_sptbr_mode__q;
    wire [3:0] _reg_sptbr_mode__d;
    DFF_POSCLK #(.width(4)) reg_sptbr_mode (
        .q(_reg_sptbr_mode__q),
        .d(_reg_sptbr_mode__d),
        .clk(clock)
    );
    wire [43:0] _reg_sptbr_ppn__q;
    wire [43:0] _reg_sptbr_ppn__d;
    DFF_POSCLK #(.width(44)) reg_sptbr_ppn (
        .q(_reg_sptbr_ppn__q),
        .d(_reg_sptbr_ppn__d),
        .clk(clock)
    );
    wire _reg_wfi__q;
    wire _reg_wfi__d;
    DFF_POSCLK #(.width(1)) reg_wfi (
        .q(_reg_wfi__q),
        .d(_reg_wfi__d),
        .clk(clock)
    );
    wire _WTEMP_143;
    MUX_UNSIGNED #(.width(1)) u_mux_1935 (
        .y(_reg_wfi__d),
        .sel(reset),
        .a(1'h0),
        .b(_WTEMP_143)
    );
    wire [4:0] _reg_fflags__q;
    wire [4:0] _reg_fflags__d;
    DFF_POSCLK #(.width(5)) reg_fflags (
        .q(_reg_fflags__q),
        .d(_reg_fflags__d),
        .clk(clock)
    );
    wire [2:0] _reg_frm__q;
    wire [2:0] _reg_frm__d;
    DFF_POSCLK #(.width(3)) reg_frm (
        .q(_reg_frm__q),
        .d(_reg_frm__d),
        .clk(clock)
    );
    wire [5:0] __T_931__q;
    wire [5:0] __T_931__d;
    DFF_POSCLK #(.width(6)) _T_931 (
        .q(__T_931__q),
        .d(__T_931__d),
        .clk(clock)
    );
    wire [5:0] _WTEMP_144;
    MUX_UNSIGNED #(.width(6)) u_mux_1936 (
        .y(__T_931__d),
        .sel(reset),
        .a(6'h0),
        .b(_WTEMP_144)
    );
    wire [6:0] _T_932;
    wire [5:0] _WTEMP_145;
    PAD_UNSIGNED #(.width(1), .n(6)) u_pad_1937 (
        .y(_WTEMP_145),
        .in(io_retire)
    );
    ADD_UNSIGNED #(.width(6)) u_add_1938 (
        .y(_T_932),
        .a(__T_931__q),
        .b(_WTEMP_145)
    );
    wire [57:0] __T_934__q;
    wire [57:0] __T_934__d;
    DFF_POSCLK #(.width(58)) _T_934 (
        .q(__T_934__q),
        .d(__T_934__d),
        .clk(clock)
    );
    wire [57:0] _WTEMP_146;
    MUX_UNSIGNED #(.width(58)) u_mux_1939 (
        .y(__T_934__d),
        .sel(reset),
        .a(58'h0),
        .b(_WTEMP_146)
    );
    wire _T_935;
    BITS #(.width(7), .high(6), .low(6)) bits_1940 (
        .y(_T_935),
        .in(_T_932)
    );
    wire [58:0] _T_937;
    wire [57:0] _WTEMP_147;
    PAD_UNSIGNED #(.width(1), .n(58)) u_pad_1941 (
        .y(_WTEMP_147),
        .in(1'h1)
    );
    ADD_UNSIGNED #(.width(58)) u_add_1942 (
        .y(_T_937),
        .a(__T_934__q),
        .b(_WTEMP_147)
    );
    wire [57:0] _T_938;
    TAIL #(.width(59), .n(1)) tail_1943 (
        .y(_T_938),
        .in(_T_937)
    );
    wire [63:0] _T_939;
    CAT #(.width_a(58), .width_b(6)) cat_1944 (
        .y(_T_939),
        .a(__T_934__q),
        .b(__T_931__q)
    );
    wire [5:0] __T_942__q;
    wire [5:0] __T_942__d;
    DFF_POSCLK #(.width(6)) _T_942 (
        .q(__T_942__q),
        .d(__T_942__d),
        .clk(clock)
    );
    wire [5:0] _WTEMP_148;
    MUX_UNSIGNED #(.width(6)) u_mux_1945 (
        .y(__T_942__d),
        .sel(reset),
        .a(6'h0),
        .b(_WTEMP_148)
    );
    wire [6:0] _T_943;
    wire [5:0] _WTEMP_149;
    PAD_UNSIGNED #(.width(1), .n(6)) u_pad_1946 (
        .y(_WTEMP_149),
        .in(1'h1)
    );
    ADD_UNSIGNED #(.width(6)) u_add_1947 (
        .y(_T_943),
        .a(__T_942__q),
        .b(_WTEMP_149)
    );
    wire [57:0] __T_945__q;
    wire [57:0] __T_945__d;
    DFF_POSCLK #(.width(58)) _T_945 (
        .q(__T_945__q),
        .d(__T_945__d),
        .clk(clock)
    );
    wire [57:0] _WTEMP_150;
    MUX_UNSIGNED #(.width(58)) u_mux_1948 (
        .y(__T_945__d),
        .sel(reset),
        .a(58'h0),
        .b(_WTEMP_150)
    );
    wire _T_946;
    BITS #(.width(7), .high(6), .low(6)) bits_1949 (
        .y(_T_946),
        .in(_T_943)
    );
    wire [58:0] _T_948;
    wire [57:0] _WTEMP_151;
    PAD_UNSIGNED #(.width(1), .n(58)) u_pad_1950 (
        .y(_WTEMP_151),
        .in(1'h1)
    );
    ADD_UNSIGNED #(.width(58)) u_add_1951 (
        .y(_T_948),
        .a(__T_945__q),
        .b(_WTEMP_151)
    );
    wire [57:0] _T_949;
    TAIL #(.width(59), .n(1)) tail_1952 (
        .y(_T_949),
        .in(_T_948)
    );
    wire [63:0] _T_950;
    CAT #(.width_a(58), .width_b(6)) cat_1953 (
        .y(_T_950),
        .a(__T_945__q),
        .b(__T_942__q)
    );
    wire _T_953;
    wire [1:0] _WTEMP_152;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_1954 (
        .y(_WTEMP_152),
        .in(1'h1)
    );
    EQ_UNSIGNED #(.width(2)) u_eq_1955 (
        .y(_T_953),
        .a(_reg_mstatus_prv__q),
        .b(_WTEMP_152)
    );
    wire _T_954;
    BITWISEOR #(.width(1)) bitwiseor_1956 (
        .y(_T_954),
        .a(1'h0),
        .b(_T_953)
    );
    wire [31:0] _T_956;
    wire [31:0] _WTEMP_153;
    PAD_UNSIGNED #(.width(3), .n(32)) u_pad_1957 (
        .y(_WTEMP_153),
        .in(3'h7)
    );
    MUX_UNSIGNED #(.width(32)) u_mux_1958 (
        .y(_T_956),
        .sel(_T_954),
        .a(_WTEMP_153),
        .b(_reg_scounteren__q)
    );
    wire [31:0] hpm_mask;
    BITWISEAND #(.width(32)) bitwiseand_1959 (
        .y(hpm_mask),
        .a(_reg_mcounteren__q),
        .b(_T_956)
    );
    wire mip_rocc;
    wire mip_meip;
    wire mip_heip;
    wire mip_seip;
    wire mip_ueip;
    wire mip_mtip;
    wire mip_htip;
    wire mip_stip;
    wire mip_utip;
    wire mip_msip;
    wire mip_hsip;
    wire mip_ssip;
    wire mip_usip;
    wire [1:0] _T_970;
    CAT #(.width_a(1), .width_b(1)) cat_1960 (
        .y(_T_970),
        .a(mip_hsip),
        .b(mip_ssip)
    );
    wire [2:0] _T_971;
    CAT #(.width_a(2), .width_b(1)) cat_1961 (
        .y(_T_971),
        .a(_T_970),
        .b(mip_usip)
    );
    wire [1:0] _T_972;
    CAT #(.width_a(1), .width_b(1)) cat_1962 (
        .y(_T_972),
        .a(mip_stip),
        .b(mip_utip)
    );
    wire [2:0] _T_973;
    CAT #(.width_a(2), .width_b(1)) cat_1963 (
        .y(_T_973),
        .a(_T_972),
        .b(mip_msip)
    );
    wire [5:0] _T_974;
    CAT #(.width_a(3), .width_b(3)) cat_1964 (
        .y(_T_974),
        .a(_T_973),
        .b(_T_971)
    );
    wire [1:0] _T_975;
    CAT #(.width_a(1), .width_b(1)) cat_1965 (
        .y(_T_975),
        .a(mip_ueip),
        .b(mip_mtip)
    );
    wire [2:0] _T_976;
    CAT #(.width_a(2), .width_b(1)) cat_1966 (
        .y(_T_976),
        .a(_T_975),
        .b(mip_htip)
    );
    wire [1:0] _T_977;
    CAT #(.width_a(1), .width_b(1)) cat_1967 (
        .y(_T_977),
        .a(mip_heip),
        .b(mip_seip)
    );
    wire [1:0] _T_978;
    CAT #(.width_a(1), .width_b(1)) cat_1968 (
        .y(_T_978),
        .a(mip_rocc),
        .b(mip_meip)
    );
    wire [3:0] _T_979;
    CAT #(.width_a(2), .width_b(2)) cat_1969 (
        .y(_T_979),
        .a(_T_978),
        .b(_T_977)
    );
    wire [6:0] _T_980;
    CAT #(.width_a(4), .width_b(3)) cat_1970 (
        .y(_T_980),
        .a(_T_979),
        .b(_T_976)
    );
    wire [12:0] _T_981;
    CAT #(.width_a(7), .width_b(6)) cat_1971 (
        .y(_T_981),
        .a(_T_980),
        .b(_T_974)
    );
    wire [12:0] read_mip;
    BITWISEAND #(.width(13)) bitwiseand_1972 (
        .y(read_mip),
        .a(_T_981),
        .b(supported_interrupts)
    );
    wire [63:0] pending_interrupts;
    wire [63:0] _WTEMP_154;
    PAD_UNSIGNED #(.width(13), .n(64)) u_pad_1973 (
        .y(_WTEMP_154),
        .in(read_mip)
    );
    BITWISEAND #(.width(64)) bitwiseand_1974 (
        .y(pending_interrupts),
        .a(_WTEMP_154),
        .b(_reg_mie__q)
    );
    wire _T_983;
    wire [1:0] _WTEMP_155;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_1975 (
        .y(_WTEMP_155),
        .in(1'h1)
    );
    LEQ_UNSIGNED #(.width(2)) u_leq_1976 (
        .y(_T_983),
        .a(_reg_mstatus_prv__q),
        .b(_WTEMP_155)
    );
    wire _T_985;
    EQ_UNSIGNED #(.width(2)) u_eq_1977 (
        .y(_T_985),
        .a(_reg_mstatus_prv__q),
        .b(2'h3)
    );
    wire _T_986;
    BITWISEAND #(.width(1)) bitwiseand_1978 (
        .y(_T_986),
        .a(_T_985),
        .b(_reg_mstatus_mie__q)
    );
    wire _T_987;
    BITWISEOR #(.width(1)) bitwiseor_1979 (
        .y(_T_987),
        .a(_T_983),
        .b(_T_986)
    );
    wire [63:0] _T_988;
    BITWISENOT #(.width(64)) bitwisenot_1980 (
        .y(_T_988),
        .in(_reg_mideleg__q)
    );
    wire [63:0] _T_989;
    BITWISEAND #(.width(64)) bitwiseand_1981 (
        .y(_T_989),
        .a(pending_interrupts),
        .b(_T_988)
    );
    wire [63:0] m_interrupts;
    wire [63:0] _WTEMP_156;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_1982 (
        .y(_WTEMP_156),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_1983 (
        .y(m_interrupts),
        .sel(_T_987),
        .a(_T_989),
        .b(_WTEMP_156)
    );
    wire _T_992;
    wire [63:0] _WTEMP_157;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_1984 (
        .y(_WTEMP_157),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(64)) u_eq_1985 (
        .y(_T_992),
        .a(m_interrupts),
        .b(_WTEMP_157)
    );
    wire _T_994;
    wire [1:0] _WTEMP_158;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_1986 (
        .y(_WTEMP_158),
        .in(1'h1)
    );
    LT_UNSIGNED #(.width(2)) u_lt_1987 (
        .y(_T_994),
        .a(_reg_mstatus_prv__q),
        .b(_WTEMP_158)
    );
    wire _T_996;
    wire [1:0] _WTEMP_159;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_1988 (
        .y(_WTEMP_159),
        .in(1'h1)
    );
    EQ_UNSIGNED #(.width(2)) u_eq_1989 (
        .y(_T_996),
        .a(_reg_mstatus_prv__q),
        .b(_WTEMP_159)
    );
    wire _T_997;
    BITWISEAND #(.width(1)) bitwiseand_1990 (
        .y(_T_997),
        .a(_T_996),
        .b(_reg_mstatus_sie__q)
    );
    wire _T_998;
    BITWISEOR #(.width(1)) bitwiseor_1991 (
        .y(_T_998),
        .a(_T_994),
        .b(_T_997)
    );
    wire _T_999;
    BITWISEAND #(.width(1)) bitwiseand_1992 (
        .y(_T_999),
        .a(_T_992),
        .b(_T_998)
    );
    wire [63:0] _T_1000;
    BITWISEAND #(.width(64)) bitwiseand_1993 (
        .y(_T_1000),
        .a(pending_interrupts),
        .b(_reg_mideleg__q)
    );
    wire [63:0] s_interrupts;
    wire [63:0] _WTEMP_160;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_1994 (
        .y(_WTEMP_160),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_1995 (
        .y(s_interrupts),
        .sel(_T_999),
        .a(_T_1000),
        .b(_WTEMP_160)
    );
    wire [63:0] all_interrupts;
    BITWISEOR #(.width(64)) bitwiseor_1996 (
        .y(all_interrupts),
        .a(m_interrupts),
        .b(s_interrupts)
    );
    wire _T_1003;
    BITS #(.width(64), .high(0), .low(0)) bits_1997 (
        .y(_T_1003),
        .in(all_interrupts)
    );
    wire _T_1004;
    BITS #(.width(64), .high(1), .low(1)) bits_1998 (
        .y(_T_1004),
        .in(all_interrupts)
    );
    wire _T_1005;
    BITS #(.width(64), .high(2), .low(2)) bits_1999 (
        .y(_T_1005),
        .in(all_interrupts)
    );
    wire _T_1006;
    BITS #(.width(64), .high(3), .low(3)) bits_2000 (
        .y(_T_1006),
        .in(all_interrupts)
    );
    wire _T_1007;
    BITS #(.width(64), .high(4), .low(4)) bits_2001 (
        .y(_T_1007),
        .in(all_interrupts)
    );
    wire _T_1008;
    BITS #(.width(64), .high(5), .low(5)) bits_2002 (
        .y(_T_1008),
        .in(all_interrupts)
    );
    wire _T_1009;
    BITS #(.width(64), .high(6), .low(6)) bits_2003 (
        .y(_T_1009),
        .in(all_interrupts)
    );
    wire _T_1010;
    BITS #(.width(64), .high(7), .low(7)) bits_2004 (
        .y(_T_1010),
        .in(all_interrupts)
    );
    wire _T_1011;
    BITS #(.width(64), .high(8), .low(8)) bits_2005 (
        .y(_T_1011),
        .in(all_interrupts)
    );
    wire _T_1012;
    BITS #(.width(64), .high(9), .low(9)) bits_2006 (
        .y(_T_1012),
        .in(all_interrupts)
    );
    wire _T_1013;
    BITS #(.width(64), .high(10), .low(10)) bits_2007 (
        .y(_T_1013),
        .in(all_interrupts)
    );
    wire _T_1014;
    BITS #(.width(64), .high(11), .low(11)) bits_2008 (
        .y(_T_1014),
        .in(all_interrupts)
    );
    wire _T_1015;
    BITS #(.width(64), .high(12), .low(12)) bits_2009 (
        .y(_T_1015),
        .in(all_interrupts)
    );
    wire _T_1016;
    BITS #(.width(64), .high(13), .low(13)) bits_2010 (
        .y(_T_1016),
        .in(all_interrupts)
    );
    wire _T_1017;
    BITS #(.width(64), .high(14), .low(14)) bits_2011 (
        .y(_T_1017),
        .in(all_interrupts)
    );
    wire _T_1018;
    BITS #(.width(64), .high(15), .low(15)) bits_2012 (
        .y(_T_1018),
        .in(all_interrupts)
    );
    wire _T_1019;
    BITS #(.width(64), .high(16), .low(16)) bits_2013 (
        .y(_T_1019),
        .in(all_interrupts)
    );
    wire _T_1020;
    BITS #(.width(64), .high(17), .low(17)) bits_2014 (
        .y(_T_1020),
        .in(all_interrupts)
    );
    wire _T_1021;
    BITS #(.width(64), .high(18), .low(18)) bits_2015 (
        .y(_T_1021),
        .in(all_interrupts)
    );
    wire _T_1022;
    BITS #(.width(64), .high(19), .low(19)) bits_2016 (
        .y(_T_1022),
        .in(all_interrupts)
    );
    wire _T_1023;
    BITS #(.width(64), .high(20), .low(20)) bits_2017 (
        .y(_T_1023),
        .in(all_interrupts)
    );
    wire _T_1024;
    BITS #(.width(64), .high(21), .low(21)) bits_2018 (
        .y(_T_1024),
        .in(all_interrupts)
    );
    wire _T_1025;
    BITS #(.width(64), .high(22), .low(22)) bits_2019 (
        .y(_T_1025),
        .in(all_interrupts)
    );
    wire _T_1026;
    BITS #(.width(64), .high(23), .low(23)) bits_2020 (
        .y(_T_1026),
        .in(all_interrupts)
    );
    wire _T_1027;
    BITS #(.width(64), .high(24), .low(24)) bits_2021 (
        .y(_T_1027),
        .in(all_interrupts)
    );
    wire _T_1028;
    BITS #(.width(64), .high(25), .low(25)) bits_2022 (
        .y(_T_1028),
        .in(all_interrupts)
    );
    wire _T_1029;
    BITS #(.width(64), .high(26), .low(26)) bits_2023 (
        .y(_T_1029),
        .in(all_interrupts)
    );
    wire _T_1030;
    BITS #(.width(64), .high(27), .low(27)) bits_2024 (
        .y(_T_1030),
        .in(all_interrupts)
    );
    wire _T_1031;
    BITS #(.width(64), .high(28), .low(28)) bits_2025 (
        .y(_T_1031),
        .in(all_interrupts)
    );
    wire _T_1032;
    BITS #(.width(64), .high(29), .low(29)) bits_2026 (
        .y(_T_1032),
        .in(all_interrupts)
    );
    wire _T_1033;
    BITS #(.width(64), .high(30), .low(30)) bits_2027 (
        .y(_T_1033),
        .in(all_interrupts)
    );
    wire _T_1034;
    BITS #(.width(64), .high(31), .low(31)) bits_2028 (
        .y(_T_1034),
        .in(all_interrupts)
    );
    wire _T_1035;
    BITS #(.width(64), .high(32), .low(32)) bits_2029 (
        .y(_T_1035),
        .in(all_interrupts)
    );
    wire _T_1036;
    BITS #(.width(64), .high(33), .low(33)) bits_2030 (
        .y(_T_1036),
        .in(all_interrupts)
    );
    wire _T_1037;
    BITS #(.width(64), .high(34), .low(34)) bits_2031 (
        .y(_T_1037),
        .in(all_interrupts)
    );
    wire _T_1038;
    BITS #(.width(64), .high(35), .low(35)) bits_2032 (
        .y(_T_1038),
        .in(all_interrupts)
    );
    wire _T_1039;
    BITS #(.width(64), .high(36), .low(36)) bits_2033 (
        .y(_T_1039),
        .in(all_interrupts)
    );
    wire _T_1040;
    BITS #(.width(64), .high(37), .low(37)) bits_2034 (
        .y(_T_1040),
        .in(all_interrupts)
    );
    wire _T_1041;
    BITS #(.width(64), .high(38), .low(38)) bits_2035 (
        .y(_T_1041),
        .in(all_interrupts)
    );
    wire _T_1042;
    BITS #(.width(64), .high(39), .low(39)) bits_2036 (
        .y(_T_1042),
        .in(all_interrupts)
    );
    wire _T_1043;
    BITS #(.width(64), .high(40), .low(40)) bits_2037 (
        .y(_T_1043),
        .in(all_interrupts)
    );
    wire _T_1044;
    BITS #(.width(64), .high(41), .low(41)) bits_2038 (
        .y(_T_1044),
        .in(all_interrupts)
    );
    wire _T_1045;
    BITS #(.width(64), .high(42), .low(42)) bits_2039 (
        .y(_T_1045),
        .in(all_interrupts)
    );
    wire _T_1046;
    BITS #(.width(64), .high(43), .low(43)) bits_2040 (
        .y(_T_1046),
        .in(all_interrupts)
    );
    wire _T_1047;
    BITS #(.width(64), .high(44), .low(44)) bits_2041 (
        .y(_T_1047),
        .in(all_interrupts)
    );
    wire _T_1048;
    BITS #(.width(64), .high(45), .low(45)) bits_2042 (
        .y(_T_1048),
        .in(all_interrupts)
    );
    wire _T_1049;
    BITS #(.width(64), .high(46), .low(46)) bits_2043 (
        .y(_T_1049),
        .in(all_interrupts)
    );
    wire _T_1050;
    BITS #(.width(64), .high(47), .low(47)) bits_2044 (
        .y(_T_1050),
        .in(all_interrupts)
    );
    wire _T_1051;
    BITS #(.width(64), .high(48), .low(48)) bits_2045 (
        .y(_T_1051),
        .in(all_interrupts)
    );
    wire _T_1052;
    BITS #(.width(64), .high(49), .low(49)) bits_2046 (
        .y(_T_1052),
        .in(all_interrupts)
    );
    wire _T_1053;
    BITS #(.width(64), .high(50), .low(50)) bits_2047 (
        .y(_T_1053),
        .in(all_interrupts)
    );
    wire _T_1054;
    BITS #(.width(64), .high(51), .low(51)) bits_2048 (
        .y(_T_1054),
        .in(all_interrupts)
    );
    wire _T_1055;
    BITS #(.width(64), .high(52), .low(52)) bits_2049 (
        .y(_T_1055),
        .in(all_interrupts)
    );
    wire _T_1056;
    BITS #(.width(64), .high(53), .low(53)) bits_2050 (
        .y(_T_1056),
        .in(all_interrupts)
    );
    wire _T_1057;
    BITS #(.width(64), .high(54), .low(54)) bits_2051 (
        .y(_T_1057),
        .in(all_interrupts)
    );
    wire _T_1058;
    BITS #(.width(64), .high(55), .low(55)) bits_2052 (
        .y(_T_1058),
        .in(all_interrupts)
    );
    wire _T_1059;
    BITS #(.width(64), .high(56), .low(56)) bits_2053 (
        .y(_T_1059),
        .in(all_interrupts)
    );
    wire _T_1060;
    BITS #(.width(64), .high(57), .low(57)) bits_2054 (
        .y(_T_1060),
        .in(all_interrupts)
    );
    wire _T_1061;
    BITS #(.width(64), .high(58), .low(58)) bits_2055 (
        .y(_T_1061),
        .in(all_interrupts)
    );
    wire _T_1062;
    BITS #(.width(64), .high(59), .low(59)) bits_2056 (
        .y(_T_1062),
        .in(all_interrupts)
    );
    wire _T_1063;
    BITS #(.width(64), .high(60), .low(60)) bits_2057 (
        .y(_T_1063),
        .in(all_interrupts)
    );
    wire _T_1064;
    BITS #(.width(64), .high(61), .low(61)) bits_2058 (
        .y(_T_1064),
        .in(all_interrupts)
    );
    wire _T_1065;
    BITS #(.width(64), .high(62), .low(62)) bits_2059 (
        .y(_T_1065),
        .in(all_interrupts)
    );
    wire _T_1066;
    BITS #(.width(64), .high(63), .low(63)) bits_2060 (
        .y(_T_1066),
        .in(all_interrupts)
    );
    wire [5:0] _T_1131;
    MUX_UNSIGNED #(.width(6)) u_mux_2061 (
        .y(_T_1131),
        .sel(_T_1065),
        .a(6'h3E),
        .b(6'h3F)
    );
    wire [5:0] _T_1132;
    MUX_UNSIGNED #(.width(6)) u_mux_2062 (
        .y(_T_1132),
        .sel(_T_1064),
        .a(6'h3D),
        .b(_T_1131)
    );
    wire [5:0] _T_1133;
    MUX_UNSIGNED #(.width(6)) u_mux_2063 (
        .y(_T_1133),
        .sel(_T_1063),
        .a(6'h3C),
        .b(_T_1132)
    );
    wire [5:0] _T_1134;
    MUX_UNSIGNED #(.width(6)) u_mux_2064 (
        .y(_T_1134),
        .sel(_T_1062),
        .a(6'h3B),
        .b(_T_1133)
    );
    wire [5:0] _T_1135;
    MUX_UNSIGNED #(.width(6)) u_mux_2065 (
        .y(_T_1135),
        .sel(_T_1061),
        .a(6'h3A),
        .b(_T_1134)
    );
    wire [5:0] _T_1136;
    MUX_UNSIGNED #(.width(6)) u_mux_2066 (
        .y(_T_1136),
        .sel(_T_1060),
        .a(6'h39),
        .b(_T_1135)
    );
    wire [5:0] _T_1137;
    MUX_UNSIGNED #(.width(6)) u_mux_2067 (
        .y(_T_1137),
        .sel(_T_1059),
        .a(6'h38),
        .b(_T_1136)
    );
    wire [5:0] _T_1138;
    MUX_UNSIGNED #(.width(6)) u_mux_2068 (
        .y(_T_1138),
        .sel(_T_1058),
        .a(6'h37),
        .b(_T_1137)
    );
    wire [5:0] _T_1139;
    MUX_UNSIGNED #(.width(6)) u_mux_2069 (
        .y(_T_1139),
        .sel(_T_1057),
        .a(6'h36),
        .b(_T_1138)
    );
    wire [5:0] _T_1140;
    MUX_UNSIGNED #(.width(6)) u_mux_2070 (
        .y(_T_1140),
        .sel(_T_1056),
        .a(6'h35),
        .b(_T_1139)
    );
    wire [5:0] _T_1141;
    MUX_UNSIGNED #(.width(6)) u_mux_2071 (
        .y(_T_1141),
        .sel(_T_1055),
        .a(6'h34),
        .b(_T_1140)
    );
    wire [5:0] _T_1142;
    MUX_UNSIGNED #(.width(6)) u_mux_2072 (
        .y(_T_1142),
        .sel(_T_1054),
        .a(6'h33),
        .b(_T_1141)
    );
    wire [5:0] _T_1143;
    MUX_UNSIGNED #(.width(6)) u_mux_2073 (
        .y(_T_1143),
        .sel(_T_1053),
        .a(6'h32),
        .b(_T_1142)
    );
    wire [5:0] _T_1144;
    MUX_UNSIGNED #(.width(6)) u_mux_2074 (
        .y(_T_1144),
        .sel(_T_1052),
        .a(6'h31),
        .b(_T_1143)
    );
    wire [5:0] _T_1145;
    MUX_UNSIGNED #(.width(6)) u_mux_2075 (
        .y(_T_1145),
        .sel(_T_1051),
        .a(6'h30),
        .b(_T_1144)
    );
    wire [5:0] _T_1146;
    MUX_UNSIGNED #(.width(6)) u_mux_2076 (
        .y(_T_1146),
        .sel(_T_1050),
        .a(6'h2F),
        .b(_T_1145)
    );
    wire [5:0] _T_1147;
    MUX_UNSIGNED #(.width(6)) u_mux_2077 (
        .y(_T_1147),
        .sel(_T_1049),
        .a(6'h2E),
        .b(_T_1146)
    );
    wire [5:0] _T_1148;
    MUX_UNSIGNED #(.width(6)) u_mux_2078 (
        .y(_T_1148),
        .sel(_T_1048),
        .a(6'h2D),
        .b(_T_1147)
    );
    wire [5:0] _T_1149;
    MUX_UNSIGNED #(.width(6)) u_mux_2079 (
        .y(_T_1149),
        .sel(_T_1047),
        .a(6'h2C),
        .b(_T_1148)
    );
    wire [5:0] _T_1150;
    MUX_UNSIGNED #(.width(6)) u_mux_2080 (
        .y(_T_1150),
        .sel(_T_1046),
        .a(6'h2B),
        .b(_T_1149)
    );
    wire [5:0] _T_1151;
    MUX_UNSIGNED #(.width(6)) u_mux_2081 (
        .y(_T_1151),
        .sel(_T_1045),
        .a(6'h2A),
        .b(_T_1150)
    );
    wire [5:0] _T_1152;
    MUX_UNSIGNED #(.width(6)) u_mux_2082 (
        .y(_T_1152),
        .sel(_T_1044),
        .a(6'h29),
        .b(_T_1151)
    );
    wire [5:0] _T_1153;
    MUX_UNSIGNED #(.width(6)) u_mux_2083 (
        .y(_T_1153),
        .sel(_T_1043),
        .a(6'h28),
        .b(_T_1152)
    );
    wire [5:0] _T_1154;
    MUX_UNSIGNED #(.width(6)) u_mux_2084 (
        .y(_T_1154),
        .sel(_T_1042),
        .a(6'h27),
        .b(_T_1153)
    );
    wire [5:0] _T_1155;
    MUX_UNSIGNED #(.width(6)) u_mux_2085 (
        .y(_T_1155),
        .sel(_T_1041),
        .a(6'h26),
        .b(_T_1154)
    );
    wire [5:0] _T_1156;
    MUX_UNSIGNED #(.width(6)) u_mux_2086 (
        .y(_T_1156),
        .sel(_T_1040),
        .a(6'h25),
        .b(_T_1155)
    );
    wire [5:0] _T_1157;
    MUX_UNSIGNED #(.width(6)) u_mux_2087 (
        .y(_T_1157),
        .sel(_T_1039),
        .a(6'h24),
        .b(_T_1156)
    );
    wire [5:0] _T_1158;
    MUX_UNSIGNED #(.width(6)) u_mux_2088 (
        .y(_T_1158),
        .sel(_T_1038),
        .a(6'h23),
        .b(_T_1157)
    );
    wire [5:0] _T_1159;
    MUX_UNSIGNED #(.width(6)) u_mux_2089 (
        .y(_T_1159),
        .sel(_T_1037),
        .a(6'h22),
        .b(_T_1158)
    );
    wire [5:0] _T_1160;
    MUX_UNSIGNED #(.width(6)) u_mux_2090 (
        .y(_T_1160),
        .sel(_T_1036),
        .a(6'h21),
        .b(_T_1159)
    );
    wire [5:0] _T_1161;
    MUX_UNSIGNED #(.width(6)) u_mux_2091 (
        .y(_T_1161),
        .sel(_T_1035),
        .a(6'h20),
        .b(_T_1160)
    );
    wire [5:0] _T_1162;
    wire [5:0] _WTEMP_161;
    PAD_UNSIGNED #(.width(5), .n(6)) u_pad_2092 (
        .y(_WTEMP_161),
        .in(5'h1F)
    );
    MUX_UNSIGNED #(.width(6)) u_mux_2093 (
        .y(_T_1162),
        .sel(_T_1034),
        .a(_WTEMP_161),
        .b(_T_1161)
    );
    wire [5:0] _T_1163;
    wire [5:0] _WTEMP_162;
    PAD_UNSIGNED #(.width(5), .n(6)) u_pad_2094 (
        .y(_WTEMP_162),
        .in(5'h1E)
    );
    MUX_UNSIGNED #(.width(6)) u_mux_2095 (
        .y(_T_1163),
        .sel(_T_1033),
        .a(_WTEMP_162),
        .b(_T_1162)
    );
    wire [5:0] _T_1164;
    wire [5:0] _WTEMP_163;
    PAD_UNSIGNED #(.width(5), .n(6)) u_pad_2096 (
        .y(_WTEMP_163),
        .in(5'h1D)
    );
    MUX_UNSIGNED #(.width(6)) u_mux_2097 (
        .y(_T_1164),
        .sel(_T_1032),
        .a(_WTEMP_163),
        .b(_T_1163)
    );
    wire [5:0] _T_1165;
    wire [5:0] _WTEMP_164;
    PAD_UNSIGNED #(.width(5), .n(6)) u_pad_2098 (
        .y(_WTEMP_164),
        .in(5'h1C)
    );
    MUX_UNSIGNED #(.width(6)) u_mux_2099 (
        .y(_T_1165),
        .sel(_T_1031),
        .a(_WTEMP_164),
        .b(_T_1164)
    );
    wire [5:0] _T_1166;
    wire [5:0] _WTEMP_165;
    PAD_UNSIGNED #(.width(5), .n(6)) u_pad_2100 (
        .y(_WTEMP_165),
        .in(5'h1B)
    );
    MUX_UNSIGNED #(.width(6)) u_mux_2101 (
        .y(_T_1166),
        .sel(_T_1030),
        .a(_WTEMP_165),
        .b(_T_1165)
    );
    wire [5:0] _T_1167;
    wire [5:0] _WTEMP_166;
    PAD_UNSIGNED #(.width(5), .n(6)) u_pad_2102 (
        .y(_WTEMP_166),
        .in(5'h1A)
    );
    MUX_UNSIGNED #(.width(6)) u_mux_2103 (
        .y(_T_1167),
        .sel(_T_1029),
        .a(_WTEMP_166),
        .b(_T_1166)
    );
    wire [5:0] _T_1168;
    wire [5:0] _WTEMP_167;
    PAD_UNSIGNED #(.width(5), .n(6)) u_pad_2104 (
        .y(_WTEMP_167),
        .in(5'h19)
    );
    MUX_UNSIGNED #(.width(6)) u_mux_2105 (
        .y(_T_1168),
        .sel(_T_1028),
        .a(_WTEMP_167),
        .b(_T_1167)
    );
    wire [5:0] _T_1169;
    wire [5:0] _WTEMP_168;
    PAD_UNSIGNED #(.width(5), .n(6)) u_pad_2106 (
        .y(_WTEMP_168),
        .in(5'h18)
    );
    MUX_UNSIGNED #(.width(6)) u_mux_2107 (
        .y(_T_1169),
        .sel(_T_1027),
        .a(_WTEMP_168),
        .b(_T_1168)
    );
    wire [5:0] _T_1170;
    wire [5:0] _WTEMP_169;
    PAD_UNSIGNED #(.width(5), .n(6)) u_pad_2108 (
        .y(_WTEMP_169),
        .in(5'h17)
    );
    MUX_UNSIGNED #(.width(6)) u_mux_2109 (
        .y(_T_1170),
        .sel(_T_1026),
        .a(_WTEMP_169),
        .b(_T_1169)
    );
    wire [5:0] _T_1171;
    wire [5:0] _WTEMP_170;
    PAD_UNSIGNED #(.width(5), .n(6)) u_pad_2110 (
        .y(_WTEMP_170),
        .in(5'h16)
    );
    MUX_UNSIGNED #(.width(6)) u_mux_2111 (
        .y(_T_1171),
        .sel(_T_1025),
        .a(_WTEMP_170),
        .b(_T_1170)
    );
    wire [5:0] _T_1172;
    wire [5:0] _WTEMP_171;
    PAD_UNSIGNED #(.width(5), .n(6)) u_pad_2112 (
        .y(_WTEMP_171),
        .in(5'h15)
    );
    MUX_UNSIGNED #(.width(6)) u_mux_2113 (
        .y(_T_1172),
        .sel(_T_1024),
        .a(_WTEMP_171),
        .b(_T_1171)
    );
    wire [5:0] _T_1173;
    wire [5:0] _WTEMP_172;
    PAD_UNSIGNED #(.width(5), .n(6)) u_pad_2114 (
        .y(_WTEMP_172),
        .in(5'h14)
    );
    MUX_UNSIGNED #(.width(6)) u_mux_2115 (
        .y(_T_1173),
        .sel(_T_1023),
        .a(_WTEMP_172),
        .b(_T_1172)
    );
    wire [5:0] _T_1174;
    wire [5:0] _WTEMP_173;
    PAD_UNSIGNED #(.width(5), .n(6)) u_pad_2116 (
        .y(_WTEMP_173),
        .in(5'h13)
    );
    MUX_UNSIGNED #(.width(6)) u_mux_2117 (
        .y(_T_1174),
        .sel(_T_1022),
        .a(_WTEMP_173),
        .b(_T_1173)
    );
    wire [5:0] _T_1175;
    wire [5:0] _WTEMP_174;
    PAD_UNSIGNED #(.width(5), .n(6)) u_pad_2118 (
        .y(_WTEMP_174),
        .in(5'h12)
    );
    MUX_UNSIGNED #(.width(6)) u_mux_2119 (
        .y(_T_1175),
        .sel(_T_1021),
        .a(_WTEMP_174),
        .b(_T_1174)
    );
    wire [5:0] _T_1176;
    wire [5:0] _WTEMP_175;
    PAD_UNSIGNED #(.width(5), .n(6)) u_pad_2120 (
        .y(_WTEMP_175),
        .in(5'h11)
    );
    MUX_UNSIGNED #(.width(6)) u_mux_2121 (
        .y(_T_1176),
        .sel(_T_1020),
        .a(_WTEMP_175),
        .b(_T_1175)
    );
    wire [5:0] _T_1177;
    wire [5:0] _WTEMP_176;
    PAD_UNSIGNED #(.width(5), .n(6)) u_pad_2122 (
        .y(_WTEMP_176),
        .in(5'h10)
    );
    MUX_UNSIGNED #(.width(6)) u_mux_2123 (
        .y(_T_1177),
        .sel(_T_1019),
        .a(_WTEMP_176),
        .b(_T_1176)
    );
    wire [5:0] _T_1178;
    wire [5:0] _WTEMP_177;
    PAD_UNSIGNED #(.width(4), .n(6)) u_pad_2124 (
        .y(_WTEMP_177),
        .in(4'hF)
    );
    MUX_UNSIGNED #(.width(6)) u_mux_2125 (
        .y(_T_1178),
        .sel(_T_1018),
        .a(_WTEMP_177),
        .b(_T_1177)
    );
    wire [5:0] _T_1179;
    wire [5:0] _WTEMP_178;
    PAD_UNSIGNED #(.width(4), .n(6)) u_pad_2126 (
        .y(_WTEMP_178),
        .in(4'hE)
    );
    MUX_UNSIGNED #(.width(6)) u_mux_2127 (
        .y(_T_1179),
        .sel(_T_1017),
        .a(_WTEMP_178),
        .b(_T_1178)
    );
    wire [5:0] _T_1180;
    wire [5:0] _WTEMP_179;
    PAD_UNSIGNED #(.width(4), .n(6)) u_pad_2128 (
        .y(_WTEMP_179),
        .in(4'hD)
    );
    MUX_UNSIGNED #(.width(6)) u_mux_2129 (
        .y(_T_1180),
        .sel(_T_1016),
        .a(_WTEMP_179),
        .b(_T_1179)
    );
    wire [5:0] _T_1181;
    wire [5:0] _WTEMP_180;
    PAD_UNSIGNED #(.width(4), .n(6)) u_pad_2130 (
        .y(_WTEMP_180),
        .in(4'hC)
    );
    MUX_UNSIGNED #(.width(6)) u_mux_2131 (
        .y(_T_1181),
        .sel(_T_1015),
        .a(_WTEMP_180),
        .b(_T_1180)
    );
    wire [5:0] _T_1182;
    wire [5:0] _WTEMP_181;
    PAD_UNSIGNED #(.width(4), .n(6)) u_pad_2132 (
        .y(_WTEMP_181),
        .in(4'hB)
    );
    MUX_UNSIGNED #(.width(6)) u_mux_2133 (
        .y(_T_1182),
        .sel(_T_1014),
        .a(_WTEMP_181),
        .b(_T_1181)
    );
    wire [5:0] _T_1183;
    wire [5:0] _WTEMP_182;
    PAD_UNSIGNED #(.width(4), .n(6)) u_pad_2134 (
        .y(_WTEMP_182),
        .in(4'hA)
    );
    MUX_UNSIGNED #(.width(6)) u_mux_2135 (
        .y(_T_1183),
        .sel(_T_1013),
        .a(_WTEMP_182),
        .b(_T_1182)
    );
    wire [5:0] _T_1184;
    wire [5:0] _WTEMP_183;
    PAD_UNSIGNED #(.width(4), .n(6)) u_pad_2136 (
        .y(_WTEMP_183),
        .in(4'h9)
    );
    MUX_UNSIGNED #(.width(6)) u_mux_2137 (
        .y(_T_1184),
        .sel(_T_1012),
        .a(_WTEMP_183),
        .b(_T_1183)
    );
    wire [5:0] _T_1185;
    wire [5:0] _WTEMP_184;
    PAD_UNSIGNED #(.width(4), .n(6)) u_pad_2138 (
        .y(_WTEMP_184),
        .in(4'h8)
    );
    MUX_UNSIGNED #(.width(6)) u_mux_2139 (
        .y(_T_1185),
        .sel(_T_1011),
        .a(_WTEMP_184),
        .b(_T_1184)
    );
    wire [5:0] _T_1186;
    wire [5:0] _WTEMP_185;
    PAD_UNSIGNED #(.width(3), .n(6)) u_pad_2140 (
        .y(_WTEMP_185),
        .in(3'h7)
    );
    MUX_UNSIGNED #(.width(6)) u_mux_2141 (
        .y(_T_1186),
        .sel(_T_1010),
        .a(_WTEMP_185),
        .b(_T_1185)
    );
    wire [5:0] _T_1187;
    wire [5:0] _WTEMP_186;
    PAD_UNSIGNED #(.width(3), .n(6)) u_pad_2142 (
        .y(_WTEMP_186),
        .in(3'h6)
    );
    MUX_UNSIGNED #(.width(6)) u_mux_2143 (
        .y(_T_1187),
        .sel(_T_1009),
        .a(_WTEMP_186),
        .b(_T_1186)
    );
    wire [5:0] _T_1188;
    wire [5:0] _WTEMP_187;
    PAD_UNSIGNED #(.width(3), .n(6)) u_pad_2144 (
        .y(_WTEMP_187),
        .in(3'h5)
    );
    MUX_UNSIGNED #(.width(6)) u_mux_2145 (
        .y(_T_1188),
        .sel(_T_1008),
        .a(_WTEMP_187),
        .b(_T_1187)
    );
    wire [5:0] _T_1189;
    wire [5:0] _WTEMP_188;
    PAD_UNSIGNED #(.width(3), .n(6)) u_pad_2146 (
        .y(_WTEMP_188),
        .in(3'h4)
    );
    MUX_UNSIGNED #(.width(6)) u_mux_2147 (
        .y(_T_1189),
        .sel(_T_1007),
        .a(_WTEMP_188),
        .b(_T_1188)
    );
    wire [5:0] _T_1190;
    wire [5:0] _WTEMP_189;
    PAD_UNSIGNED #(.width(2), .n(6)) u_pad_2148 (
        .y(_WTEMP_189),
        .in(2'h3)
    );
    MUX_UNSIGNED #(.width(6)) u_mux_2149 (
        .y(_T_1190),
        .sel(_T_1006),
        .a(_WTEMP_189),
        .b(_T_1189)
    );
    wire [5:0] _T_1191;
    wire [5:0] _WTEMP_190;
    PAD_UNSIGNED #(.width(2), .n(6)) u_pad_2150 (
        .y(_WTEMP_190),
        .in(2'h2)
    );
    MUX_UNSIGNED #(.width(6)) u_mux_2151 (
        .y(_T_1191),
        .sel(_T_1005),
        .a(_WTEMP_190),
        .b(_T_1190)
    );
    wire [5:0] _T_1192;
    wire [5:0] _WTEMP_191;
    PAD_UNSIGNED #(.width(1), .n(6)) u_pad_2152 (
        .y(_WTEMP_191),
        .in(1'h1)
    );
    MUX_UNSIGNED #(.width(6)) u_mux_2153 (
        .y(_T_1192),
        .sel(_T_1004),
        .a(_WTEMP_191),
        .b(_T_1191)
    );
    wire [5:0] _T_1193;
    wire [5:0] _WTEMP_192;
    PAD_UNSIGNED #(.width(1), .n(6)) u_pad_2154 (
        .y(_WTEMP_192),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(6)) u_mux_2155 (
        .y(_T_1193),
        .sel(_T_1003),
        .a(_WTEMP_192),
        .b(_T_1192)
    );
    wire [64:0] _T_1194;
    wire [63:0] _WTEMP_193;
    PAD_UNSIGNED #(.width(6), .n(64)) u_pad_2156 (
        .y(_WTEMP_193),
        .in(_T_1193)
    );
    ADD_UNSIGNED #(.width(64)) u_add_2157 (
        .y(_T_1194),
        .a(64'h8000000000000000),
        .b(_WTEMP_193)
    );
    wire [63:0] interruptCause;
    TAIL #(.width(65), .n(1)) tail_2158 (
        .y(interruptCause),
        .in(_T_1194)
    );
    wire _T_1196;
    wire [63:0] _WTEMP_194;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_2159 (
        .y(_WTEMP_194),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(64)) u_neq_2160 (
        .y(_T_1196),
        .a(all_interrupts),
        .b(_WTEMP_194)
    );
    wire _T_1198;
    EQ_UNSIGNED #(.width(1)) u_eq_2161 (
        .y(_T_1198),
        .a(_reg_debug__q),
        .b(1'h0)
    );
    wire _T_1199;
    BITWISEAND #(.width(1)) bitwiseand_2162 (
        .y(_T_1199),
        .a(_T_1196),
        .b(_T_1198)
    );
    wire _T_1201;
    EQ_UNSIGNED #(.width(1)) u_eq_2163 (
        .y(_T_1201),
        .a(io_singleStep),
        .b(1'h0)
    );
    wire _T_1202;
    BITWISEAND #(.width(1)) bitwiseand_2164 (
        .y(_T_1202),
        .a(_T_1199),
        .b(_T_1201)
    );
    wire _T_1203;
    BITWISEOR #(.width(1)) bitwiseor_2165 (
        .y(_T_1203),
        .a(_T_1202),
        .b(_reg_singleStepped__q)
    );
    wire _T_1205;
    BITWISEAND #(.width(1)) bitwiseand_2166 (
        .y(_T_1205),
        .a(1'h1),
        .b(_reg_dcsr_debugint__q)
    );
    wire _T_1207;
    EQ_UNSIGNED #(.width(1)) u_eq_2167 (
        .y(_T_1207),
        .a(_reg_debug__q),
        .b(1'h0)
    );
    wire _T_1208;
    BITWISEAND #(.width(1)) bitwiseand_2168 (
        .y(_T_1208),
        .a(_T_1205),
        .b(_T_1207)
    );
    wire [64:0] _T_1226;
    assign _T_1226 = 65'h800000000000000D;
    wire [63:0] _T_1227;
    assign _T_1227 = 64'h800000000000000D;
    wire [63:0] _reg_misa__q;
    wire [63:0] _reg_misa__d;
    DFF_POSCLK #(.width(64)) reg_misa (
        .q(_reg_misa__q),
        .d(_reg_misa__d),
        .clk(clock)
    );
    wire [63:0] _WTEMP_195;
    MUX_UNSIGNED #(.width(64)) u_mux_2169 (
        .y(_reg_misa__d),
        .sel(reset),
        .a(64'h800000000014112D),
        .b(_WTEMP_195)
    );
    wire [1:0] _T_1229;
    CAT #(.width_a(1), .width_b(1)) cat_2170 (
        .y(_T_1229),
        .a(io_status_hie),
        .b(io_status_sie)
    );
    wire [2:0] _T_1230;
    CAT #(.width_a(2), .width_b(1)) cat_2171 (
        .y(_T_1230),
        .a(_T_1229),
        .b(io_status_uie)
    );
    wire [1:0] _T_1231;
    CAT #(.width_a(1), .width_b(1)) cat_2172 (
        .y(_T_1231),
        .a(io_status_upie),
        .b(io_status_mie)
    );
    wire [1:0] _T_1232;
    CAT #(.width_a(1), .width_b(1)) cat_2173 (
        .y(_T_1232),
        .a(io_status_hpie),
        .b(io_status_spie)
    );
    wire [3:0] _T_1233;
    CAT #(.width_a(2), .width_b(2)) cat_2174 (
        .y(_T_1233),
        .a(_T_1232),
        .b(_T_1231)
    );
    wire [6:0] _T_1234;
    CAT #(.width_a(4), .width_b(3)) cat_2175 (
        .y(_T_1234),
        .a(_T_1233),
        .b(_T_1230)
    );
    wire [2:0] _T_1235;
    CAT #(.width_a(2), .width_b(1)) cat_2176 (
        .y(_T_1235),
        .a(io_status_hpp),
        .b(io_status_spp)
    );
    wire [3:0] _T_1236;
    CAT #(.width_a(3), .width_b(1)) cat_2177 (
        .y(_T_1236),
        .a(_T_1235),
        .b(io_status_mpie)
    );
    wire [3:0] _T_1237;
    CAT #(.width_a(2), .width_b(2)) cat_2178 (
        .y(_T_1237),
        .a(io_status_fs),
        .b(io_status_mpp)
    );
    wire [2:0] _T_1238;
    CAT #(.width_a(1), .width_b(2)) cat_2179 (
        .y(_T_1238),
        .a(io_status_mprv),
        .b(io_status_xs)
    );
    wire [6:0] _T_1239;
    CAT #(.width_a(3), .width_b(4)) cat_2180 (
        .y(_T_1239),
        .a(_T_1238),
        .b(_T_1237)
    );
    wire [10:0] _T_1240;
    CAT #(.width_a(7), .width_b(4)) cat_2181 (
        .y(_T_1240),
        .a(_T_1239),
        .b(_T_1236)
    );
    wire [17:0] _T_1241;
    CAT #(.width_a(11), .width_b(7)) cat_2182 (
        .y(_T_1241),
        .a(_T_1240),
        .b(_T_1234)
    );
    wire [1:0] _T_1242;
    CAT #(.width_a(1), .width_b(1)) cat_2183 (
        .y(_T_1242),
        .a(io_status_tvm),
        .b(io_status_mxr)
    );
    wire [2:0] _T_1243;
    CAT #(.width_a(2), .width_b(1)) cat_2184 (
        .y(_T_1243),
        .a(_T_1242),
        .b(io_status_pum)
    );
    wire [1:0] _T_1244;
    CAT #(.width_a(1), .width_b(1)) cat_2185 (
        .y(_T_1244),
        .a(io_status_tsr),
        .b(io_status_tw)
    );
    wire [8:0] _T_1245;
    CAT #(.width_a(1), .width_b(8)) cat_2186 (
        .y(_T_1245),
        .a(io_status_sd_rv32),
        .b(io_status_zero1)
    );
    wire [10:0] _T_1246;
    CAT #(.width_a(9), .width_b(2)) cat_2187 (
        .y(_T_1246),
        .a(_T_1245),
        .b(_T_1244)
    );
    wire [13:0] _T_1247;
    CAT #(.width_a(11), .width_b(3)) cat_2188 (
        .y(_T_1247),
        .a(_T_1246),
        .b(_T_1243)
    );
    wire [28:0] _T_1248;
    CAT #(.width_a(27), .width_b(2)) cat_2189 (
        .y(_T_1248),
        .a(io_status_zero2),
        .b(io_status_sxl)
    );
    wire [30:0] _T_1249;
    CAT #(.width_a(29), .width_b(2)) cat_2190 (
        .y(_T_1249),
        .a(_T_1248),
        .b(io_status_uxl)
    );
    wire [2:0] _T_1250;
    CAT #(.width_a(2), .width_b(1)) cat_2191 (
        .y(_T_1250),
        .a(io_status_prv),
        .b(io_status_sd)
    );
    wire [32:0] _T_1251;
    CAT #(.width_a(1), .width_b(32)) cat_2192 (
        .y(_T_1251),
        .a(io_status_debug),
        .b(io_status_isa)
    );
    wire [35:0] _T_1252;
    CAT #(.width_a(33), .width_b(3)) cat_2193 (
        .y(_T_1252),
        .a(_T_1251),
        .b(_T_1250)
    );
    wire [66:0] _T_1253;
    CAT #(.width_a(36), .width_b(31)) cat_2194 (
        .y(_T_1253),
        .a(_T_1252),
        .b(_T_1249)
    );
    wire [80:0] _T_1254;
    CAT #(.width_a(67), .width_b(14)) cat_2195 (
        .y(_T_1254),
        .a(_T_1253),
        .b(_T_1247)
    );
    wire [98:0] _T_1255;
    CAT #(.width_a(81), .width_b(18)) cat_2196 (
        .y(_T_1255),
        .a(_T_1254),
        .b(_T_1241)
    );
    wire [63:0] read_mstatus;
    BITS #(.width(99), .high(63), .low(0)) bits_2197 (
        .y(read_mstatus),
        .in(_T_1255)
    );
    wire [1:0] _T_1291;
    CAT #(.width_a(1), .width_b(1)) cat_2198 (
        .y(_T_1291),
        .a(_reg_bp_0_control_x__q),
        .b(_reg_bp_0_control_w__q)
    );
    wire [2:0] _T_1292;
    CAT #(.width_a(2), .width_b(1)) cat_2199 (
        .y(_T_1292),
        .a(_T_1291),
        .b(_reg_bp_0_control_r__q)
    );
    wire [1:0] _T_1293;
    CAT #(.width_a(1), .width_b(1)) cat_2200 (
        .y(_T_1293),
        .a(_reg_bp_0_control_s__q),
        .b(_reg_bp_0_control_u__q)
    );
    wire [1:0] _T_1294;
    CAT #(.width_a(1), .width_b(1)) cat_2201 (
        .y(_T_1294),
        .a(_reg_bp_0_control_m__q),
        .b(1'h0)
    );
    wire [3:0] _T_1295;
    CAT #(.width_a(2), .width_b(2)) cat_2202 (
        .y(_T_1295),
        .a(_T_1294),
        .b(_T_1293)
    );
    wire [6:0] _T_1296;
    CAT #(.width_a(4), .width_b(3)) cat_2203 (
        .y(_T_1296),
        .a(_T_1295),
        .b(_T_1292)
    );
    wire [3:0] _T_1297;
    CAT #(.width_a(2), .width_b(2)) cat_2204 (
        .y(_T_1297),
        .a(2'h0),
        .b(_reg_bp_0_control_tmatch__q)
    );
    wire [1:0] _T_1298;
    CAT #(.width_a(1), .width_b(1)) cat_2205 (
        .y(_T_1298),
        .a(_reg_bp_0_control_action__q),
        .b(1'h0)
    );
    wire [5:0] _T_1299;
    CAT #(.width_a(2), .width_b(4)) cat_2206 (
        .y(_T_1299),
        .a(_T_1298),
        .b(_T_1297)
    );
    wire [4:0] _T_1301;
    CAT #(.width_a(4), .width_b(1)) cat_2207 (
        .y(_T_1301),
        .a(4'h2),
        .b(_reg_bp_0_control_dmode__q)
    );
    wire [50:0] _T_1302;
    CAT #(.width_a(5), .width_b(46)) cat_2208 (
        .y(_T_1302),
        .a(_T_1301),
        .b(46'h40000000000)
    );
    wire [56:0] _T_1303;
    CAT #(.width_a(51), .width_b(6)) cat_2209 (
        .y(_T_1303),
        .a(_T_1302),
        .b(_T_1299)
    );
    wire [63:0] _T_1304;
    CAT #(.width_a(57), .width_b(7)) cat_2210 (
        .y(_T_1304),
        .a(_T_1303),
        .b(_T_1296)
    );
    wire _T_1340;
    BITS #(.width(39), .high(38), .low(38)) bits_2211 (
        .y(_T_1340),
        .in(_reg_bp_0_address__q)
    );
    wire _T_1341;
    BITS #(.width(1), .high(0), .low(0)) bits_2212 (
        .y(_T_1341),
        .in(_T_1340)
    );
    wire [24:0] _T_1344;
    MUX_UNSIGNED #(.width(25)) u_mux_2213 (
        .y(_T_1344),
        .sel(_T_1341),
        .a(25'h1FFFFFF),
        .b(25'h0)
    );
    wire [63:0] _T_1345;
    CAT #(.width_a(25), .width_b(39)) cat_2214 (
        .y(_T_1345),
        .a(_T_1344),
        .b(_reg_bp_0_address__q)
    );
    wire _T_1349;
    BITS #(.width(40), .high(39), .low(39)) bits_2215 (
        .y(_T_1349),
        .in(_reg_mepc__q)
    );
    wire _T_1350;
    BITS #(.width(1), .high(0), .low(0)) bits_2216 (
        .y(_T_1350),
        .in(_T_1349)
    );
    wire [23:0] _T_1353;
    MUX_UNSIGNED #(.width(24)) u_mux_2217 (
        .y(_T_1353),
        .sel(_T_1350),
        .a(24'hFFFFFF),
        .b(24'h0)
    );
    wire [63:0] _T_1354;
    CAT #(.width_a(24), .width_b(40)) cat_2218 (
        .y(_T_1354),
        .a(_T_1353),
        .b(_reg_mepc__q)
    );
    wire _T_1355;
    BITS #(.width(40), .high(39), .low(39)) bits_2219 (
        .y(_T_1355),
        .in(_reg_mbadaddr__q)
    );
    wire _T_1356;
    BITS #(.width(1), .high(0), .low(0)) bits_2220 (
        .y(_T_1356),
        .in(_T_1355)
    );
    wire [23:0] _T_1359;
    MUX_UNSIGNED #(.width(24)) u_mux_2221 (
        .y(_T_1359),
        .sel(_T_1356),
        .a(24'hFFFFFF),
        .b(24'h0)
    );
    wire [63:0] _T_1360;
    CAT #(.width_a(24), .width_b(40)) cat_2222 (
        .y(_T_1360),
        .a(_T_1359),
        .b(_reg_mbadaddr__q)
    );
    wire [2:0] _T_1361;
    CAT #(.width_a(1), .width_b(2)) cat_2223 (
        .y(_T_1361),
        .a(_reg_dcsr_step__q),
        .b(_reg_dcsr_prv__q)
    );
    wire [1:0] _T_1362;
    CAT #(.width_a(1), .width_b(1)) cat_2224 (
        .y(_T_1362),
        .a(1'h0),
        .b(_reg_dcsr_halt__q)
    );
    wire [4:0] _T_1363;
    CAT #(.width_a(2), .width_b(3)) cat_2225 (
        .y(_T_1363),
        .a(_T_1362),
        .b(_T_1361)
    );
    wire [3:0] _T_1364;
    CAT #(.width_a(3), .width_b(1)) cat_2226 (
        .y(_T_1364),
        .a(_reg_dcsr_cause__q),
        .b(_reg_dcsr_debugint__q)
    );
    wire [1:0] _T_1365;
    assign _T_1365 = 2'h0;
    wire [5:0] _T_1366;
    CAT #(.width_a(2), .width_b(4)) cat_2227 (
        .y(_T_1366),
        .a(_T_1365),
        .b(_T_1364)
    );
    wire [10:0] _T_1367;
    CAT #(.width_a(6), .width_b(5)) cat_2228 (
        .y(_T_1367),
        .a(_T_1366),
        .b(_T_1363)
    );
    wire [1:0] _T_1368;
    CAT #(.width_a(1), .width_b(1)) cat_2229 (
        .y(_T_1368),
        .a(_reg_dcsr_ebreaku__q),
        .b(1'h0)
    );
    wire [1:0] _T_1369;
    CAT #(.width_a(1), .width_b(1)) cat_2230 (
        .y(_T_1369),
        .a(1'h0),
        .b(_reg_dcsr_ebreaks__q)
    );
    wire [3:0] _T_1370;
    CAT #(.width_a(2), .width_b(2)) cat_2231 (
        .y(_T_1370),
        .a(_T_1369),
        .b(_T_1368)
    );
    wire [12:0] _T_1371;
    CAT #(.width_a(12), .width_b(1)) cat_2232 (
        .y(_T_1371),
        .a(12'h0),
        .b(_reg_dcsr_ebreakm__q)
    );
    wire [2:0] _T_1372;
    assign _T_1372 = 3'h2;
    wire [3:0] _T_1373;
    assign _T_1373 = 4'h4;
    wire [16:0] _T_1374;
    CAT #(.width_a(4), .width_b(13)) cat_2233 (
        .y(_T_1374),
        .a(_T_1373),
        .b(_T_1371)
    );
    wire [20:0] _T_1375;
    CAT #(.width_a(17), .width_b(4)) cat_2234 (
        .y(_T_1375),
        .a(_T_1374),
        .b(_T_1370)
    );
    wire [31:0] _T_1376;
    CAT #(.width_a(21), .width_b(11)) cat_2235 (
        .y(_T_1376),
        .a(_T_1375),
        .b(_T_1367)
    );
    wire [7:0] _T_1377;
    CAT #(.width_a(3), .width_b(5)) cat_2236 (
        .y(_T_1377),
        .a(_reg_frm__q),
        .b(_reg_fflags__q)
    );
    wire [63:0] _T_1380;
    BITWISEAND #(.width(64)) bitwiseand_2237 (
        .y(_T_1380),
        .a(_reg_mie__q),
        .b(_reg_mideleg__q)
    );
    wire [63:0] _T_1381;
    wire [63:0] _WTEMP_196;
    PAD_UNSIGNED #(.width(13), .n(64)) u_pad_2238 (
        .y(_WTEMP_196),
        .in(read_mip)
    );
    BITWISEAND #(.width(64)) bitwiseand_2239 (
        .y(_T_1381),
        .a(_WTEMP_196),
        .b(_reg_mideleg__q)
    );
    wire _T_1382_debug;
    wire [31:0] _T_1382_isa;
    wire [1:0] _T_1382_prv;
    wire _T_1382_sd;
    wire [26:0] _T_1382_zero2;
    wire [1:0] _T_1382_sxl;
    wire [1:0] _T_1382_uxl;
    wire _T_1382_sd_rv32;
    wire [7:0] _T_1382_zero1;
    wire _T_1382_tsr;
    wire _T_1382_tw;
    wire _T_1382_tvm;
    wire _T_1382_mxr;
    wire _T_1382_pum;
    wire _T_1382_mprv;
    wire [1:0] _T_1382_xs;
    wire [1:0] _T_1382_fs;
    wire [1:0] _T_1382_mpp;
    wire [1:0] _T_1382_hpp;
    wire _T_1382_spp;
    wire _T_1382_mpie;
    wire _T_1382_hpie;
    wire _T_1382_spie;
    wire _T_1382_upie;
    wire _T_1382_mie;
    wire _T_1382_hie;
    wire _T_1382_sie;
    wire _T_1382_uie;
    wire [1:0] _T_1418;
    CAT #(.width_a(1), .width_b(1)) cat_2240 (
        .y(_T_1418),
        .a(_T_1382_hie),
        .b(_T_1382_sie)
    );
    wire [2:0] _T_1419;
    CAT #(.width_a(2), .width_b(1)) cat_2241 (
        .y(_T_1419),
        .a(_T_1418),
        .b(_T_1382_uie)
    );
    wire [1:0] _T_1420;
    CAT #(.width_a(1), .width_b(1)) cat_2242 (
        .y(_T_1420),
        .a(_T_1382_upie),
        .b(_T_1382_mie)
    );
    wire [1:0] _T_1421;
    CAT #(.width_a(1), .width_b(1)) cat_2243 (
        .y(_T_1421),
        .a(_T_1382_hpie),
        .b(_T_1382_spie)
    );
    wire [3:0] _T_1422;
    CAT #(.width_a(2), .width_b(2)) cat_2244 (
        .y(_T_1422),
        .a(_T_1421),
        .b(_T_1420)
    );
    wire [6:0] _T_1423;
    CAT #(.width_a(4), .width_b(3)) cat_2245 (
        .y(_T_1423),
        .a(_T_1422),
        .b(_T_1419)
    );
    wire [2:0] _T_1424;
    CAT #(.width_a(2), .width_b(1)) cat_2246 (
        .y(_T_1424),
        .a(_T_1382_hpp),
        .b(_T_1382_spp)
    );
    wire [3:0] _T_1425;
    CAT #(.width_a(3), .width_b(1)) cat_2247 (
        .y(_T_1425),
        .a(_T_1424),
        .b(_T_1382_mpie)
    );
    wire [3:0] _T_1426;
    CAT #(.width_a(2), .width_b(2)) cat_2248 (
        .y(_T_1426),
        .a(_T_1382_fs),
        .b(_T_1382_mpp)
    );
    wire [2:0] _T_1427;
    CAT #(.width_a(1), .width_b(2)) cat_2249 (
        .y(_T_1427),
        .a(_T_1382_mprv),
        .b(_T_1382_xs)
    );
    wire [6:0] _T_1428;
    CAT #(.width_a(3), .width_b(4)) cat_2250 (
        .y(_T_1428),
        .a(_T_1427),
        .b(_T_1426)
    );
    wire [10:0] _T_1429;
    CAT #(.width_a(7), .width_b(4)) cat_2251 (
        .y(_T_1429),
        .a(_T_1428),
        .b(_T_1425)
    );
    wire [17:0] _T_1430;
    CAT #(.width_a(11), .width_b(7)) cat_2252 (
        .y(_T_1430),
        .a(_T_1429),
        .b(_T_1423)
    );
    wire [1:0] _T_1431;
    CAT #(.width_a(1), .width_b(1)) cat_2253 (
        .y(_T_1431),
        .a(_T_1382_tvm),
        .b(_T_1382_mxr)
    );
    wire [2:0] _T_1432;
    CAT #(.width_a(2), .width_b(1)) cat_2254 (
        .y(_T_1432),
        .a(_T_1431),
        .b(_T_1382_pum)
    );
    wire [1:0] _T_1433;
    CAT #(.width_a(1), .width_b(1)) cat_2255 (
        .y(_T_1433),
        .a(_T_1382_tsr),
        .b(_T_1382_tw)
    );
    wire [8:0] _T_1434;
    CAT #(.width_a(1), .width_b(8)) cat_2256 (
        .y(_T_1434),
        .a(_T_1382_sd_rv32),
        .b(_T_1382_zero1)
    );
    wire [10:0] _T_1435;
    CAT #(.width_a(9), .width_b(2)) cat_2257 (
        .y(_T_1435),
        .a(_T_1434),
        .b(_T_1433)
    );
    wire [13:0] _T_1436;
    CAT #(.width_a(11), .width_b(3)) cat_2258 (
        .y(_T_1436),
        .a(_T_1435),
        .b(_T_1432)
    );
    wire [28:0] _T_1437;
    CAT #(.width_a(27), .width_b(2)) cat_2259 (
        .y(_T_1437),
        .a(_T_1382_zero2),
        .b(_T_1382_sxl)
    );
    wire [30:0] _T_1438;
    CAT #(.width_a(29), .width_b(2)) cat_2260 (
        .y(_T_1438),
        .a(_T_1437),
        .b(_T_1382_uxl)
    );
    wire [2:0] _T_1439;
    CAT #(.width_a(2), .width_b(1)) cat_2261 (
        .y(_T_1439),
        .a(_T_1382_prv),
        .b(_T_1382_sd)
    );
    wire [32:0] _T_1440;
    CAT #(.width_a(1), .width_b(32)) cat_2262 (
        .y(_T_1440),
        .a(_T_1382_debug),
        .b(_T_1382_isa)
    );
    wire [35:0] _T_1441;
    CAT #(.width_a(33), .width_b(3)) cat_2263 (
        .y(_T_1441),
        .a(_T_1440),
        .b(_T_1439)
    );
    wire [66:0] _T_1442;
    CAT #(.width_a(36), .width_b(31)) cat_2264 (
        .y(_T_1442),
        .a(_T_1441),
        .b(_T_1438)
    );
    wire [80:0] _T_1443;
    CAT #(.width_a(67), .width_b(14)) cat_2265 (
        .y(_T_1443),
        .a(_T_1442),
        .b(_T_1436)
    );
    wire [98:0] _T_1444;
    CAT #(.width_a(81), .width_b(18)) cat_2266 (
        .y(_T_1444),
        .a(_T_1443),
        .b(_T_1430)
    );
    wire [63:0] _T_1445;
    BITS #(.width(99), .high(63), .low(0)) bits_2267 (
        .y(_T_1445),
        .in(_T_1444)
    );
    wire _T_1446;
    BITS #(.width(40), .high(39), .low(39)) bits_2268 (
        .y(_T_1446),
        .in(_reg_sbadaddr__q)
    );
    wire _T_1447;
    BITS #(.width(1), .high(0), .low(0)) bits_2269 (
        .y(_T_1447),
        .in(_T_1446)
    );
    wire [23:0] _T_1450;
    MUX_UNSIGNED #(.width(24)) u_mux_2270 (
        .y(_T_1450),
        .sel(_T_1447),
        .a(24'hFFFFFF),
        .b(24'h0)
    );
    wire [63:0] _T_1451;
    CAT #(.width_a(24), .width_b(40)) cat_2271 (
        .y(_T_1451),
        .a(_T_1450),
        .b(_reg_sbadaddr__q)
    );
    wire [19:0] _T_1452;
    CAT #(.width_a(4), .width_b(16)) cat_2272 (
        .y(_T_1452),
        .a(_reg_sptbr_mode__q),
        .b(16'h0)
    );
    wire [63:0] _T_1453;
    CAT #(.width_a(20), .width_b(44)) cat_2273 (
        .y(_T_1453),
        .a(_T_1452),
        .b(_reg_sptbr_ppn__q)
    );
    wire _T_1454;
    BITS #(.width(40), .high(39), .low(39)) bits_2274 (
        .y(_T_1454),
        .in(_reg_sepc__q)
    );
    wire _T_1455;
    BITS #(.width(1), .high(0), .low(0)) bits_2275 (
        .y(_T_1455),
        .in(_T_1454)
    );
    wire [23:0] _T_1458;
    MUX_UNSIGNED #(.width(24)) u_mux_2276 (
        .y(_T_1458),
        .sel(_T_1455),
        .a(24'hFFFFFF),
        .b(24'h0)
    );
    wire [63:0] _T_1459;
    CAT #(.width_a(24), .width_b(40)) cat_2277 (
        .y(_T_1459),
        .a(_T_1458),
        .b(_reg_sepc__q)
    );
    wire _T_1460;
    BITS #(.width(39), .high(38), .low(38)) bits_2278 (
        .y(_T_1460),
        .in(_reg_stvec__q)
    );
    wire _T_1461;
    BITS #(.width(1), .high(0), .low(0)) bits_2279 (
        .y(_T_1461),
        .in(_T_1460)
    );
    wire [24:0] _T_1464;
    MUX_UNSIGNED #(.width(25)) u_mux_2280 (
        .y(_T_1464),
        .sel(_T_1461),
        .a(25'h1FFFFFF),
        .b(25'h0)
    );
    wire [63:0] _T_1465;
    CAT #(.width_a(25), .width_b(39)) cat_2281 (
        .y(_T_1465),
        .a(_T_1464),
        .b(_reg_stvec__q)
    );
    wire _T_1467;
    wire [11:0] _WTEMP_197;
    PAD_UNSIGNED #(.width(11), .n(12)) u_pad_2282 (
        .y(_WTEMP_197),
        .in(11'h7A0)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2283 (
        .y(_T_1467),
        .a(io_rw_addr),
        .b(_WTEMP_197)
    );
    wire _T_1469;
    wire [11:0] _WTEMP_198;
    PAD_UNSIGNED #(.width(11), .n(12)) u_pad_2284 (
        .y(_WTEMP_198),
        .in(11'h7A1)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2285 (
        .y(_T_1469),
        .a(io_rw_addr),
        .b(_WTEMP_198)
    );
    wire _T_1471;
    wire [11:0] _WTEMP_199;
    PAD_UNSIGNED #(.width(11), .n(12)) u_pad_2286 (
        .y(_WTEMP_199),
        .in(11'h7A2)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2287 (
        .y(_T_1471),
        .a(io_rw_addr),
        .b(_WTEMP_199)
    );
    wire _T_1473;
    EQ_UNSIGNED #(.width(12)) u_eq_2288 (
        .y(_T_1473),
        .a(io_rw_addr),
        .b(12'hF13)
    );
    wire _T_1475;
    EQ_UNSIGNED #(.width(12)) u_eq_2289 (
        .y(_T_1475),
        .a(io_rw_addr),
        .b(12'hF12)
    );
    wire _T_1477;
    EQ_UNSIGNED #(.width(12)) u_eq_2290 (
        .y(_T_1477),
        .a(io_rw_addr),
        .b(12'hF11)
    );
    wire _T_1479;
    EQ_UNSIGNED #(.width(12)) u_eq_2291 (
        .y(_T_1479),
        .a(io_rw_addr),
        .b(12'hB00)
    );
    wire _T_1481;
    EQ_UNSIGNED #(.width(12)) u_eq_2292 (
        .y(_T_1481),
        .a(io_rw_addr),
        .b(12'hB02)
    );
    wire _T_1483;
    wire [11:0] _WTEMP_200;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2293 (
        .y(_WTEMP_200),
        .in(10'h301)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2294 (
        .y(_T_1483),
        .a(io_rw_addr),
        .b(_WTEMP_200)
    );
    wire _T_1485;
    wire [11:0] _WTEMP_201;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2295 (
        .y(_WTEMP_201),
        .in(10'h300)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2296 (
        .y(_T_1485),
        .a(io_rw_addr),
        .b(_WTEMP_201)
    );
    wire _T_1487;
    wire [11:0] _WTEMP_202;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2297 (
        .y(_WTEMP_202),
        .in(10'h305)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2298 (
        .y(_T_1487),
        .a(io_rw_addr),
        .b(_WTEMP_202)
    );
    wire _T_1489;
    wire [11:0] _WTEMP_203;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2299 (
        .y(_WTEMP_203),
        .in(10'h344)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2300 (
        .y(_T_1489),
        .a(io_rw_addr),
        .b(_WTEMP_203)
    );
    wire _T_1491;
    wire [11:0] _WTEMP_204;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2301 (
        .y(_WTEMP_204),
        .in(10'h304)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2302 (
        .y(_T_1491),
        .a(io_rw_addr),
        .b(_WTEMP_204)
    );
    wire _T_1493;
    wire [11:0] _WTEMP_205;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2303 (
        .y(_WTEMP_205),
        .in(10'h303)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2304 (
        .y(_T_1493),
        .a(io_rw_addr),
        .b(_WTEMP_205)
    );
    wire _T_1495;
    wire [11:0] _WTEMP_206;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2305 (
        .y(_WTEMP_206),
        .in(10'h302)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2306 (
        .y(_T_1495),
        .a(io_rw_addr),
        .b(_WTEMP_206)
    );
    wire _T_1497;
    wire [11:0] _WTEMP_207;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2307 (
        .y(_WTEMP_207),
        .in(10'h340)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2308 (
        .y(_T_1497),
        .a(io_rw_addr),
        .b(_WTEMP_207)
    );
    wire _T_1499;
    wire [11:0] _WTEMP_208;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2309 (
        .y(_WTEMP_208),
        .in(10'h341)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2310 (
        .y(_T_1499),
        .a(io_rw_addr),
        .b(_WTEMP_208)
    );
    wire _T_1501;
    wire [11:0] _WTEMP_209;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2311 (
        .y(_WTEMP_209),
        .in(10'h343)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2312 (
        .y(_T_1501),
        .a(io_rw_addr),
        .b(_WTEMP_209)
    );
    wire _T_1503;
    wire [11:0] _WTEMP_210;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2313 (
        .y(_WTEMP_210),
        .in(10'h342)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2314 (
        .y(_T_1503),
        .a(io_rw_addr),
        .b(_WTEMP_210)
    );
    wire _T_1505;
    EQ_UNSIGNED #(.width(12)) u_eq_2315 (
        .y(_T_1505),
        .a(io_rw_addr),
        .b(12'hF14)
    );
    wire _T_1507;
    wire [11:0] _WTEMP_211;
    PAD_UNSIGNED #(.width(11), .n(12)) u_pad_2316 (
        .y(_WTEMP_211),
        .in(11'h7B0)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2317 (
        .y(_T_1507),
        .a(io_rw_addr),
        .b(_WTEMP_211)
    );
    wire _T_1509;
    wire [11:0] _WTEMP_212;
    PAD_UNSIGNED #(.width(11), .n(12)) u_pad_2318 (
        .y(_WTEMP_212),
        .in(11'h7B1)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2319 (
        .y(_T_1509),
        .a(io_rw_addr),
        .b(_WTEMP_212)
    );
    wire _T_1511;
    wire [11:0] _WTEMP_213;
    PAD_UNSIGNED #(.width(11), .n(12)) u_pad_2320 (
        .y(_WTEMP_213),
        .in(11'h7B2)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2321 (
        .y(_T_1511),
        .a(io_rw_addr),
        .b(_WTEMP_213)
    );
    wire _T_1513;
    wire [11:0] _WTEMP_214;
    PAD_UNSIGNED #(.width(1), .n(12)) u_pad_2322 (
        .y(_WTEMP_214),
        .in(1'h1)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2323 (
        .y(_T_1513),
        .a(io_rw_addr),
        .b(_WTEMP_214)
    );
    wire _T_1515;
    wire [11:0] _WTEMP_215;
    PAD_UNSIGNED #(.width(2), .n(12)) u_pad_2324 (
        .y(_WTEMP_215),
        .in(2'h2)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2325 (
        .y(_T_1515),
        .a(io_rw_addr),
        .b(_WTEMP_215)
    );
    wire _T_1517;
    wire [11:0] _WTEMP_216;
    PAD_UNSIGNED #(.width(2), .n(12)) u_pad_2326 (
        .y(_WTEMP_216),
        .in(2'h3)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2327 (
        .y(_T_1517),
        .a(io_rw_addr),
        .b(_WTEMP_216)
    );
    wire _T_1519;
    wire [11:0] _WTEMP_217;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2328 (
        .y(_WTEMP_217),
        .in(10'h323)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2329 (
        .y(_T_1519),
        .a(io_rw_addr),
        .b(_WTEMP_217)
    );
    wire _T_1521;
    EQ_UNSIGNED #(.width(12)) u_eq_2330 (
        .y(_T_1521),
        .a(io_rw_addr),
        .b(12'hB03)
    );
    wire _T_1523;
    EQ_UNSIGNED #(.width(12)) u_eq_2331 (
        .y(_T_1523),
        .a(io_rw_addr),
        .b(12'hC03)
    );
    wire _T_1525;
    wire [11:0] _WTEMP_218;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2332 (
        .y(_WTEMP_218),
        .in(10'h324)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2333 (
        .y(_T_1525),
        .a(io_rw_addr),
        .b(_WTEMP_218)
    );
    wire _T_1527;
    EQ_UNSIGNED #(.width(12)) u_eq_2334 (
        .y(_T_1527),
        .a(io_rw_addr),
        .b(12'hB04)
    );
    wire _T_1529;
    EQ_UNSIGNED #(.width(12)) u_eq_2335 (
        .y(_T_1529),
        .a(io_rw_addr),
        .b(12'hC04)
    );
    wire _T_1531;
    wire [11:0] _WTEMP_219;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2336 (
        .y(_WTEMP_219),
        .in(10'h325)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2337 (
        .y(_T_1531),
        .a(io_rw_addr),
        .b(_WTEMP_219)
    );
    wire _T_1533;
    EQ_UNSIGNED #(.width(12)) u_eq_2338 (
        .y(_T_1533),
        .a(io_rw_addr),
        .b(12'hB05)
    );
    wire _T_1535;
    EQ_UNSIGNED #(.width(12)) u_eq_2339 (
        .y(_T_1535),
        .a(io_rw_addr),
        .b(12'hC05)
    );
    wire _T_1537;
    wire [11:0] _WTEMP_220;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2340 (
        .y(_WTEMP_220),
        .in(10'h326)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2341 (
        .y(_T_1537),
        .a(io_rw_addr),
        .b(_WTEMP_220)
    );
    wire _T_1539;
    EQ_UNSIGNED #(.width(12)) u_eq_2342 (
        .y(_T_1539),
        .a(io_rw_addr),
        .b(12'hB06)
    );
    wire _T_1541;
    EQ_UNSIGNED #(.width(12)) u_eq_2343 (
        .y(_T_1541),
        .a(io_rw_addr),
        .b(12'hC06)
    );
    wire _T_1543;
    wire [11:0] _WTEMP_221;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2344 (
        .y(_WTEMP_221),
        .in(10'h327)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2345 (
        .y(_T_1543),
        .a(io_rw_addr),
        .b(_WTEMP_221)
    );
    wire _T_1545;
    EQ_UNSIGNED #(.width(12)) u_eq_2346 (
        .y(_T_1545),
        .a(io_rw_addr),
        .b(12'hB07)
    );
    wire _T_1547;
    EQ_UNSIGNED #(.width(12)) u_eq_2347 (
        .y(_T_1547),
        .a(io_rw_addr),
        .b(12'hC07)
    );
    wire _T_1549;
    wire [11:0] _WTEMP_222;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2348 (
        .y(_WTEMP_222),
        .in(10'h328)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2349 (
        .y(_T_1549),
        .a(io_rw_addr),
        .b(_WTEMP_222)
    );
    wire _T_1551;
    EQ_UNSIGNED #(.width(12)) u_eq_2350 (
        .y(_T_1551),
        .a(io_rw_addr),
        .b(12'hB08)
    );
    wire _T_1553;
    EQ_UNSIGNED #(.width(12)) u_eq_2351 (
        .y(_T_1553),
        .a(io_rw_addr),
        .b(12'hC08)
    );
    wire _T_1555;
    wire [11:0] _WTEMP_223;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2352 (
        .y(_WTEMP_223),
        .in(10'h329)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2353 (
        .y(_T_1555),
        .a(io_rw_addr),
        .b(_WTEMP_223)
    );
    wire _T_1557;
    EQ_UNSIGNED #(.width(12)) u_eq_2354 (
        .y(_T_1557),
        .a(io_rw_addr),
        .b(12'hB09)
    );
    wire _T_1559;
    EQ_UNSIGNED #(.width(12)) u_eq_2355 (
        .y(_T_1559),
        .a(io_rw_addr),
        .b(12'hC09)
    );
    wire _T_1561;
    wire [11:0] _WTEMP_224;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2356 (
        .y(_WTEMP_224),
        .in(10'h32A)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2357 (
        .y(_T_1561),
        .a(io_rw_addr),
        .b(_WTEMP_224)
    );
    wire _T_1563;
    EQ_UNSIGNED #(.width(12)) u_eq_2358 (
        .y(_T_1563),
        .a(io_rw_addr),
        .b(12'hB0A)
    );
    wire _T_1565;
    EQ_UNSIGNED #(.width(12)) u_eq_2359 (
        .y(_T_1565),
        .a(io_rw_addr),
        .b(12'hC0A)
    );
    wire _T_1567;
    wire [11:0] _WTEMP_225;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2360 (
        .y(_WTEMP_225),
        .in(10'h32B)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2361 (
        .y(_T_1567),
        .a(io_rw_addr),
        .b(_WTEMP_225)
    );
    wire _T_1569;
    EQ_UNSIGNED #(.width(12)) u_eq_2362 (
        .y(_T_1569),
        .a(io_rw_addr),
        .b(12'hB0B)
    );
    wire _T_1571;
    EQ_UNSIGNED #(.width(12)) u_eq_2363 (
        .y(_T_1571),
        .a(io_rw_addr),
        .b(12'hC0B)
    );
    wire _T_1573;
    wire [11:0] _WTEMP_226;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2364 (
        .y(_WTEMP_226),
        .in(10'h32C)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2365 (
        .y(_T_1573),
        .a(io_rw_addr),
        .b(_WTEMP_226)
    );
    wire _T_1575;
    EQ_UNSIGNED #(.width(12)) u_eq_2366 (
        .y(_T_1575),
        .a(io_rw_addr),
        .b(12'hB0C)
    );
    wire _T_1577;
    EQ_UNSIGNED #(.width(12)) u_eq_2367 (
        .y(_T_1577),
        .a(io_rw_addr),
        .b(12'hC0C)
    );
    wire _T_1579;
    wire [11:0] _WTEMP_227;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2368 (
        .y(_WTEMP_227),
        .in(10'h32D)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2369 (
        .y(_T_1579),
        .a(io_rw_addr),
        .b(_WTEMP_227)
    );
    wire _T_1581;
    EQ_UNSIGNED #(.width(12)) u_eq_2370 (
        .y(_T_1581),
        .a(io_rw_addr),
        .b(12'hB0D)
    );
    wire _T_1583;
    EQ_UNSIGNED #(.width(12)) u_eq_2371 (
        .y(_T_1583),
        .a(io_rw_addr),
        .b(12'hC0D)
    );
    wire _T_1585;
    wire [11:0] _WTEMP_228;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2372 (
        .y(_WTEMP_228),
        .in(10'h32E)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2373 (
        .y(_T_1585),
        .a(io_rw_addr),
        .b(_WTEMP_228)
    );
    wire _T_1587;
    EQ_UNSIGNED #(.width(12)) u_eq_2374 (
        .y(_T_1587),
        .a(io_rw_addr),
        .b(12'hB0E)
    );
    wire _T_1589;
    EQ_UNSIGNED #(.width(12)) u_eq_2375 (
        .y(_T_1589),
        .a(io_rw_addr),
        .b(12'hC0E)
    );
    wire _T_1591;
    wire [11:0] _WTEMP_229;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2376 (
        .y(_WTEMP_229),
        .in(10'h32F)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2377 (
        .y(_T_1591),
        .a(io_rw_addr),
        .b(_WTEMP_229)
    );
    wire _T_1593;
    EQ_UNSIGNED #(.width(12)) u_eq_2378 (
        .y(_T_1593),
        .a(io_rw_addr),
        .b(12'hB0F)
    );
    wire _T_1595;
    EQ_UNSIGNED #(.width(12)) u_eq_2379 (
        .y(_T_1595),
        .a(io_rw_addr),
        .b(12'hC0F)
    );
    wire _T_1597;
    wire [11:0] _WTEMP_230;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2380 (
        .y(_WTEMP_230),
        .in(10'h330)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2381 (
        .y(_T_1597),
        .a(io_rw_addr),
        .b(_WTEMP_230)
    );
    wire _T_1599;
    EQ_UNSIGNED #(.width(12)) u_eq_2382 (
        .y(_T_1599),
        .a(io_rw_addr),
        .b(12'hB10)
    );
    wire _T_1601;
    EQ_UNSIGNED #(.width(12)) u_eq_2383 (
        .y(_T_1601),
        .a(io_rw_addr),
        .b(12'hC10)
    );
    wire _T_1603;
    wire [11:0] _WTEMP_231;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2384 (
        .y(_WTEMP_231),
        .in(10'h331)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2385 (
        .y(_T_1603),
        .a(io_rw_addr),
        .b(_WTEMP_231)
    );
    wire _T_1605;
    EQ_UNSIGNED #(.width(12)) u_eq_2386 (
        .y(_T_1605),
        .a(io_rw_addr),
        .b(12'hB11)
    );
    wire _T_1607;
    EQ_UNSIGNED #(.width(12)) u_eq_2387 (
        .y(_T_1607),
        .a(io_rw_addr),
        .b(12'hC11)
    );
    wire _T_1609;
    wire [11:0] _WTEMP_232;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2388 (
        .y(_WTEMP_232),
        .in(10'h332)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2389 (
        .y(_T_1609),
        .a(io_rw_addr),
        .b(_WTEMP_232)
    );
    wire _T_1611;
    EQ_UNSIGNED #(.width(12)) u_eq_2390 (
        .y(_T_1611),
        .a(io_rw_addr),
        .b(12'hB12)
    );
    wire _T_1613;
    EQ_UNSIGNED #(.width(12)) u_eq_2391 (
        .y(_T_1613),
        .a(io_rw_addr),
        .b(12'hC12)
    );
    wire _T_1615;
    wire [11:0] _WTEMP_233;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2392 (
        .y(_WTEMP_233),
        .in(10'h333)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2393 (
        .y(_T_1615),
        .a(io_rw_addr),
        .b(_WTEMP_233)
    );
    wire _T_1617;
    EQ_UNSIGNED #(.width(12)) u_eq_2394 (
        .y(_T_1617),
        .a(io_rw_addr),
        .b(12'hB13)
    );
    wire _T_1619;
    EQ_UNSIGNED #(.width(12)) u_eq_2395 (
        .y(_T_1619),
        .a(io_rw_addr),
        .b(12'hC13)
    );
    wire _T_1621;
    wire [11:0] _WTEMP_234;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2396 (
        .y(_WTEMP_234),
        .in(10'h334)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2397 (
        .y(_T_1621),
        .a(io_rw_addr),
        .b(_WTEMP_234)
    );
    wire _T_1623;
    EQ_UNSIGNED #(.width(12)) u_eq_2398 (
        .y(_T_1623),
        .a(io_rw_addr),
        .b(12'hB14)
    );
    wire _T_1625;
    EQ_UNSIGNED #(.width(12)) u_eq_2399 (
        .y(_T_1625),
        .a(io_rw_addr),
        .b(12'hC14)
    );
    wire _T_1627;
    wire [11:0] _WTEMP_235;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2400 (
        .y(_WTEMP_235),
        .in(10'h335)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2401 (
        .y(_T_1627),
        .a(io_rw_addr),
        .b(_WTEMP_235)
    );
    wire _T_1629;
    EQ_UNSIGNED #(.width(12)) u_eq_2402 (
        .y(_T_1629),
        .a(io_rw_addr),
        .b(12'hB15)
    );
    wire _T_1631;
    EQ_UNSIGNED #(.width(12)) u_eq_2403 (
        .y(_T_1631),
        .a(io_rw_addr),
        .b(12'hC15)
    );
    wire _T_1633;
    wire [11:0] _WTEMP_236;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2404 (
        .y(_WTEMP_236),
        .in(10'h336)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2405 (
        .y(_T_1633),
        .a(io_rw_addr),
        .b(_WTEMP_236)
    );
    wire _T_1635;
    EQ_UNSIGNED #(.width(12)) u_eq_2406 (
        .y(_T_1635),
        .a(io_rw_addr),
        .b(12'hB16)
    );
    wire _T_1637;
    EQ_UNSIGNED #(.width(12)) u_eq_2407 (
        .y(_T_1637),
        .a(io_rw_addr),
        .b(12'hC16)
    );
    wire _T_1639;
    wire [11:0] _WTEMP_237;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2408 (
        .y(_WTEMP_237),
        .in(10'h337)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2409 (
        .y(_T_1639),
        .a(io_rw_addr),
        .b(_WTEMP_237)
    );
    wire _T_1641;
    EQ_UNSIGNED #(.width(12)) u_eq_2410 (
        .y(_T_1641),
        .a(io_rw_addr),
        .b(12'hB17)
    );
    wire _T_1643;
    EQ_UNSIGNED #(.width(12)) u_eq_2411 (
        .y(_T_1643),
        .a(io_rw_addr),
        .b(12'hC17)
    );
    wire _T_1645;
    wire [11:0] _WTEMP_238;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2412 (
        .y(_WTEMP_238),
        .in(10'h338)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2413 (
        .y(_T_1645),
        .a(io_rw_addr),
        .b(_WTEMP_238)
    );
    wire _T_1647;
    EQ_UNSIGNED #(.width(12)) u_eq_2414 (
        .y(_T_1647),
        .a(io_rw_addr),
        .b(12'hB18)
    );
    wire _T_1649;
    EQ_UNSIGNED #(.width(12)) u_eq_2415 (
        .y(_T_1649),
        .a(io_rw_addr),
        .b(12'hC18)
    );
    wire _T_1651;
    wire [11:0] _WTEMP_239;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2416 (
        .y(_WTEMP_239),
        .in(10'h339)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2417 (
        .y(_T_1651),
        .a(io_rw_addr),
        .b(_WTEMP_239)
    );
    wire _T_1653;
    EQ_UNSIGNED #(.width(12)) u_eq_2418 (
        .y(_T_1653),
        .a(io_rw_addr),
        .b(12'hB19)
    );
    wire _T_1655;
    EQ_UNSIGNED #(.width(12)) u_eq_2419 (
        .y(_T_1655),
        .a(io_rw_addr),
        .b(12'hC19)
    );
    wire _T_1657;
    wire [11:0] _WTEMP_240;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2420 (
        .y(_WTEMP_240),
        .in(10'h33A)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2421 (
        .y(_T_1657),
        .a(io_rw_addr),
        .b(_WTEMP_240)
    );
    wire _T_1659;
    EQ_UNSIGNED #(.width(12)) u_eq_2422 (
        .y(_T_1659),
        .a(io_rw_addr),
        .b(12'hB1A)
    );
    wire _T_1661;
    EQ_UNSIGNED #(.width(12)) u_eq_2423 (
        .y(_T_1661),
        .a(io_rw_addr),
        .b(12'hC1A)
    );
    wire _T_1663;
    wire [11:0] _WTEMP_241;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2424 (
        .y(_WTEMP_241),
        .in(10'h33B)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2425 (
        .y(_T_1663),
        .a(io_rw_addr),
        .b(_WTEMP_241)
    );
    wire _T_1665;
    EQ_UNSIGNED #(.width(12)) u_eq_2426 (
        .y(_T_1665),
        .a(io_rw_addr),
        .b(12'hB1B)
    );
    wire _T_1667;
    EQ_UNSIGNED #(.width(12)) u_eq_2427 (
        .y(_T_1667),
        .a(io_rw_addr),
        .b(12'hC1B)
    );
    wire _T_1669;
    wire [11:0] _WTEMP_242;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2428 (
        .y(_WTEMP_242),
        .in(10'h33C)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2429 (
        .y(_T_1669),
        .a(io_rw_addr),
        .b(_WTEMP_242)
    );
    wire _T_1671;
    EQ_UNSIGNED #(.width(12)) u_eq_2430 (
        .y(_T_1671),
        .a(io_rw_addr),
        .b(12'hB1C)
    );
    wire _T_1673;
    EQ_UNSIGNED #(.width(12)) u_eq_2431 (
        .y(_T_1673),
        .a(io_rw_addr),
        .b(12'hC1C)
    );
    wire _T_1675;
    wire [11:0] _WTEMP_243;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2432 (
        .y(_WTEMP_243),
        .in(10'h33D)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2433 (
        .y(_T_1675),
        .a(io_rw_addr),
        .b(_WTEMP_243)
    );
    wire _T_1677;
    EQ_UNSIGNED #(.width(12)) u_eq_2434 (
        .y(_T_1677),
        .a(io_rw_addr),
        .b(12'hB1D)
    );
    wire _T_1679;
    EQ_UNSIGNED #(.width(12)) u_eq_2435 (
        .y(_T_1679),
        .a(io_rw_addr),
        .b(12'hC1D)
    );
    wire _T_1681;
    wire [11:0] _WTEMP_244;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2436 (
        .y(_WTEMP_244),
        .in(10'h33E)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2437 (
        .y(_T_1681),
        .a(io_rw_addr),
        .b(_WTEMP_244)
    );
    wire _T_1683;
    EQ_UNSIGNED #(.width(12)) u_eq_2438 (
        .y(_T_1683),
        .a(io_rw_addr),
        .b(12'hB1E)
    );
    wire _T_1685;
    EQ_UNSIGNED #(.width(12)) u_eq_2439 (
        .y(_T_1685),
        .a(io_rw_addr),
        .b(12'hC1E)
    );
    wire _T_1687;
    wire [11:0] _WTEMP_245;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2440 (
        .y(_WTEMP_245),
        .in(10'h33F)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2441 (
        .y(_T_1687),
        .a(io_rw_addr),
        .b(_WTEMP_245)
    );
    wire _T_1689;
    EQ_UNSIGNED #(.width(12)) u_eq_2442 (
        .y(_T_1689),
        .a(io_rw_addr),
        .b(12'hB1F)
    );
    wire _T_1691;
    EQ_UNSIGNED #(.width(12)) u_eq_2443 (
        .y(_T_1691),
        .a(io_rw_addr),
        .b(12'hC1F)
    );
    wire _T_1693;
    wire [11:0] _WTEMP_246;
    PAD_UNSIGNED #(.width(9), .n(12)) u_pad_2444 (
        .y(_WTEMP_246),
        .in(9'h100)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2445 (
        .y(_T_1693),
        .a(io_rw_addr),
        .b(_WTEMP_246)
    );
    wire _T_1695;
    wire [11:0] _WTEMP_247;
    PAD_UNSIGNED #(.width(9), .n(12)) u_pad_2446 (
        .y(_WTEMP_247),
        .in(9'h144)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2447 (
        .y(_T_1695),
        .a(io_rw_addr),
        .b(_WTEMP_247)
    );
    wire _T_1697;
    wire [11:0] _WTEMP_248;
    PAD_UNSIGNED #(.width(9), .n(12)) u_pad_2448 (
        .y(_WTEMP_248),
        .in(9'h104)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2449 (
        .y(_T_1697),
        .a(io_rw_addr),
        .b(_WTEMP_248)
    );
    wire _T_1699;
    wire [11:0] _WTEMP_249;
    PAD_UNSIGNED #(.width(9), .n(12)) u_pad_2450 (
        .y(_WTEMP_249),
        .in(9'h140)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2451 (
        .y(_T_1699),
        .a(io_rw_addr),
        .b(_WTEMP_249)
    );
    wire _T_1701;
    wire [11:0] _WTEMP_250;
    PAD_UNSIGNED #(.width(9), .n(12)) u_pad_2452 (
        .y(_WTEMP_250),
        .in(9'h142)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2453 (
        .y(_T_1701),
        .a(io_rw_addr),
        .b(_WTEMP_250)
    );
    wire _T_1703;
    wire [11:0] _WTEMP_251;
    PAD_UNSIGNED #(.width(9), .n(12)) u_pad_2454 (
        .y(_WTEMP_251),
        .in(9'h143)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2455 (
        .y(_T_1703),
        .a(io_rw_addr),
        .b(_WTEMP_251)
    );
    wire _T_1705;
    wire [11:0] _WTEMP_252;
    PAD_UNSIGNED #(.width(9), .n(12)) u_pad_2456 (
        .y(_WTEMP_252),
        .in(9'h180)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2457 (
        .y(_T_1705),
        .a(io_rw_addr),
        .b(_WTEMP_252)
    );
    wire _T_1707;
    wire [11:0] _WTEMP_253;
    PAD_UNSIGNED #(.width(9), .n(12)) u_pad_2458 (
        .y(_WTEMP_253),
        .in(9'h141)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2459 (
        .y(_T_1707),
        .a(io_rw_addr),
        .b(_WTEMP_253)
    );
    wire _T_1709;
    wire [11:0] _WTEMP_254;
    PAD_UNSIGNED #(.width(9), .n(12)) u_pad_2460 (
        .y(_WTEMP_254),
        .in(9'h105)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2461 (
        .y(_T_1709),
        .a(io_rw_addr),
        .b(_WTEMP_254)
    );
    wire _T_1711;
    wire [11:0] _WTEMP_255;
    PAD_UNSIGNED #(.width(9), .n(12)) u_pad_2462 (
        .y(_WTEMP_255),
        .in(9'h106)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2463 (
        .y(_T_1711),
        .a(io_rw_addr),
        .b(_WTEMP_255)
    );
    wire _T_1713;
    wire [11:0] _WTEMP_256;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2464 (
        .y(_WTEMP_256),
        .in(10'h306)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2465 (
        .y(_T_1713),
        .a(io_rw_addr),
        .b(_WTEMP_256)
    );
    wire _T_1715;
    EQ_UNSIGNED #(.width(12)) u_eq_2466 (
        .y(_T_1715),
        .a(io_rw_addr),
        .b(12'hC00)
    );
    wire _T_1717;
    EQ_UNSIGNED #(.width(12)) u_eq_2467 (
        .y(_T_1717),
        .a(io_rw_addr),
        .b(12'hC02)
    );
    wire _T_1720;
    EQ_UNSIGNED #(.width(3)) u_eq_2468 (
        .y(_T_1720),
        .a(io_rw_cmd),
        .b(3'h2)
    );
    wire _T_1721;
    EQ_UNSIGNED #(.width(3)) u_eq_2469 (
        .y(_T_1721),
        .a(io_rw_cmd),
        .b(3'h3)
    );
    wire _T_1722;
    BITWISEOR #(.width(1)) bitwiseor_2470 (
        .y(_T_1722),
        .a(_T_1720),
        .b(_T_1721)
    );
    wire [63:0] _T_1724;
    wire [63:0] _WTEMP_257;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_2471 (
        .y(_WTEMP_257),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_2472 (
        .y(_T_1724),
        .sel(_T_1722),
        .a(io_rw_rdata),
        .b(_WTEMP_257)
    );
    wire [63:0] _T_1725;
    BITWISEOR #(.width(64)) bitwiseor_2473 (
        .y(_T_1725),
        .a(_T_1724),
        .b(io_rw_wdata)
    );
    wire _T_1727;
    EQ_UNSIGNED #(.width(3)) u_eq_2474 (
        .y(_T_1727),
        .a(io_rw_cmd),
        .b(3'h3)
    );
    wire [63:0] _T_1729;
    wire [63:0] _WTEMP_258;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_2475 (
        .y(_WTEMP_258),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_2476 (
        .y(_T_1729),
        .sel(_T_1727),
        .a(io_rw_wdata),
        .b(_WTEMP_258)
    );
    wire [63:0] _T_1730;
    BITWISENOT #(.width(64)) bitwisenot_2477 (
        .y(_T_1730),
        .in(_T_1729)
    );
    wire [63:0] wdata;
    BITWISEAND #(.width(64)) bitwiseand_2478 (
        .y(wdata),
        .a(_T_1725),
        .b(_T_1730)
    );
    wire system_insn;
    EQ_UNSIGNED #(.width(3)) u_eq_2479 (
        .y(system_insn),
        .a(io_rw_cmd),
        .b(3'h4)
    );
    wire [2:0] _T_1733;
    BITS #(.width(12), .high(2), .low(0)) bits_2480 (
        .y(_T_1733),
        .in(io_rw_addr)
    );
    wire [7:0] opcode;
    DSHL_UNSIGNED #(.width_in(1), .width_n(3)) u_dshl_2481 (
        .y(opcode),
        .in(1'h1),
        .n(_T_1733)
    );
    wire insn_rs2;
    BITS #(.width(12), .high(5), .low(5)) bits_2482 (
        .y(insn_rs2),
        .in(io_rw_addr)
    );
    wire _T_1735;
    EQ_UNSIGNED #(.width(1)) u_eq_2483 (
        .y(_T_1735),
        .a(insn_rs2),
        .b(1'h0)
    );
    wire _T_1736;
    BITWISEAND #(.width(1)) bitwiseand_2484 (
        .y(_T_1736),
        .a(system_insn),
        .b(_T_1735)
    );
    wire _T_1737;
    BITS #(.width(8), .high(0), .low(0)) bits_2485 (
        .y(_T_1737),
        .in(opcode)
    );
    wire insn_call;
    BITWISEAND #(.width(1)) bitwiseand_2486 (
        .y(insn_call),
        .a(_T_1736),
        .b(_T_1737)
    );
    wire _T_1738;
    BITS #(.width(8), .high(1), .low(1)) bits_2487 (
        .y(_T_1738),
        .in(opcode)
    );
    wire insn_break;
    BITWISEAND #(.width(1)) bitwiseand_2488 (
        .y(insn_break),
        .a(system_insn),
        .b(_T_1738)
    );
    wire _T_1739;
    BITS #(.width(8), .high(2), .low(2)) bits_2489 (
        .y(_T_1739),
        .in(opcode)
    );
    wire insn_ret;
    BITWISEAND #(.width(1)) bitwiseand_2490 (
        .y(insn_ret),
        .a(system_insn),
        .b(_T_1739)
    );
    wire _T_1740;
    BITS #(.width(8), .high(5), .low(5)) bits_2491 (
        .y(_T_1740),
        .in(opcode)
    );
    wire insn_wfi;
    BITWISEAND #(.width(1)) bitwiseand_2492 (
        .y(insn_wfi),
        .a(system_insn),
        .b(_T_1740)
    );
    wire insn_sfence_vma;
    BITWISEAND #(.width(1)) bitwiseand_2493 (
        .y(insn_sfence_vma),
        .a(system_insn),
        .b(insn_rs2)
    );
    wire _T_1743;
    wire [2:0] _WTEMP_259;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_2494 (
        .y(_WTEMP_259),
        .in(1'h1)
    );
    GT_UNSIGNED #(.width(3)) u_gt_2495 (
        .y(_T_1743),
        .a(effective_prv),
        .b(_WTEMP_259)
    );
    wire _T_1744;
    BITWISEOR #(.width(1)) bitwiseor_2496 (
        .y(_T_1744),
        .a(1'h0),
        .b(_T_1743)
    );
    wire _T_1746;
    EQ_UNSIGNED #(.width(1)) u_eq_2497 (
        .y(_T_1746),
        .a(_reg_mstatus_tw__q),
        .b(1'h0)
    );
    wire allow_wfi;
    BITWISEOR #(.width(1)) bitwiseor_2498 (
        .y(allow_wfi),
        .a(_T_1744),
        .b(_T_1746)
    );
    wire _T_1749;
    wire [2:0] _WTEMP_260;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_2499 (
        .y(_WTEMP_260),
        .in(1'h1)
    );
    GT_UNSIGNED #(.width(3)) u_gt_2500 (
        .y(_T_1749),
        .a(effective_prv),
        .b(_WTEMP_260)
    );
    wire _T_1750;
    BITWISEOR #(.width(1)) bitwiseor_2501 (
        .y(_T_1750),
        .a(1'h0),
        .b(_T_1749)
    );
    wire _T_1752;
    EQ_UNSIGNED #(.width(1)) u_eq_2502 (
        .y(_T_1752),
        .a(_reg_mstatus_tvm__q),
        .b(1'h0)
    );
    wire allow_sfence_vma;
    BITWISEOR #(.width(1)) bitwiseor_2503 (
        .y(allow_sfence_vma),
        .a(_T_1750),
        .b(_T_1752)
    );
    wire _T_1755;
    wire [2:0] _WTEMP_261;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_2504 (
        .y(_WTEMP_261),
        .in(1'h1)
    );
    GT_UNSIGNED #(.width(3)) u_gt_2505 (
        .y(_T_1755),
        .a(effective_prv),
        .b(_WTEMP_261)
    );
    wire _T_1756;
    BITWISEOR #(.width(1)) bitwiseor_2506 (
        .y(_T_1756),
        .a(1'h0),
        .b(_T_1755)
    );
    wire _T_1758;
    EQ_UNSIGNED #(.width(1)) u_eq_2507 (
        .y(_T_1758),
        .a(_reg_mstatus_tsr__q),
        .b(1'h0)
    );
    wire allow_sret;
    BITWISEOR #(.width(1)) bitwiseor_2508 (
        .y(allow_sret),
        .a(_T_1756),
        .b(_T_1758)
    );
    wire _T_1760;
    wire [1:0] _WTEMP_262;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2509 (
        .y(_WTEMP_262),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(2)) u_eq_2510 (
        .y(_T_1760),
        .a(io_status_fs),
        .b(_WTEMP_262)
    );
    wire _T_1761;
    BITS #(.width(64), .high(5), .low(5)) bits_2511 (
        .y(_T_1761),
        .in(_reg_misa__q)
    );
    wire _T_1763;
    EQ_UNSIGNED #(.width(1)) u_eq_2512 (
        .y(_T_1763),
        .a(_T_1761),
        .b(1'h0)
    );
    wire _T_1764;
    BITWISEOR #(.width(1)) bitwiseor_2513 (
        .y(_T_1764),
        .a(_T_1760),
        .b(_T_1763)
    );
    wire _T_1766;
    wire [1:0] _WTEMP_263;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2514 (
        .y(_WTEMP_263),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(2)) u_eq_2515 (
        .y(_T_1766),
        .a(io_status_xs),
        .b(_WTEMP_263)
    );
    wire _T_1767;
    BITS #(.width(64), .high(23), .low(23)) bits_2516 (
        .y(_T_1767),
        .in(_reg_misa__q)
    );
    wire _T_1769;
    EQ_UNSIGNED #(.width(1)) u_eq_2517 (
        .y(_T_1769),
        .a(_T_1767),
        .b(1'h0)
    );
    wire _T_1770;
    BITWISEOR #(.width(1)) bitwiseor_2518 (
        .y(_T_1770),
        .a(_T_1766),
        .b(_T_1769)
    );
    wire [1:0] _T_1771;
    BITS #(.width(12), .high(9), .low(8)) bits_2519 (
        .y(_T_1771),
        .in(io_decode_csr)
    );
    wire _T_1772;
    wire [2:0] _WTEMP_264;
    PAD_UNSIGNED #(.width(2), .n(3)) u_pad_2520 (
        .y(_WTEMP_264),
        .in(_T_1771)
    );
    LT_UNSIGNED #(.width(3)) u_lt_2521 (
        .y(_T_1772),
        .a(effective_prv),
        .b(_WTEMP_264)
    );
    wire _T_1774;
    wire [11:0] _WTEMP_265;
    PAD_UNSIGNED #(.width(11), .n(12)) u_pad_2522 (
        .y(_WTEMP_265),
        .in(11'h7A0)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2523 (
        .y(_T_1774),
        .a(io_decode_csr),
        .b(_WTEMP_265)
    );
    wire _T_1776;
    wire [11:0] _WTEMP_266;
    PAD_UNSIGNED #(.width(11), .n(12)) u_pad_2524 (
        .y(_WTEMP_266),
        .in(11'h7A1)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2525 (
        .y(_T_1776),
        .a(io_decode_csr),
        .b(_WTEMP_266)
    );
    wire _T_1778;
    wire [11:0] _WTEMP_267;
    PAD_UNSIGNED #(.width(11), .n(12)) u_pad_2526 (
        .y(_WTEMP_267),
        .in(11'h7A2)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2527 (
        .y(_T_1778),
        .a(io_decode_csr),
        .b(_WTEMP_267)
    );
    wire _T_1780;
    EQ_UNSIGNED #(.width(12)) u_eq_2528 (
        .y(_T_1780),
        .a(io_decode_csr),
        .b(12'hF13)
    );
    wire _T_1782;
    EQ_UNSIGNED #(.width(12)) u_eq_2529 (
        .y(_T_1782),
        .a(io_decode_csr),
        .b(12'hF12)
    );
    wire _T_1784;
    EQ_UNSIGNED #(.width(12)) u_eq_2530 (
        .y(_T_1784),
        .a(io_decode_csr),
        .b(12'hF11)
    );
    wire _T_1786;
    EQ_UNSIGNED #(.width(12)) u_eq_2531 (
        .y(_T_1786),
        .a(io_decode_csr),
        .b(12'hB00)
    );
    wire _T_1788;
    EQ_UNSIGNED #(.width(12)) u_eq_2532 (
        .y(_T_1788),
        .a(io_decode_csr),
        .b(12'hB02)
    );
    wire _T_1790;
    wire [11:0] _WTEMP_268;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2533 (
        .y(_WTEMP_268),
        .in(10'h301)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2534 (
        .y(_T_1790),
        .a(io_decode_csr),
        .b(_WTEMP_268)
    );
    wire _T_1792;
    wire [11:0] _WTEMP_269;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2535 (
        .y(_WTEMP_269),
        .in(10'h300)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2536 (
        .y(_T_1792),
        .a(io_decode_csr),
        .b(_WTEMP_269)
    );
    wire _T_1794;
    wire [11:0] _WTEMP_270;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2537 (
        .y(_WTEMP_270),
        .in(10'h305)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2538 (
        .y(_T_1794),
        .a(io_decode_csr),
        .b(_WTEMP_270)
    );
    wire _T_1796;
    wire [11:0] _WTEMP_271;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2539 (
        .y(_WTEMP_271),
        .in(10'h344)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2540 (
        .y(_T_1796),
        .a(io_decode_csr),
        .b(_WTEMP_271)
    );
    wire _T_1798;
    wire [11:0] _WTEMP_272;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2541 (
        .y(_WTEMP_272),
        .in(10'h304)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2542 (
        .y(_T_1798),
        .a(io_decode_csr),
        .b(_WTEMP_272)
    );
    wire _T_1800;
    wire [11:0] _WTEMP_273;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2543 (
        .y(_WTEMP_273),
        .in(10'h303)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2544 (
        .y(_T_1800),
        .a(io_decode_csr),
        .b(_WTEMP_273)
    );
    wire _T_1802;
    wire [11:0] _WTEMP_274;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2545 (
        .y(_WTEMP_274),
        .in(10'h302)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2546 (
        .y(_T_1802),
        .a(io_decode_csr),
        .b(_WTEMP_274)
    );
    wire _T_1804;
    wire [11:0] _WTEMP_275;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2547 (
        .y(_WTEMP_275),
        .in(10'h340)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2548 (
        .y(_T_1804),
        .a(io_decode_csr),
        .b(_WTEMP_275)
    );
    wire _T_1806;
    wire [11:0] _WTEMP_276;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2549 (
        .y(_WTEMP_276),
        .in(10'h341)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2550 (
        .y(_T_1806),
        .a(io_decode_csr),
        .b(_WTEMP_276)
    );
    wire _T_1808;
    wire [11:0] _WTEMP_277;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2551 (
        .y(_WTEMP_277),
        .in(10'h343)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2552 (
        .y(_T_1808),
        .a(io_decode_csr),
        .b(_WTEMP_277)
    );
    wire _T_1810;
    wire [11:0] _WTEMP_278;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2553 (
        .y(_WTEMP_278),
        .in(10'h342)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2554 (
        .y(_T_1810),
        .a(io_decode_csr),
        .b(_WTEMP_278)
    );
    wire _T_1812;
    EQ_UNSIGNED #(.width(12)) u_eq_2555 (
        .y(_T_1812),
        .a(io_decode_csr),
        .b(12'hF14)
    );
    wire _T_1814;
    wire [11:0] _WTEMP_279;
    PAD_UNSIGNED #(.width(11), .n(12)) u_pad_2556 (
        .y(_WTEMP_279),
        .in(11'h7B0)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2557 (
        .y(_T_1814),
        .a(io_decode_csr),
        .b(_WTEMP_279)
    );
    wire _T_1816;
    wire [11:0] _WTEMP_280;
    PAD_UNSIGNED #(.width(11), .n(12)) u_pad_2558 (
        .y(_WTEMP_280),
        .in(11'h7B1)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2559 (
        .y(_T_1816),
        .a(io_decode_csr),
        .b(_WTEMP_280)
    );
    wire _T_1818;
    wire [11:0] _WTEMP_281;
    PAD_UNSIGNED #(.width(11), .n(12)) u_pad_2560 (
        .y(_WTEMP_281),
        .in(11'h7B2)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2561 (
        .y(_T_1818),
        .a(io_decode_csr),
        .b(_WTEMP_281)
    );
    wire _T_1820;
    wire [11:0] _WTEMP_282;
    PAD_UNSIGNED #(.width(1), .n(12)) u_pad_2562 (
        .y(_WTEMP_282),
        .in(1'h1)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2563 (
        .y(_T_1820),
        .a(io_decode_csr),
        .b(_WTEMP_282)
    );
    wire _T_1822;
    wire [11:0] _WTEMP_283;
    PAD_UNSIGNED #(.width(2), .n(12)) u_pad_2564 (
        .y(_WTEMP_283),
        .in(2'h2)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2565 (
        .y(_T_1822),
        .a(io_decode_csr),
        .b(_WTEMP_283)
    );
    wire _T_1824;
    wire [11:0] _WTEMP_284;
    PAD_UNSIGNED #(.width(2), .n(12)) u_pad_2566 (
        .y(_WTEMP_284),
        .in(2'h3)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2567 (
        .y(_T_1824),
        .a(io_decode_csr),
        .b(_WTEMP_284)
    );
    wire _T_1826;
    wire [11:0] _WTEMP_285;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2568 (
        .y(_WTEMP_285),
        .in(10'h323)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2569 (
        .y(_T_1826),
        .a(io_decode_csr),
        .b(_WTEMP_285)
    );
    wire _T_1828;
    EQ_UNSIGNED #(.width(12)) u_eq_2570 (
        .y(_T_1828),
        .a(io_decode_csr),
        .b(12'hB03)
    );
    wire _T_1830;
    EQ_UNSIGNED #(.width(12)) u_eq_2571 (
        .y(_T_1830),
        .a(io_decode_csr),
        .b(12'hC03)
    );
    wire _T_1832;
    wire [11:0] _WTEMP_286;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2572 (
        .y(_WTEMP_286),
        .in(10'h324)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2573 (
        .y(_T_1832),
        .a(io_decode_csr),
        .b(_WTEMP_286)
    );
    wire _T_1834;
    EQ_UNSIGNED #(.width(12)) u_eq_2574 (
        .y(_T_1834),
        .a(io_decode_csr),
        .b(12'hB04)
    );
    wire _T_1836;
    EQ_UNSIGNED #(.width(12)) u_eq_2575 (
        .y(_T_1836),
        .a(io_decode_csr),
        .b(12'hC04)
    );
    wire _T_1838;
    wire [11:0] _WTEMP_287;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2576 (
        .y(_WTEMP_287),
        .in(10'h325)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2577 (
        .y(_T_1838),
        .a(io_decode_csr),
        .b(_WTEMP_287)
    );
    wire _T_1840;
    EQ_UNSIGNED #(.width(12)) u_eq_2578 (
        .y(_T_1840),
        .a(io_decode_csr),
        .b(12'hB05)
    );
    wire _T_1842;
    EQ_UNSIGNED #(.width(12)) u_eq_2579 (
        .y(_T_1842),
        .a(io_decode_csr),
        .b(12'hC05)
    );
    wire _T_1844;
    wire [11:0] _WTEMP_288;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2580 (
        .y(_WTEMP_288),
        .in(10'h326)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2581 (
        .y(_T_1844),
        .a(io_decode_csr),
        .b(_WTEMP_288)
    );
    wire _T_1846;
    EQ_UNSIGNED #(.width(12)) u_eq_2582 (
        .y(_T_1846),
        .a(io_decode_csr),
        .b(12'hB06)
    );
    wire _T_1848;
    EQ_UNSIGNED #(.width(12)) u_eq_2583 (
        .y(_T_1848),
        .a(io_decode_csr),
        .b(12'hC06)
    );
    wire _T_1850;
    wire [11:0] _WTEMP_289;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2584 (
        .y(_WTEMP_289),
        .in(10'h327)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2585 (
        .y(_T_1850),
        .a(io_decode_csr),
        .b(_WTEMP_289)
    );
    wire _T_1852;
    EQ_UNSIGNED #(.width(12)) u_eq_2586 (
        .y(_T_1852),
        .a(io_decode_csr),
        .b(12'hB07)
    );
    wire _T_1854;
    EQ_UNSIGNED #(.width(12)) u_eq_2587 (
        .y(_T_1854),
        .a(io_decode_csr),
        .b(12'hC07)
    );
    wire _T_1856;
    wire [11:0] _WTEMP_290;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2588 (
        .y(_WTEMP_290),
        .in(10'h328)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2589 (
        .y(_T_1856),
        .a(io_decode_csr),
        .b(_WTEMP_290)
    );
    wire _T_1858;
    EQ_UNSIGNED #(.width(12)) u_eq_2590 (
        .y(_T_1858),
        .a(io_decode_csr),
        .b(12'hB08)
    );
    wire _T_1860;
    EQ_UNSIGNED #(.width(12)) u_eq_2591 (
        .y(_T_1860),
        .a(io_decode_csr),
        .b(12'hC08)
    );
    wire _T_1862;
    wire [11:0] _WTEMP_291;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2592 (
        .y(_WTEMP_291),
        .in(10'h329)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2593 (
        .y(_T_1862),
        .a(io_decode_csr),
        .b(_WTEMP_291)
    );
    wire _T_1864;
    EQ_UNSIGNED #(.width(12)) u_eq_2594 (
        .y(_T_1864),
        .a(io_decode_csr),
        .b(12'hB09)
    );
    wire _T_1866;
    EQ_UNSIGNED #(.width(12)) u_eq_2595 (
        .y(_T_1866),
        .a(io_decode_csr),
        .b(12'hC09)
    );
    wire _T_1868;
    wire [11:0] _WTEMP_292;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2596 (
        .y(_WTEMP_292),
        .in(10'h32A)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2597 (
        .y(_T_1868),
        .a(io_decode_csr),
        .b(_WTEMP_292)
    );
    wire _T_1870;
    EQ_UNSIGNED #(.width(12)) u_eq_2598 (
        .y(_T_1870),
        .a(io_decode_csr),
        .b(12'hB0A)
    );
    wire _T_1872;
    EQ_UNSIGNED #(.width(12)) u_eq_2599 (
        .y(_T_1872),
        .a(io_decode_csr),
        .b(12'hC0A)
    );
    wire _T_1874;
    wire [11:0] _WTEMP_293;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2600 (
        .y(_WTEMP_293),
        .in(10'h32B)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2601 (
        .y(_T_1874),
        .a(io_decode_csr),
        .b(_WTEMP_293)
    );
    wire _T_1876;
    EQ_UNSIGNED #(.width(12)) u_eq_2602 (
        .y(_T_1876),
        .a(io_decode_csr),
        .b(12'hB0B)
    );
    wire _T_1878;
    EQ_UNSIGNED #(.width(12)) u_eq_2603 (
        .y(_T_1878),
        .a(io_decode_csr),
        .b(12'hC0B)
    );
    wire _T_1880;
    wire [11:0] _WTEMP_294;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2604 (
        .y(_WTEMP_294),
        .in(10'h32C)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2605 (
        .y(_T_1880),
        .a(io_decode_csr),
        .b(_WTEMP_294)
    );
    wire _T_1882;
    EQ_UNSIGNED #(.width(12)) u_eq_2606 (
        .y(_T_1882),
        .a(io_decode_csr),
        .b(12'hB0C)
    );
    wire _T_1884;
    EQ_UNSIGNED #(.width(12)) u_eq_2607 (
        .y(_T_1884),
        .a(io_decode_csr),
        .b(12'hC0C)
    );
    wire _T_1886;
    wire [11:0] _WTEMP_295;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2608 (
        .y(_WTEMP_295),
        .in(10'h32D)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2609 (
        .y(_T_1886),
        .a(io_decode_csr),
        .b(_WTEMP_295)
    );
    wire _T_1888;
    EQ_UNSIGNED #(.width(12)) u_eq_2610 (
        .y(_T_1888),
        .a(io_decode_csr),
        .b(12'hB0D)
    );
    wire _T_1890;
    EQ_UNSIGNED #(.width(12)) u_eq_2611 (
        .y(_T_1890),
        .a(io_decode_csr),
        .b(12'hC0D)
    );
    wire _T_1892;
    wire [11:0] _WTEMP_296;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2612 (
        .y(_WTEMP_296),
        .in(10'h32E)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2613 (
        .y(_T_1892),
        .a(io_decode_csr),
        .b(_WTEMP_296)
    );
    wire _T_1894;
    EQ_UNSIGNED #(.width(12)) u_eq_2614 (
        .y(_T_1894),
        .a(io_decode_csr),
        .b(12'hB0E)
    );
    wire _T_1896;
    EQ_UNSIGNED #(.width(12)) u_eq_2615 (
        .y(_T_1896),
        .a(io_decode_csr),
        .b(12'hC0E)
    );
    wire _T_1898;
    wire [11:0] _WTEMP_297;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2616 (
        .y(_WTEMP_297),
        .in(10'h32F)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2617 (
        .y(_T_1898),
        .a(io_decode_csr),
        .b(_WTEMP_297)
    );
    wire _T_1900;
    EQ_UNSIGNED #(.width(12)) u_eq_2618 (
        .y(_T_1900),
        .a(io_decode_csr),
        .b(12'hB0F)
    );
    wire _T_1902;
    EQ_UNSIGNED #(.width(12)) u_eq_2619 (
        .y(_T_1902),
        .a(io_decode_csr),
        .b(12'hC0F)
    );
    wire _T_1904;
    wire [11:0] _WTEMP_298;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2620 (
        .y(_WTEMP_298),
        .in(10'h330)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2621 (
        .y(_T_1904),
        .a(io_decode_csr),
        .b(_WTEMP_298)
    );
    wire _T_1906;
    EQ_UNSIGNED #(.width(12)) u_eq_2622 (
        .y(_T_1906),
        .a(io_decode_csr),
        .b(12'hB10)
    );
    wire _T_1908;
    EQ_UNSIGNED #(.width(12)) u_eq_2623 (
        .y(_T_1908),
        .a(io_decode_csr),
        .b(12'hC10)
    );
    wire _T_1910;
    wire [11:0] _WTEMP_299;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2624 (
        .y(_WTEMP_299),
        .in(10'h331)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2625 (
        .y(_T_1910),
        .a(io_decode_csr),
        .b(_WTEMP_299)
    );
    wire _T_1912;
    EQ_UNSIGNED #(.width(12)) u_eq_2626 (
        .y(_T_1912),
        .a(io_decode_csr),
        .b(12'hB11)
    );
    wire _T_1914;
    EQ_UNSIGNED #(.width(12)) u_eq_2627 (
        .y(_T_1914),
        .a(io_decode_csr),
        .b(12'hC11)
    );
    wire _T_1916;
    wire [11:0] _WTEMP_300;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2628 (
        .y(_WTEMP_300),
        .in(10'h332)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2629 (
        .y(_T_1916),
        .a(io_decode_csr),
        .b(_WTEMP_300)
    );
    wire _T_1918;
    EQ_UNSIGNED #(.width(12)) u_eq_2630 (
        .y(_T_1918),
        .a(io_decode_csr),
        .b(12'hB12)
    );
    wire _T_1920;
    EQ_UNSIGNED #(.width(12)) u_eq_2631 (
        .y(_T_1920),
        .a(io_decode_csr),
        .b(12'hC12)
    );
    wire _T_1922;
    wire [11:0] _WTEMP_301;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2632 (
        .y(_WTEMP_301),
        .in(10'h333)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2633 (
        .y(_T_1922),
        .a(io_decode_csr),
        .b(_WTEMP_301)
    );
    wire _T_1924;
    EQ_UNSIGNED #(.width(12)) u_eq_2634 (
        .y(_T_1924),
        .a(io_decode_csr),
        .b(12'hB13)
    );
    wire _T_1926;
    EQ_UNSIGNED #(.width(12)) u_eq_2635 (
        .y(_T_1926),
        .a(io_decode_csr),
        .b(12'hC13)
    );
    wire _T_1928;
    wire [11:0] _WTEMP_302;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2636 (
        .y(_WTEMP_302),
        .in(10'h334)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2637 (
        .y(_T_1928),
        .a(io_decode_csr),
        .b(_WTEMP_302)
    );
    wire _T_1930;
    EQ_UNSIGNED #(.width(12)) u_eq_2638 (
        .y(_T_1930),
        .a(io_decode_csr),
        .b(12'hB14)
    );
    wire _T_1932;
    EQ_UNSIGNED #(.width(12)) u_eq_2639 (
        .y(_T_1932),
        .a(io_decode_csr),
        .b(12'hC14)
    );
    wire _T_1934;
    wire [11:0] _WTEMP_303;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2640 (
        .y(_WTEMP_303),
        .in(10'h335)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2641 (
        .y(_T_1934),
        .a(io_decode_csr),
        .b(_WTEMP_303)
    );
    wire _T_1936;
    EQ_UNSIGNED #(.width(12)) u_eq_2642 (
        .y(_T_1936),
        .a(io_decode_csr),
        .b(12'hB15)
    );
    wire _T_1938;
    EQ_UNSIGNED #(.width(12)) u_eq_2643 (
        .y(_T_1938),
        .a(io_decode_csr),
        .b(12'hC15)
    );
    wire _T_1940;
    wire [11:0] _WTEMP_304;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2644 (
        .y(_WTEMP_304),
        .in(10'h336)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2645 (
        .y(_T_1940),
        .a(io_decode_csr),
        .b(_WTEMP_304)
    );
    wire _T_1942;
    EQ_UNSIGNED #(.width(12)) u_eq_2646 (
        .y(_T_1942),
        .a(io_decode_csr),
        .b(12'hB16)
    );
    wire _T_1944;
    EQ_UNSIGNED #(.width(12)) u_eq_2647 (
        .y(_T_1944),
        .a(io_decode_csr),
        .b(12'hC16)
    );
    wire _T_1946;
    wire [11:0] _WTEMP_305;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2648 (
        .y(_WTEMP_305),
        .in(10'h337)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2649 (
        .y(_T_1946),
        .a(io_decode_csr),
        .b(_WTEMP_305)
    );
    wire _T_1948;
    EQ_UNSIGNED #(.width(12)) u_eq_2650 (
        .y(_T_1948),
        .a(io_decode_csr),
        .b(12'hB17)
    );
    wire _T_1950;
    EQ_UNSIGNED #(.width(12)) u_eq_2651 (
        .y(_T_1950),
        .a(io_decode_csr),
        .b(12'hC17)
    );
    wire _T_1952;
    wire [11:0] _WTEMP_306;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2652 (
        .y(_WTEMP_306),
        .in(10'h338)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2653 (
        .y(_T_1952),
        .a(io_decode_csr),
        .b(_WTEMP_306)
    );
    wire _T_1954;
    EQ_UNSIGNED #(.width(12)) u_eq_2654 (
        .y(_T_1954),
        .a(io_decode_csr),
        .b(12'hB18)
    );
    wire _T_1956;
    EQ_UNSIGNED #(.width(12)) u_eq_2655 (
        .y(_T_1956),
        .a(io_decode_csr),
        .b(12'hC18)
    );
    wire _T_1958;
    wire [11:0] _WTEMP_307;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2656 (
        .y(_WTEMP_307),
        .in(10'h339)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2657 (
        .y(_T_1958),
        .a(io_decode_csr),
        .b(_WTEMP_307)
    );
    wire _T_1960;
    EQ_UNSIGNED #(.width(12)) u_eq_2658 (
        .y(_T_1960),
        .a(io_decode_csr),
        .b(12'hB19)
    );
    wire _T_1962;
    EQ_UNSIGNED #(.width(12)) u_eq_2659 (
        .y(_T_1962),
        .a(io_decode_csr),
        .b(12'hC19)
    );
    wire _T_1964;
    wire [11:0] _WTEMP_308;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2660 (
        .y(_WTEMP_308),
        .in(10'h33A)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2661 (
        .y(_T_1964),
        .a(io_decode_csr),
        .b(_WTEMP_308)
    );
    wire _T_1966;
    EQ_UNSIGNED #(.width(12)) u_eq_2662 (
        .y(_T_1966),
        .a(io_decode_csr),
        .b(12'hB1A)
    );
    wire _T_1968;
    EQ_UNSIGNED #(.width(12)) u_eq_2663 (
        .y(_T_1968),
        .a(io_decode_csr),
        .b(12'hC1A)
    );
    wire _T_1970;
    wire [11:0] _WTEMP_309;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2664 (
        .y(_WTEMP_309),
        .in(10'h33B)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2665 (
        .y(_T_1970),
        .a(io_decode_csr),
        .b(_WTEMP_309)
    );
    wire _T_1972;
    EQ_UNSIGNED #(.width(12)) u_eq_2666 (
        .y(_T_1972),
        .a(io_decode_csr),
        .b(12'hB1B)
    );
    wire _T_1974;
    EQ_UNSIGNED #(.width(12)) u_eq_2667 (
        .y(_T_1974),
        .a(io_decode_csr),
        .b(12'hC1B)
    );
    wire _T_1976;
    wire [11:0] _WTEMP_310;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2668 (
        .y(_WTEMP_310),
        .in(10'h33C)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2669 (
        .y(_T_1976),
        .a(io_decode_csr),
        .b(_WTEMP_310)
    );
    wire _T_1978;
    EQ_UNSIGNED #(.width(12)) u_eq_2670 (
        .y(_T_1978),
        .a(io_decode_csr),
        .b(12'hB1C)
    );
    wire _T_1980;
    EQ_UNSIGNED #(.width(12)) u_eq_2671 (
        .y(_T_1980),
        .a(io_decode_csr),
        .b(12'hC1C)
    );
    wire _T_1982;
    wire [11:0] _WTEMP_311;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2672 (
        .y(_WTEMP_311),
        .in(10'h33D)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2673 (
        .y(_T_1982),
        .a(io_decode_csr),
        .b(_WTEMP_311)
    );
    wire _T_1984;
    EQ_UNSIGNED #(.width(12)) u_eq_2674 (
        .y(_T_1984),
        .a(io_decode_csr),
        .b(12'hB1D)
    );
    wire _T_1986;
    EQ_UNSIGNED #(.width(12)) u_eq_2675 (
        .y(_T_1986),
        .a(io_decode_csr),
        .b(12'hC1D)
    );
    wire _T_1988;
    wire [11:0] _WTEMP_312;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2676 (
        .y(_WTEMP_312),
        .in(10'h33E)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2677 (
        .y(_T_1988),
        .a(io_decode_csr),
        .b(_WTEMP_312)
    );
    wire _T_1990;
    EQ_UNSIGNED #(.width(12)) u_eq_2678 (
        .y(_T_1990),
        .a(io_decode_csr),
        .b(12'hB1E)
    );
    wire _T_1992;
    EQ_UNSIGNED #(.width(12)) u_eq_2679 (
        .y(_T_1992),
        .a(io_decode_csr),
        .b(12'hC1E)
    );
    wire _T_1994;
    wire [11:0] _WTEMP_313;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2680 (
        .y(_WTEMP_313),
        .in(10'h33F)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2681 (
        .y(_T_1994),
        .a(io_decode_csr),
        .b(_WTEMP_313)
    );
    wire _T_1996;
    EQ_UNSIGNED #(.width(12)) u_eq_2682 (
        .y(_T_1996),
        .a(io_decode_csr),
        .b(12'hB1F)
    );
    wire _T_1998;
    EQ_UNSIGNED #(.width(12)) u_eq_2683 (
        .y(_T_1998),
        .a(io_decode_csr),
        .b(12'hC1F)
    );
    wire _T_2000;
    wire [11:0] _WTEMP_314;
    PAD_UNSIGNED #(.width(9), .n(12)) u_pad_2684 (
        .y(_WTEMP_314),
        .in(9'h100)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2685 (
        .y(_T_2000),
        .a(io_decode_csr),
        .b(_WTEMP_314)
    );
    wire _T_2002;
    wire [11:0] _WTEMP_315;
    PAD_UNSIGNED #(.width(9), .n(12)) u_pad_2686 (
        .y(_WTEMP_315),
        .in(9'h144)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2687 (
        .y(_T_2002),
        .a(io_decode_csr),
        .b(_WTEMP_315)
    );
    wire _T_2004;
    wire [11:0] _WTEMP_316;
    PAD_UNSIGNED #(.width(9), .n(12)) u_pad_2688 (
        .y(_WTEMP_316),
        .in(9'h104)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2689 (
        .y(_T_2004),
        .a(io_decode_csr),
        .b(_WTEMP_316)
    );
    wire _T_2006;
    wire [11:0] _WTEMP_317;
    PAD_UNSIGNED #(.width(9), .n(12)) u_pad_2690 (
        .y(_WTEMP_317),
        .in(9'h140)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2691 (
        .y(_T_2006),
        .a(io_decode_csr),
        .b(_WTEMP_317)
    );
    wire _T_2008;
    wire [11:0] _WTEMP_318;
    PAD_UNSIGNED #(.width(9), .n(12)) u_pad_2692 (
        .y(_WTEMP_318),
        .in(9'h142)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2693 (
        .y(_T_2008),
        .a(io_decode_csr),
        .b(_WTEMP_318)
    );
    wire _T_2010;
    wire [11:0] _WTEMP_319;
    PAD_UNSIGNED #(.width(9), .n(12)) u_pad_2694 (
        .y(_WTEMP_319),
        .in(9'h143)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2695 (
        .y(_T_2010),
        .a(io_decode_csr),
        .b(_WTEMP_319)
    );
    wire _T_2012;
    wire [11:0] _WTEMP_320;
    PAD_UNSIGNED #(.width(9), .n(12)) u_pad_2696 (
        .y(_WTEMP_320),
        .in(9'h180)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2697 (
        .y(_T_2012),
        .a(io_decode_csr),
        .b(_WTEMP_320)
    );
    wire _T_2014;
    wire [11:0] _WTEMP_321;
    PAD_UNSIGNED #(.width(9), .n(12)) u_pad_2698 (
        .y(_WTEMP_321),
        .in(9'h141)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2699 (
        .y(_T_2014),
        .a(io_decode_csr),
        .b(_WTEMP_321)
    );
    wire _T_2016;
    wire [11:0] _WTEMP_322;
    PAD_UNSIGNED #(.width(9), .n(12)) u_pad_2700 (
        .y(_WTEMP_322),
        .in(9'h105)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2701 (
        .y(_T_2016),
        .a(io_decode_csr),
        .b(_WTEMP_322)
    );
    wire _T_2018;
    wire [11:0] _WTEMP_323;
    PAD_UNSIGNED #(.width(9), .n(12)) u_pad_2702 (
        .y(_WTEMP_323),
        .in(9'h106)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2703 (
        .y(_T_2018),
        .a(io_decode_csr),
        .b(_WTEMP_323)
    );
    wire _T_2020;
    wire [11:0] _WTEMP_324;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2704 (
        .y(_WTEMP_324),
        .in(10'h306)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2705 (
        .y(_T_2020),
        .a(io_decode_csr),
        .b(_WTEMP_324)
    );
    wire _T_2022;
    EQ_UNSIGNED #(.width(12)) u_eq_2706 (
        .y(_T_2022),
        .a(io_decode_csr),
        .b(12'hC00)
    );
    wire _T_2024;
    EQ_UNSIGNED #(.width(12)) u_eq_2707 (
        .y(_T_2024),
        .a(io_decode_csr),
        .b(12'hC02)
    );
    wire _T_2025;
    BITWISEOR #(.width(1)) bitwiseor_2708 (
        .y(_T_2025),
        .a(_T_1952),
        .b(_T_1820)
    );
    wire _T_2026;
    BITWISEOR #(.width(1)) bitwiseor_2709 (
        .y(_T_2026),
        .a(_T_2025),
        .b(_T_1864)
    );
    wire _T_2027;
    BITWISEOR #(.width(1)) bitwiseor_2710 (
        .y(_T_2027),
        .a(_T_2026),
        .b(_T_2006)
    );
    wire _T_2028;
    BITWISEOR #(.width(1)) bitwiseor_2711 (
        .y(_T_2028),
        .a(_T_2027),
        .b(_T_1978)
    );
    wire _T_2029;
    BITWISEOR #(.width(1)) bitwiseor_2712 (
        .y(_T_2029),
        .a(_T_2028),
        .b(_T_1946)
    );
    wire _T_2030;
    BITWISEOR #(.width(1)) bitwiseor_2713 (
        .y(_T_2030),
        .a(_T_2029),
        .b(_T_1832)
    );
    wire _T_2031;
    BITWISEOR #(.width(1)) bitwiseor_2714 (
        .y(_T_2031),
        .a(_T_2030),
        .b(_T_1800)
    );
    wire _T_2032;
    BITWISEOR #(.width(1)) bitwiseor_2715 (
        .y(_T_2032),
        .a(_T_2031),
        .b(_T_2020)
    );
    wire _T_2033;
    BITWISEOR #(.width(1)) bitwiseor_2716 (
        .y(_T_2033),
        .a(_T_2032),
        .b(_T_1914)
    );
    wire _T_2034;
    BITWISEOR #(.width(1)) bitwiseor_2717 (
        .y(_T_2034),
        .a(_T_2033),
        .b(_T_1876)
    );
    wire _T_2035;
    BITWISEOR #(.width(1)) bitwiseor_2718 (
        .y(_T_2035),
        .a(_T_2034),
        .b(_T_1920)
    );
    wire _T_2036;
    BITWISEOR #(.width(1)) bitwiseor_2719 (
        .y(_T_2036),
        .a(_T_2035),
        .b(_T_1788)
    );
    wire _T_2037;
    BITWISEOR #(.width(1)) bitwiseor_2720 (
        .y(_T_2037),
        .a(_T_2036),
        .b(_T_1844)
    );
    wire _T_2038;
    BITWISEOR #(.width(1)) bitwiseor_2721 (
        .y(_T_2038),
        .a(_T_2037),
        .b(_T_1888)
    );
    wire _T_2039;
    BITWISEOR #(.width(1)) bitwiseor_2722 (
        .y(_T_2039),
        .a(_T_2038),
        .b(_T_1872)
    );
    wire _T_2040;
    BITWISEOR #(.width(1)) bitwiseor_2723 (
        .y(_T_2040),
        .a(_T_2039),
        .b(_T_1988)
    );
    wire _T_2041;
    BITWISEOR #(.width(1)) bitwiseor_2724 (
        .y(_T_2041),
        .a(_T_2040),
        .b(_T_1910)
    );
    wire _T_2042;
    BITWISEOR #(.width(1)) bitwiseor_2725 (
        .y(_T_2042),
        .a(_T_2041),
        .b(_T_1924)
    );
    wire _T_2043;
    BITWISEOR #(.width(1)) bitwiseor_2726 (
        .y(_T_2043),
        .a(_T_2042),
        .b(_T_1776)
    );
    wire _T_2044;
    BITWISEOR #(.width(1)) bitwiseor_2727 (
        .y(_T_2044),
        .a(_T_2043),
        .b(_T_1808)
    );
    wire _T_2045;
    BITWISEOR #(.width(1)) bitwiseor_2728 (
        .y(_T_2045),
        .a(_T_2044),
        .b(_T_1892)
    );
    wire _T_2046;
    BITWISEOR #(.width(1)) bitwiseor_2729 (
        .y(_T_2046),
        .a(_T_2045),
        .b(_T_1840)
    );
    wire _T_2047;
    BITWISEOR #(.width(1)) bitwiseor_2730 (
        .y(_T_2047),
        .a(_T_2046),
        .b(_T_1956)
    );
    wire _T_2048;
    BITWISEOR #(.width(1)) bitwiseor_2731 (
        .y(_T_2048),
        .a(_T_2047),
        .b(_T_2010)
    );
    wire _T_2049;
    BITWISEOR #(.width(1)) bitwiseor_2732 (
        .y(_T_2049),
        .a(_T_2048),
        .b(_T_1868)
    );
    wire _T_2050;
    BITWISEOR #(.width(1)) bitwiseor_2733 (
        .y(_T_2050),
        .a(_T_2049),
        .b(_T_2000)
    );
    wire _T_2051;
    BITWISEOR #(.width(1)) bitwiseor_2734 (
        .y(_T_2051),
        .a(_T_2050),
        .b(_T_1878)
    );
    wire _T_2052;
    BITWISEOR #(.width(1)) bitwiseor_2735 (
        .y(_T_2052),
        .a(_T_2051),
        .b(_T_1942)
    );
    wire _T_2053;
    BITWISEOR #(.width(1)) bitwiseor_2736 (
        .y(_T_2053),
        .a(_T_2052),
        .b(_T_1812)
    );
    wire _T_2054;
    BITWISEOR #(.width(1)) bitwiseor_2737 (
        .y(_T_2054),
        .a(_T_2053),
        .b(_T_1974)
    );
    wire _T_2055;
    BITWISEOR #(.width(1)) bitwiseor_2738 (
        .y(_T_2055),
        .a(_T_2054),
        .b(_T_1968)
    );
    wire _T_2056;
    BITWISEOR #(.width(1)) bitwiseor_2739 (
        .y(_T_2056),
        .a(_T_2055),
        .b(_T_1780)
    );
    wire _T_2057;
    BITWISEOR #(.width(1)) bitwiseor_2740 (
        .y(_T_2057),
        .a(_T_2056),
        .b(_T_1836)
    );
    wire _T_2058;
    BITWISEOR #(.width(1)) bitwiseor_2741 (
        .y(_T_2058),
        .a(_T_2057),
        .b(_T_1996)
    );
    wire _T_2059;
    BITWISEOR #(.width(1)) bitwiseor_2742 (
        .y(_T_2059),
        .a(_T_2058),
        .b(_T_1814)
    );
    wire _T_2060;
    BITWISEOR #(.width(1)) bitwiseor_2743 (
        .y(_T_2060),
        .a(_T_2059),
        .b(_T_1900)
    );
    wire _T_2061;
    BITWISEOR #(.width(1)) bitwiseor_2744 (
        .y(_T_2061),
        .a(_T_2060),
        .b(_T_1846)
    );
    wire _T_2062;
    BITWISEOR #(.width(1)) bitwiseor_2745 (
        .y(_T_2062),
        .a(_T_2061),
        .b(_T_1932)
    );
    wire _T_2063;
    BITWISEOR #(.width(1)) bitwiseor_2746 (
        .y(_T_2063),
        .a(_T_2062),
        .b(_T_1964)
    );
    wire _T_2064;
    BITWISEOR #(.width(1)) bitwiseor_2747 (
        .y(_T_2064),
        .a(_T_2063),
        .b(_T_1782)
    );
    wire _T_2065;
    BITWISEOR #(.width(1)) bitwiseor_2748 (
        .y(_T_2065),
        .a(_T_2064),
        .b(_T_1904)
    );
    wire _T_2066;
    BITWISEOR #(.width(1)) bitwiseor_2749 (
        .y(_T_2066),
        .a(_T_2065),
        .b(_T_1992)
    );
    wire _T_2067;
    BITWISEOR #(.width(1)) bitwiseor_2750 (
        .y(_T_2067),
        .a(_T_2066),
        .b(_T_1860)
    );
    wire _T_2068;
    BITWISEOR #(.width(1)) bitwiseor_2751 (
        .y(_T_2068),
        .a(_T_2067),
        .b(_T_1804)
    );
    wire _T_2069;
    BITWISEOR #(.width(1)) bitwiseor_2752 (
        .y(_T_2069),
        .a(_T_2068),
        .b(_T_1936)
    );
    wire _T_2070;
    BITWISEOR #(.width(1)) bitwiseor_2753 (
        .y(_T_2070),
        .a(_T_2069),
        .b(_T_1960)
    );
    wire _T_2071;
    BITWISEOR #(.width(1)) bitwiseor_2754 (
        .y(_T_2071),
        .a(_T_2070),
        .b(_T_1828)
    );
    wire _T_2072;
    BITWISEOR #(.width(1)) bitwiseor_2755 (
        .y(_T_2072),
        .a(_T_2071),
        .b(_T_1908)
    );
    wire _T_2073;
    BITWISEOR #(.width(1)) bitwiseor_2756 (
        .y(_T_2073),
        .a(_T_2072),
        .b(_T_2024)
    );
    wire _T_2074;
    BITWISEOR #(.width(1)) bitwiseor_2757 (
        .y(_T_2074),
        .a(_T_2073),
        .b(_T_2004)
    );
    wire _T_2075;
    BITWISEOR #(.width(1)) bitwiseor_2758 (
        .y(_T_2075),
        .a(_T_2074),
        .b(_T_1856)
    );
    wire _T_2076;
    BITWISEOR #(.width(1)) bitwiseor_2759 (
        .y(_T_2076),
        .a(_T_2075),
        .b(_T_1940)
    );
    wire _T_2077;
    BITWISEOR #(.width(1)) bitwiseor_2760 (
        .y(_T_2077),
        .a(_T_2076),
        .b(_T_1792)
    );
    wire _T_2078;
    BITWISEOR #(.width(1)) bitwiseor_2761 (
        .y(_T_2078),
        .a(_T_2077),
        .b(_T_1972)
    );
    wire _T_2079;
    BITWISEOR #(.width(1)) bitwiseor_2762 (
        .y(_T_2079),
        .a(_T_2078),
        .b(_T_1824)
    );
    wire _T_2080;
    BITWISEOR #(.width(1)) bitwiseor_2763 (
        .y(_T_2080),
        .a(_T_2079),
        .b(_T_1896)
    );
    wire _T_2081;
    BITWISEOR #(.width(1)) bitwiseor_2764 (
        .y(_T_2081),
        .a(_T_2080),
        .b(_T_1928)
    );
    wire _T_2082;
    BITWISEOR #(.width(1)) bitwiseor_2765 (
        .y(_T_2082),
        .a(_T_2081),
        .b(_T_1796)
    );
    wire _T_2083;
    BITWISEOR #(.width(1)) bitwiseor_2766 (
        .y(_T_2083),
        .a(_T_2082),
        .b(_T_1918)
    );
    wire _T_2084;
    BITWISEOR #(.width(1)) bitwiseor_2767 (
        .y(_T_2084),
        .a(_T_2083),
        .b(_T_1786)
    );
    wire _T_2085;
    BITWISEOR #(.width(1)) bitwiseor_2768 (
        .y(_T_2085),
        .a(_T_2084),
        .b(_T_1980)
    );
    wire _T_2086;
    BITWISEOR #(.width(1)) bitwiseor_2769 (
        .y(_T_2086),
        .a(_T_2085),
        .b(_T_1774)
    );
    wire _T_2087;
    BITWISEOR #(.width(1)) bitwiseor_2770 (
        .y(_T_2087),
        .a(_T_2086),
        .b(_T_1830)
    );
    wire _T_2088;
    BITWISEOR #(.width(1)) bitwiseor_2771 (
        .y(_T_2088),
        .a(_T_2087),
        .b(_T_1890)
    );
    wire _T_2089;
    BITWISEOR #(.width(1)) bitwiseor_2772 (
        .y(_T_2089),
        .a(_T_2088),
        .b(_T_2018)
    );
    wire _T_2090;
    BITWISEOR #(.width(1)) bitwiseor_2773 (
        .y(_T_2090),
        .a(_T_2089),
        .b(_T_1916)
    );
    wire _T_2091;
    BITWISEOR #(.width(1)) bitwiseor_2774 (
        .y(_T_2091),
        .a(_T_2090),
        .b(_T_1884)
    );
    wire _T_2092;
    BITWISEOR #(.width(1)) bitwiseor_2775 (
        .y(_T_2092),
        .a(_T_2091),
        .b(_T_1862)
    );
    wire _T_2093;
    BITWISEOR #(.width(1)) bitwiseor_2776 (
        .y(_T_2093),
        .a(_T_2092),
        .b(_T_1948)
    );
    wire _T_2094;
    BITWISEOR #(.width(1)) bitwiseor_2777 (
        .y(_T_2094),
        .a(_T_2093),
        .b(_T_1798)
    );
    wire _T_2095;
    BITWISEOR #(.width(1)) bitwiseor_2778 (
        .y(_T_2095),
        .a(_T_2094),
        .b(_T_1976)
    );
    wire _T_2096;
    BITWISEOR #(.width(1)) bitwiseor_2779 (
        .y(_T_2096),
        .a(_T_2095),
        .b(_T_1886)
    );
    wire _T_2097;
    BITWISEOR #(.width(1)) bitwiseor_2780 (
        .y(_T_2097),
        .a(_T_2096),
        .b(_T_1950)
    );
    wire _T_2098;
    BITWISEOR #(.width(1)) bitwiseor_2781 (
        .y(_T_2098),
        .a(_T_2097),
        .b(_T_1818)
    );
    wire _T_2099;
    BITWISEOR #(.width(1)) bitwiseor_2782 (
        .y(_T_2099),
        .a(_T_2098),
        .b(_T_1982)
    );
    wire _T_2100;
    BITWISEOR #(.width(1)) bitwiseor_2783 (
        .y(_T_2100),
        .a(_T_2099),
        .b(_T_1850)
    );
    wire _T_2101;
    BITWISEOR #(.width(1)) bitwiseor_2784 (
        .y(_T_2101),
        .a(_T_2100),
        .b(_T_1810)
    );
    wire _T_2102;
    BITWISEOR #(.width(1)) bitwiseor_2785 (
        .y(_T_2102),
        .a(_T_2101),
        .b(_T_1944)
    );
    wire _T_2103;
    BITWISEOR #(.width(1)) bitwiseor_2786 (
        .y(_T_2103),
        .a(_T_2102),
        .b(_T_2014)
    );
    wire _T_2104;
    BITWISEOR #(.width(1)) bitwiseor_2787 (
        .y(_T_2104),
        .a(_T_2103),
        .b(_T_1838)
    );
    wire _T_2105;
    BITWISEOR #(.width(1)) bitwiseor_2788 (
        .y(_T_2105),
        .a(_T_2104),
        .b(_T_1954)
    );
    wire _T_2106;
    BITWISEOR #(.width(1)) bitwiseor_2789 (
        .y(_T_2106),
        .a(_T_2105),
        .b(_T_1870)
    );
    wire _T_2107;
    BITWISEOR #(.width(1)) bitwiseor_2790 (
        .y(_T_2107),
        .a(_T_2106),
        .b(_T_1986)
    );
    wire _T_2108;
    BITWISEOR #(.width(1)) bitwiseor_2791 (
        .y(_T_2108),
        .a(_T_2107),
        .b(_T_2008)
    );
    wire _T_2109;
    BITWISEOR #(.width(1)) bitwiseor_2792 (
        .y(_T_2109),
        .a(_T_2108),
        .b(_T_1922)
    );
    wire _T_2110;
    BITWISEOR #(.width(1)) bitwiseor_2793 (
        .y(_T_2110),
        .a(_T_2109),
        .b(_T_1778)
    );
    wire _T_2111;
    BITWISEOR #(.width(1)) bitwiseor_2794 (
        .y(_T_2111),
        .a(_T_2110),
        .b(_T_1806)
    );
    wire _T_2112;
    BITWISEOR #(.width(1)) bitwiseor_2795 (
        .y(_T_2112),
        .a(_T_2111),
        .b(_T_1842)
    );
    wire _T_2113;
    BITWISEOR #(.width(1)) bitwiseor_2796 (
        .y(_T_2113),
        .a(_T_2112),
        .b(_T_1874)
    );
    wire _T_2114;
    BITWISEOR #(.width(1)) bitwiseor_2797 (
        .y(_T_2114),
        .a(_T_2113),
        .b(_T_1880)
    );
    wire _T_2115;
    BITWISEOR #(.width(1)) bitwiseor_2798 (
        .y(_T_2115),
        .a(_T_2114),
        .b(_T_2012)
    );
    wire _T_2116;
    BITWISEOR #(.width(1)) bitwiseor_2799 (
        .y(_T_2116),
        .a(_T_2115),
        .b(_T_1912)
    );
    wire _T_2117;
    BITWISEOR #(.width(1)) bitwiseor_2800 (
        .y(_T_2117),
        .a(_T_2116),
        .b(_T_1802)
    );
    wire _T_2118;
    BITWISEOR #(.width(1)) bitwiseor_2801 (
        .y(_T_2118),
        .a(_T_2117),
        .b(_T_1934)
    );
    wire _T_2119;
    BITWISEOR #(.width(1)) bitwiseor_2802 (
        .y(_T_2119),
        .a(_T_2118),
        .b(_T_1848)
    );
    wire _T_2120;
    BITWISEOR #(.width(1)) bitwiseor_2803 (
        .y(_T_2120),
        .a(_T_2119),
        .b(_T_1962)
    );
    wire _T_2121;
    BITWISEOR #(.width(1)) bitwiseor_2804 (
        .y(_T_2121),
        .a(_T_2120),
        .b(_T_1784)
    );
    wire _T_2122;
    BITWISEOR #(.width(1)) bitwiseor_2805 (
        .y(_T_2122),
        .a(_T_2121),
        .b(_T_1902)
    );
    wire _T_2123;
    BITWISEOR #(.width(1)) bitwiseor_2806 (
        .y(_T_2123),
        .a(_T_2122),
        .b(_T_1994)
    );
    wire _T_2124;
    BITWISEOR #(.width(1)) bitwiseor_2807 (
        .y(_T_2124),
        .a(_T_2123),
        .b(_T_2016)
    );
    wire _T_2125;
    BITWISEOR #(.width(1)) bitwiseor_2808 (
        .y(_T_2125),
        .a(_T_2124),
        .b(_T_1930)
    );
    wire _T_2126;
    BITWISEOR #(.width(1)) bitwiseor_2809 (
        .y(_T_2126),
        .a(_T_2125),
        .b(_T_1816)
    );
    wire _T_2127;
    BITWISEOR #(.width(1)) bitwiseor_2810 (
        .y(_T_2127),
        .a(_T_2126),
        .b(_T_1834)
    );
    wire _T_2128;
    BITWISEOR #(.width(1)) bitwiseor_2811 (
        .y(_T_2128),
        .a(_T_2127),
        .b(_T_1966)
    );
    wire _T_2129;
    BITWISEOR #(.width(1)) bitwiseor_2812 (
        .y(_T_2129),
        .a(_T_2128),
        .b(_T_1898)
    );
    wire _T_2130;
    BITWISEOR #(.width(1)) bitwiseor_2813 (
        .y(_T_2130),
        .a(_T_2129),
        .b(_T_1866)
    );
    wire _T_2131;
    BITWISEOR #(.width(1)) bitwiseor_2814 (
        .y(_T_2131),
        .a(_T_2130),
        .b(_T_1998)
    );
    wire _T_2132;
    BITWISEOR #(.width(1)) bitwiseor_2815 (
        .y(_T_2132),
        .a(_T_2131),
        .b(_T_1926)
    );
    wire _T_2133;
    BITWISEOR #(.width(1)) bitwiseor_2816 (
        .y(_T_2133),
        .a(_T_2132),
        .b(_T_1794)
    );
    wire _T_2134;
    BITWISEOR #(.width(1)) bitwiseor_2817 (
        .y(_T_2134),
        .a(_T_2133),
        .b(_T_1882)
    );
    wire _T_2135;
    BITWISEOR #(.width(1)) bitwiseor_2818 (
        .y(_T_2135),
        .a(_T_2134),
        .b(_T_1970)
    );
    wire _T_2136;
    BITWISEOR #(.width(1)) bitwiseor_2819 (
        .y(_T_2136),
        .a(_T_2135),
        .b(_T_1822)
    );
    wire _T_2137;
    BITWISEOR #(.width(1)) bitwiseor_2820 (
        .y(_T_2137),
        .a(_T_2136),
        .b(_T_1894)
    );
    wire _T_2138;
    BITWISEOR #(.width(1)) bitwiseor_2821 (
        .y(_T_2138),
        .a(_T_2137),
        .b(_T_2002)
    );
    wire _T_2139;
    BITWISEOR #(.width(1)) bitwiseor_2822 (
        .y(_T_2139),
        .a(_T_2138),
        .b(_T_1854)
    );
    wire _T_2140;
    BITWISEOR #(.width(1)) bitwiseor_2823 (
        .y(_T_2140),
        .a(_T_2139),
        .b(_T_1938)
    );
    wire _T_2141;
    BITWISEOR #(.width(1)) bitwiseor_2824 (
        .y(_T_2141),
        .a(_T_2140),
        .b(_T_1984)
    );
    wire _T_2142;
    BITWISEOR #(.width(1)) bitwiseor_2825 (
        .y(_T_2142),
        .a(_T_2141),
        .b(_T_1790)
    );
    wire _T_2143;
    BITWISEOR #(.width(1)) bitwiseor_2826 (
        .y(_T_2143),
        .a(_T_2142),
        .b(_T_1852)
    );
    wire _T_2144;
    BITWISEOR #(.width(1)) bitwiseor_2827 (
        .y(_T_2144),
        .a(_T_2143),
        .b(_T_1958)
    );
    wire _T_2145;
    BITWISEOR #(.width(1)) bitwiseor_2828 (
        .y(_T_2145),
        .a(_T_2144),
        .b(_T_1826)
    );
    wire _T_2146;
    BITWISEOR #(.width(1)) bitwiseor_2829 (
        .y(_T_2146),
        .a(_T_2145),
        .b(_T_2022)
    );
    wire _T_2147;
    BITWISEOR #(.width(1)) bitwiseor_2830 (
        .y(_T_2147),
        .a(_T_2146),
        .b(_T_1906)
    );
    wire _T_2148;
    BITWISEOR #(.width(1)) bitwiseor_2831 (
        .y(_T_2148),
        .a(_T_2147),
        .b(_T_1990)
    );
    wire _T_2149;
    BITWISEOR #(.width(1)) bitwiseor_2832 (
        .y(_T_2149),
        .a(_T_2148),
        .b(_T_1858)
    );
    wire _T_2151;
    EQ_UNSIGNED #(.width(1)) u_eq_2833 (
        .y(_T_2151),
        .a(_T_2149),
        .b(1'h0)
    );
    wire _T_2152;
    BITWISEOR #(.width(1)) bitwiseor_2834 (
        .y(_T_2152),
        .a(_T_1772),
        .b(_T_2151)
    );
    wire _T_2154;
    wire [11:0] _WTEMP_325;
    PAD_UNSIGNED #(.width(9), .n(12)) u_pad_2835 (
        .y(_WTEMP_325),
        .in(9'h180)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2836 (
        .y(_T_2154),
        .a(io_decode_csr),
        .b(_WTEMP_325)
    );
    wire _T_2156;
    EQ_UNSIGNED #(.width(1)) u_eq_2837 (
        .y(_T_2156),
        .a(allow_sfence_vma),
        .b(1'h0)
    );
    wire _T_2157;
    BITWISEAND #(.width(1)) bitwiseand_2838 (
        .y(_T_2157),
        .a(_T_2154),
        .b(_T_2156)
    );
    wire _T_2158;
    BITWISEOR #(.width(1)) bitwiseor_2839 (
        .y(_T_2158),
        .a(_T_2152),
        .b(_T_2157)
    );
    wire _T_2161;
    GEQ_UNSIGNED #(.width(12)) u_geq_2840 (
        .y(_T_2161),
        .a(io_decode_csr),
        .b(12'hC00)
    );
    wire _T_2162;
    LT_UNSIGNED #(.width(12)) u_lt_2841 (
        .y(_T_2162),
        .a(io_decode_csr),
        .b(12'hC20)
    );
    wire _T_2163;
    BITWISEAND #(.width(1)) bitwiseand_2842 (
        .y(_T_2163),
        .a(_T_2161),
        .b(_T_2162)
    );
    wire _T_2166;
    GEQ_UNSIGNED #(.width(12)) u_geq_2843 (
        .y(_T_2166),
        .a(io_decode_csr),
        .b(12'hC80)
    );
    wire _T_2167;
    LT_UNSIGNED #(.width(12)) u_lt_2844 (
        .y(_T_2167),
        .a(io_decode_csr),
        .b(12'hCA0)
    );
    wire _T_2168;
    BITWISEAND #(.width(1)) bitwiseand_2845 (
        .y(_T_2168),
        .a(_T_2166),
        .b(_T_2167)
    );
    wire _T_2169;
    BITWISEOR #(.width(1)) bitwiseor_2846 (
        .y(_T_2169),
        .a(_T_2163),
        .b(_T_2168)
    );
    wire _T_2171;
    wire [2:0] _WTEMP_326;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_2847 (
        .y(_WTEMP_326),
        .in(1'h1)
    );
    LEQ_UNSIGNED #(.width(3)) u_leq_2848 (
        .y(_T_2171),
        .a(effective_prv),
        .b(_WTEMP_326)
    );
    wire _T_2172;
    BITWISEAND #(.width(1)) bitwiseand_2849 (
        .y(_T_2172),
        .a(_T_2169),
        .b(_T_2171)
    );
    wire [11:0] _T_2173;
    BITS #(.width(12), .high(11), .low(0)) bits_2850 (
        .y(_T_2173),
        .in(io_decode_csr)
    );
    wire [31:0] _T_2174;
    DSHR_UNSIGNED #(.width_in(32), .width_n(12)) u_dshr_2851 (
        .y(_T_2174),
        .in(hpm_mask),
        .n(_T_2173)
    );
    wire _T_2175;
    BITS #(.width(32), .high(0), .low(0)) bits_2852 (
        .y(_T_2175),
        .in(_T_2174)
    );
    wire _T_2176;
    BITWISEAND #(.width(1)) bitwiseand_2853 (
        .y(_T_2176),
        .a(_T_2172),
        .b(_T_2175)
    );
    wire _T_2177;
    BITWISEOR #(.width(1)) bitwiseor_2854 (
        .y(_T_2177),
        .a(_T_2158),
        .b(_T_2176)
    );
    wire _T_2180;
    EQ_UNSIGNED #(.width(1)) u_eq_2855 (
        .y(_T_2180),
        .a(_reg_debug__q),
        .b(1'h0)
    );
    wire _T_2181;
    BITWISEAND #(.width(1)) bitwiseand_2856 (
        .y(_T_2181),
        .a(1'h1),
        .b(_T_2180)
    );
    wire _T_2183;
    wire [11:0] _WTEMP_327;
    PAD_UNSIGNED #(.width(11), .n(12)) u_pad_2857 (
        .y(_WTEMP_327),
        .in(11'h7B0)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2858 (
        .y(_T_2183),
        .a(io_decode_csr),
        .b(_WTEMP_327)
    );
    wire _T_2185;
    wire [11:0] _WTEMP_328;
    PAD_UNSIGNED #(.width(11), .n(12)) u_pad_2859 (
        .y(_WTEMP_328),
        .in(11'h7B1)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2860 (
        .y(_T_2185),
        .a(io_decode_csr),
        .b(_WTEMP_328)
    );
    wire _T_2187;
    wire [11:0] _WTEMP_329;
    PAD_UNSIGNED #(.width(11), .n(12)) u_pad_2861 (
        .y(_WTEMP_329),
        .in(11'h7B2)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2862 (
        .y(_T_2187),
        .a(io_decode_csr),
        .b(_WTEMP_329)
    );
    wire _T_2188;
    BITWISEOR #(.width(1)) bitwiseor_2863 (
        .y(_T_2188),
        .a(_T_2183),
        .b(_T_2185)
    );
    wire _T_2189;
    BITWISEOR #(.width(1)) bitwiseor_2864 (
        .y(_T_2189),
        .a(_T_2188),
        .b(_T_2187)
    );
    wire _T_2190;
    BITWISEAND #(.width(1)) bitwiseand_2865 (
        .y(_T_2190),
        .a(_T_2181),
        .b(_T_2189)
    );
    wire _T_2191;
    BITWISEOR #(.width(1)) bitwiseor_2866 (
        .y(_T_2191),
        .a(_T_2177),
        .b(_T_2190)
    );
    wire _T_2194;
    wire [11:0] _WTEMP_330;
    PAD_UNSIGNED #(.width(1), .n(12)) u_pad_2867 (
        .y(_WTEMP_330),
        .in(1'h1)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2868 (
        .y(_T_2194),
        .a(io_decode_csr),
        .b(_WTEMP_330)
    );
    wire _T_2196;
    wire [11:0] _WTEMP_331;
    PAD_UNSIGNED #(.width(2), .n(12)) u_pad_2869 (
        .y(_WTEMP_331),
        .in(2'h2)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2870 (
        .y(_T_2196),
        .a(io_decode_csr),
        .b(_WTEMP_331)
    );
    wire _T_2198;
    wire [11:0] _WTEMP_332;
    PAD_UNSIGNED #(.width(2), .n(12)) u_pad_2871 (
        .y(_WTEMP_332),
        .in(2'h3)
    );
    EQ_UNSIGNED #(.width(12)) u_eq_2872 (
        .y(_T_2198),
        .a(io_decode_csr),
        .b(_WTEMP_332)
    );
    wire _T_2199;
    BITWISEOR #(.width(1)) bitwiseor_2873 (
        .y(_T_2199),
        .a(_T_2194),
        .b(_T_2196)
    );
    wire _T_2200;
    BITWISEOR #(.width(1)) bitwiseor_2874 (
        .y(_T_2200),
        .a(_T_2199),
        .b(_T_2198)
    );
    wire _T_2201;
    BITWISEAND #(.width(1)) bitwiseand_2875 (
        .y(_T_2201),
        .a(1'h1),
        .b(_T_2200)
    );
    wire _T_2202;
    BITWISEAND #(.width(1)) bitwiseand_2876 (
        .y(_T_2202),
        .a(_T_2201),
        .b(io_decode_fp_illegal)
    );
    wire _T_2203;
    BITWISEOR #(.width(1)) bitwiseor_2877 (
        .y(_T_2203),
        .a(_T_2191),
        .b(_T_2202)
    );
    wire [1:0] _T_2204;
    BITS #(.width(12), .high(11), .low(10)) bits_2878 (
        .y(_T_2204),
        .in(io_decode_csr)
    );
    wire [1:0] _T_2205;
    BITWISENOT #(.width(2)) bitwisenot_2879 (
        .y(_T_2205),
        .in(_T_2204)
    );
    wire _T_2207;
    wire [1:0] _WTEMP_333;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2880 (
        .y(_WTEMP_333),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(2)) u_eq_2881 (
        .y(_T_2207),
        .a(_T_2205),
        .b(_WTEMP_333)
    );
    wire _T_2209;
    wire [11:0] _WTEMP_334;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2882 (
        .y(_WTEMP_334),
        .in(10'h340)
    );
    GEQ_UNSIGNED #(.width(12)) u_geq_2883 (
        .y(_T_2209),
        .a(io_decode_csr),
        .b(_WTEMP_334)
    );
    wire _T_2211;
    wire [11:0] _WTEMP_335;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2884 (
        .y(_WTEMP_335),
        .in(10'h343)
    );
    LEQ_UNSIGNED #(.width(12)) u_leq_2885 (
        .y(_T_2211),
        .a(io_decode_csr),
        .b(_WTEMP_335)
    );
    wire _T_2212;
    BITWISEAND #(.width(1)) bitwiseand_2886 (
        .y(_T_2212),
        .a(_T_2209),
        .b(_T_2211)
    );
    wire _T_2214;
    wire [11:0] _WTEMP_336;
    PAD_UNSIGNED #(.width(9), .n(12)) u_pad_2887 (
        .y(_WTEMP_336),
        .in(9'h140)
    );
    GEQ_UNSIGNED #(.width(12)) u_geq_2888 (
        .y(_T_2214),
        .a(io_decode_csr),
        .b(_WTEMP_336)
    );
    wire _T_2216;
    wire [11:0] _WTEMP_337;
    PAD_UNSIGNED #(.width(9), .n(12)) u_pad_2889 (
        .y(_WTEMP_337),
        .in(9'h143)
    );
    LEQ_UNSIGNED #(.width(12)) u_leq_2890 (
        .y(_T_2216),
        .a(io_decode_csr),
        .b(_WTEMP_337)
    );
    wire _T_2217;
    BITWISEAND #(.width(1)) bitwiseand_2891 (
        .y(_T_2217),
        .a(_T_2214),
        .b(_T_2216)
    );
    wire _T_2218;
    BITWISEOR #(.width(1)) bitwiseor_2892 (
        .y(_T_2218),
        .a(_T_2212),
        .b(_T_2217)
    );
    wire _T_2220;
    EQ_UNSIGNED #(.width(1)) u_eq_2893 (
        .y(_T_2220),
        .a(_T_2218),
        .b(1'h0)
    );
    wire [1:0] _T_2221;
    BITS #(.width(12), .high(9), .low(8)) bits_2894 (
        .y(_T_2221),
        .in(io_decode_csr)
    );
    wire _T_2222;
    wire [2:0] _WTEMP_338;
    PAD_UNSIGNED #(.width(2), .n(3)) u_pad_2895 (
        .y(_WTEMP_338),
        .in(_T_2221)
    );
    LT_UNSIGNED #(.width(3)) u_lt_2896 (
        .y(_T_2222),
        .a(effective_prv),
        .b(_WTEMP_338)
    );
    wire _T_2223;
    BITS #(.width(12), .high(5), .low(5)) bits_2897 (
        .y(_T_2223),
        .in(io_decode_csr)
    );
    wire _T_2225;
    EQ_UNSIGNED #(.width(1)) u_eq_2898 (
        .y(_T_2225),
        .a(_T_2223),
        .b(1'h0)
    );
    wire _T_2226;
    BITS #(.width(12), .high(2), .low(2)) bits_2899 (
        .y(_T_2226),
        .in(io_decode_csr)
    );
    wire _T_2227;
    BITWISEAND #(.width(1)) bitwiseand_2900 (
        .y(_T_2227),
        .a(_T_2225),
        .b(_T_2226)
    );
    wire _T_2229;
    EQ_UNSIGNED #(.width(1)) u_eq_2901 (
        .y(_T_2229),
        .a(allow_wfi),
        .b(1'h0)
    );
    wire _T_2230;
    BITWISEAND #(.width(1)) bitwiseand_2902 (
        .y(_T_2230),
        .a(_T_2227),
        .b(_T_2229)
    );
    wire _T_2231;
    BITWISEOR #(.width(1)) bitwiseor_2903 (
        .y(_T_2231),
        .a(_T_2222),
        .b(_T_2230)
    );
    wire _T_2232;
    BITS #(.width(12), .high(5), .low(5)) bits_2904 (
        .y(_T_2232),
        .in(io_decode_csr)
    );
    wire _T_2234;
    EQ_UNSIGNED #(.width(1)) u_eq_2905 (
        .y(_T_2234),
        .a(_T_2232),
        .b(1'h0)
    );
    wire _T_2235;
    BITS #(.width(12), .high(1), .low(1)) bits_2906 (
        .y(_T_2235),
        .in(io_decode_csr)
    );
    wire _T_2236;
    BITWISEAND #(.width(1)) bitwiseand_2907 (
        .y(_T_2236),
        .a(_T_2234),
        .b(_T_2235)
    );
    wire _T_2238;
    EQ_UNSIGNED #(.width(1)) u_eq_2908 (
        .y(_T_2238),
        .a(allow_sret),
        .b(1'h0)
    );
    wire _T_2239;
    BITWISEAND #(.width(1)) bitwiseand_2909 (
        .y(_T_2239),
        .a(_T_2236),
        .b(_T_2238)
    );
    wire _T_2240;
    BITWISEOR #(.width(1)) bitwiseor_2910 (
        .y(_T_2240),
        .a(_T_2231),
        .b(_T_2239)
    );
    wire _T_2241;
    BITS #(.width(12), .high(5), .low(5)) bits_2911 (
        .y(_T_2241),
        .in(io_decode_csr)
    );
    wire _T_2243;
    EQ_UNSIGNED #(.width(1)) u_eq_2912 (
        .y(_T_2243),
        .a(allow_sfence_vma),
        .b(1'h0)
    );
    wire _T_2244;
    BITWISEAND #(.width(1)) bitwiseand_2913 (
        .y(_T_2244),
        .a(_T_2241),
        .b(_T_2243)
    );
    wire _T_2245;
    BITWISEOR #(.width(1)) bitwiseor_2914 (
        .y(_T_2245),
        .a(_T_2240),
        .b(_T_2244)
    );
    wire [4:0] _T_2247;
    wire [3:0] _WTEMP_339;
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_2915 (
        .y(_WTEMP_339),
        .in(_reg_mstatus_prv__q)
    );
    ADD_UNSIGNED #(.width(4)) u_add_2916 (
        .y(_T_2247),
        .a(_WTEMP_339),
        .b(4'h8)
    );
    wire [3:0] _T_2248;
    TAIL #(.width(5), .n(1)) tail_2917 (
        .y(_T_2248),
        .in(_T_2247)
    );
    wire [63:0] _T_2250;
    wire [63:0] _WTEMP_340;
    PAD_UNSIGNED #(.width(2), .n(64)) u_pad_2918 (
        .y(_WTEMP_340),
        .in(2'h3)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_2919 (
        .y(_T_2250),
        .sel(insn_break),
        .a(_WTEMP_340),
        .b(io_cause)
    );
    wire [63:0] cause;
    wire [63:0] _WTEMP_341;
    PAD_UNSIGNED #(.width(4), .n(64)) u_pad_2920 (
        .y(_WTEMP_341),
        .in(_T_2248)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_2921 (
        .y(cause),
        .sel(insn_call),
        .a(_WTEMP_341),
        .b(_T_2250)
    );
    wire [5:0] cause_lsbs;
    BITS #(.width(64), .high(5), .low(0)) bits_2922 (
        .y(cause_lsbs),
        .in(cause)
    );
    wire _T_2251;
    BITS #(.width(64), .high(63), .low(63)) bits_2923 (
        .y(_T_2251),
        .in(cause)
    );
    wire _T_2267;
    wire [5:0] _WTEMP_342;
    PAD_UNSIGNED #(.width(4), .n(6)) u_pad_2924 (
        .y(_WTEMP_342),
        .in(4'hD)
    );
    EQ_UNSIGNED #(.width(6)) u_eq_2925 (
        .y(_T_2267),
        .a(cause_lsbs),
        .b(_WTEMP_342)
    );
    wire causeIsDebugInt;
    BITWISEAND #(.width(1)) bitwiseand_2926 (
        .y(causeIsDebugInt),
        .a(_T_2251),
        .b(_T_2267)
    );
    wire _T_2268;
    BITS #(.width(64), .high(63), .low(63)) bits_2927 (
        .y(_T_2268),
        .in(cause)
    );
    wire _T_2270;
    EQ_UNSIGNED #(.width(1)) u_eq_2928 (
        .y(_T_2270),
        .a(_T_2268),
        .b(1'h0)
    );
    wire _T_2300;
    wire [5:0] _WTEMP_343;
    PAD_UNSIGNED #(.width(4), .n(6)) u_pad_2929 (
        .y(_WTEMP_343),
        .in(4'hD)
    );
    EQ_UNSIGNED #(.width(6)) u_eq_2930 (
        .y(_T_2300),
        .a(cause_lsbs),
        .b(_WTEMP_343)
    );
    wire causeIsDebugTrigger;
    BITWISEAND #(.width(1)) bitwiseand_2931 (
        .y(causeIsDebugTrigger),
        .a(_T_2270),
        .b(_T_2300)
    );
    wire _T_2301;
    BITS #(.width(64), .high(63), .low(63)) bits_2932 (
        .y(_T_2301),
        .in(cause)
    );
    wire _T_2303;
    EQ_UNSIGNED #(.width(1)) u_eq_2933 (
        .y(_T_2303),
        .a(_T_2301),
        .b(1'h0)
    );
    wire _T_2304;
    BITWISEAND #(.width(1)) bitwiseand_2934 (
        .y(_T_2304),
        .a(_T_2303),
        .b(insn_break)
    );
    wire [1:0] _T_2305;
    CAT #(.width_a(1), .width_b(1)) cat_2935 (
        .y(_T_2305),
        .a(_reg_dcsr_ebreaks__q),
        .b(_reg_dcsr_ebreaku__q)
    );
    wire [1:0] _T_2306;
    CAT #(.width_a(1), .width_b(1)) cat_2936 (
        .y(_T_2306),
        .a(_reg_dcsr_ebreakm__q),
        .b(1'h0)
    );
    wire [3:0] _T_2307;
    CAT #(.width_a(2), .width_b(2)) cat_2937 (
        .y(_T_2307),
        .a(_T_2306),
        .b(_T_2305)
    );
    wire [3:0] _T_2308;
    DSHR_UNSIGNED #(.width_in(4), .width_n(2)) u_dshr_2938 (
        .y(_T_2308),
        .in(_T_2307),
        .n(_reg_mstatus_prv__q)
    );
    wire _T_2309;
    BITS #(.width(4), .high(0), .low(0)) bits_2939 (
        .y(_T_2309),
        .in(_T_2308)
    );
    wire causeIsDebugBreak;
    BITWISEAND #(.width(1)) bitwiseand_2940 (
        .y(causeIsDebugBreak),
        .a(_T_2304),
        .b(_T_2309)
    );
    wire _T_2311;
    BITWISEOR #(.width(1)) bitwiseor_2941 (
        .y(_T_2311),
        .a(_reg_singleStepped__q),
        .b(causeIsDebugInt)
    );
    wire _T_2312;
    BITWISEOR #(.width(1)) bitwiseor_2942 (
        .y(_T_2312),
        .a(_T_2311),
        .b(causeIsDebugTrigger)
    );
    wire _T_2313;
    BITWISEOR #(.width(1)) bitwiseor_2943 (
        .y(_T_2313),
        .a(_T_2312),
        .b(causeIsDebugBreak)
    );
    wire _T_2314;
    BITWISEOR #(.width(1)) bitwiseor_2944 (
        .y(_T_2314),
        .a(_T_2313),
        .b(_reg_debug__q)
    );
    wire trapToDebug;
    BITWISEAND #(.width(1)) bitwiseand_2945 (
        .y(trapToDebug),
        .a(1'h1),
        .b(_T_2314)
    );
    wire _T_2317;
    wire [1:0] _WTEMP_344;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2946 (
        .y(_WTEMP_344),
        .in(1'h1)
    );
    LEQ_UNSIGNED #(.width(2)) u_leq_2947 (
        .y(_T_2317),
        .a(_reg_mstatus_prv__q),
        .b(_WTEMP_344)
    );
    wire _T_2318;
    BITWISEAND #(.width(1)) bitwiseand_2948 (
        .y(_T_2318),
        .a(1'h1),
        .b(_T_2317)
    );
    wire _T_2319;
    BITS #(.width(64), .high(63), .low(63)) bits_2949 (
        .y(_T_2319),
        .in(cause)
    );
    wire [63:0] _T_2320;
    DSHR_UNSIGNED #(.width_in(64), .width_n(6)) u_dshr_2950 (
        .y(_T_2320),
        .in(_reg_mideleg__q),
        .n(cause_lsbs)
    );
    wire _T_2321;
    BITS #(.width(64), .high(0), .low(0)) bits_2951 (
        .y(_T_2321),
        .in(_T_2320)
    );
    wire [63:0] _T_2322;
    DSHR_UNSIGNED #(.width_in(64), .width_n(6)) u_dshr_2952 (
        .y(_T_2322),
        .in(_reg_medeleg__q),
        .n(cause_lsbs)
    );
    wire _T_2323;
    BITS #(.width(64), .high(0), .low(0)) bits_2953 (
        .y(_T_2323),
        .in(_T_2322)
    );
    wire _T_2324;
    MUX_UNSIGNED #(.width(1)) u_mux_2954 (
        .y(_T_2324),
        .sel(_T_2319),
        .a(_T_2321),
        .b(_T_2323)
    );
    wire delegate;
    BITWISEAND #(.width(1)) bitwiseand_2955 (
        .y(delegate),
        .a(_T_2318),
        .b(_T_2324)
    );
    wire [11:0] debugTVec;
    MUX_UNSIGNED #(.width(12)) u_mux_2956 (
        .y(debugTVec),
        .sel(_reg_debug__q),
        .a(12'h808),
        .b(12'h800)
    );
    wire _T_2327;
    BITS #(.width(39), .high(38), .low(38)) bits_2957 (
        .y(_T_2327),
        .in(_reg_stvec__q)
    );
    wire [39:0] _T_2328;
    CAT #(.width_a(1), .width_b(39)) cat_2958 (
        .y(_T_2328),
        .a(_T_2327),
        .b(_reg_stvec__q)
    );
    wire [39:0] _T_2329;
    wire [39:0] _WTEMP_345;
    PAD_UNSIGNED #(.width(32), .n(40)) u_pad_2959 (
        .y(_WTEMP_345),
        .in(_reg_mtvec__q)
    );
    MUX_UNSIGNED #(.width(40)) u_mux_2960 (
        .y(_T_2329),
        .sel(delegate),
        .a(_T_2328),
        .b(_WTEMP_345)
    );
    wire [39:0] tvec;
    wire [39:0] _WTEMP_346;
    PAD_UNSIGNED #(.width(12), .n(40)) u_pad_2961 (
        .y(_WTEMP_346),
        .in(debugTVec)
    );
    MUX_UNSIGNED #(.width(40)) u_mux_2962 (
        .y(tvec),
        .sel(trapToDebug),
        .a(_WTEMP_346),
        .b(_T_2329)
    );
    wire _T_2330;
    BITWISEOR #(.width(1)) bitwiseor_2963 (
        .y(_T_2330),
        .a(insn_call),
        .b(insn_break)
    );
    wire _T_2331;
    BITWISEOR #(.width(1)) bitwiseor_2964 (
        .y(_T_2331),
        .a(_T_2330),
        .b(insn_ret)
    );
    wire _T_2333;
    EQ_UNSIGNED #(.width(1)) u_eq_2965 (
        .y(_T_2333),
        .a(_reg_debug__q),
        .b(1'h0)
    );
    wire _T_2334;
    BITWISEAND #(.width(1)) bitwiseand_2966 (
        .y(_T_2334),
        .a(_reg_dcsr_step__q),
        .b(_T_2333)
    );
    wire [1:0] _T_2335;
    BITWISENOT #(.width(2)) bitwisenot_2967 (
        .y(_T_2335),
        .in(io_status_fs)
    );
    wire _T_2337;
    wire [1:0] _WTEMP_347;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2968 (
        .y(_WTEMP_347),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(2)) u_eq_2969 (
        .y(_T_2337),
        .a(_T_2335),
        .b(_WTEMP_347)
    );
    wire [1:0] _T_2338;
    BITWISENOT #(.width(2)) bitwisenot_2970 (
        .y(_T_2338),
        .in(io_status_xs)
    );
    wire _T_2340;
    wire [1:0] _WTEMP_348;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2971 (
        .y(_WTEMP_348),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(2)) u_eq_2972 (
        .y(_T_2340),
        .a(_T_2338),
        .b(_WTEMP_348)
    );
    wire _T_2341;
    BITWISEOR #(.width(1)) bitwiseor_2973 (
        .y(_T_2341),
        .a(_T_2337),
        .b(_T_2340)
    );
    wire _T_2344;
    BITWISEOR #(.width(1)) bitwiseor_2974 (
        .y(_T_2344),
        .a(insn_call),
        .b(insn_break)
    );
    wire exception;
    BITWISEOR #(.width(1)) bitwiseor_2975 (
        .y(exception),
        .a(_T_2344),
        .b(io_exception)
    );
    wire [1:0] _T_2345;
    ADD_UNSIGNED #(.width(1)) u_add_2976 (
        .y(_T_2345),
        .a(insn_ret),
        .b(insn_call)
    );
    wire [1:0] _T_2346;
    ADD_UNSIGNED #(.width(1)) u_add_2977 (
        .y(_T_2346),
        .a(insn_break),
        .b(io_exception)
    );
    wire [2:0] _T_2347;
    ADD_UNSIGNED #(.width(2)) u_add_2978 (
        .y(_T_2347),
        .a(_T_2345),
        .b(_T_2346)
    );
    wire _T_2349;
    wire [2:0] _WTEMP_349;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_2979 (
        .y(_WTEMP_349),
        .in(1'h1)
    );
    LEQ_UNSIGNED #(.width(3)) u_leq_2980 (
        .y(_T_2349),
        .a(_T_2347),
        .b(_WTEMP_349)
    );
    wire _T_2350;
    BITWISEOR #(.width(1)) bitwiseor_2981 (
        .y(_T_2350),
        .a(_T_2349),
        .b(reset)
    );
    wire _T_2352;
    EQ_UNSIGNED #(.width(1)) u_eq_2982 (
        .y(_T_2352),
        .a(_T_2350),
        .b(1'h0)
    );
    wire _T_2355;
    wire [63:0] _WTEMP_350;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_2983 (
        .y(_WTEMP_350),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(64)) u_neq_2984 (
        .y(_T_2355),
        .a(pending_interrupts),
        .b(_WTEMP_350)
    );
    wire _T_2356;
    BITWISEOR #(.width(1)) bitwiseor_2985 (
        .y(_T_2356),
        .a(_T_2355),
        .b(exception)
    );
    wire _node_8;
    MUX_UNSIGNED #(.width(1)) u_mux_2986 (
        .y(_node_8),
        .sel(insn_wfi),
        .a(1'h1),
        .b(_reg_wfi__q)
    );
    wire _T_2359;
    EQ_UNSIGNED #(.width(1)) u_eq_2987 (
        .y(_T_2359),
        .a(_reg_wfi__q),
        .b(1'h0)
    );
    wire _T_2361;
    EQ_UNSIGNED #(.width(1)) u_eq_2988 (
        .y(_T_2361),
        .a(io_retire),
        .b(1'h0)
    );
    wire _T_2362;
    BITWISEOR #(.width(1)) bitwiseor_2989 (
        .y(_T_2362),
        .a(_T_2359),
        .b(_T_2361)
    );
    wire _T_2363;
    BITWISEOR #(.width(1)) bitwiseor_2990 (
        .y(_T_2363),
        .a(_T_2362),
        .b(reset)
    );
    wire _T_2365;
    EQ_UNSIGNED #(.width(1)) u_eq_2991 (
        .y(_T_2365),
        .a(_T_2363),
        .b(1'h0)
    );
    wire _T_2366;
    BITS #(.width(1), .high(0), .low(0)) bits_2992 (
        .y(_T_2366),
        .in(io_retire)
    );
    wire _T_2369;
    EQ_UNSIGNED #(.width(1)) u_eq_2993 (
        .y(_T_2369),
        .a(io_singleStep),
        .b(1'h0)
    );
    wire _node_9;
    MUX_UNSIGNED #(.width(1)) u_mux_2994 (
        .y(_node_9),
        .sel(_T_2366),
        .a(1'h1),
        .b(_reg_singleStepped__q)
    );
    wire _T_2372;
    EQ_UNSIGNED #(.width(1)) u_eq_2995 (
        .y(_T_2372),
        .a(io_singleStep),
        .b(1'h0)
    );
    wire _T_2374;
    LEQ_UNSIGNED #(.width(1)) u_leq_2996 (
        .y(_T_2374),
        .a(io_retire),
        .b(1'h1)
    );
    wire _T_2375;
    BITWISEOR #(.width(1)) bitwiseor_2997 (
        .y(_T_2375),
        .a(_T_2372),
        .b(_T_2374)
    );
    wire _T_2376;
    BITWISEOR #(.width(1)) bitwiseor_2998 (
        .y(_T_2376),
        .a(_T_2375),
        .b(reset)
    );
    wire _T_2378;
    EQ_UNSIGNED #(.width(1)) u_eq_2999 (
        .y(_T_2378),
        .a(_T_2376),
        .b(1'h0)
    );
    wire _T_2380;
    EQ_UNSIGNED #(.width(1)) u_eq_3000 (
        .y(_T_2380),
        .a(_reg_singleStepped__q),
        .b(1'h0)
    );
    wire _T_2382;
    EQ_UNSIGNED #(.width(1)) u_eq_3001 (
        .y(_T_2382),
        .a(io_retire),
        .b(1'h0)
    );
    wire _T_2383;
    BITWISEOR #(.width(1)) bitwiseor_3002 (
        .y(_T_2383),
        .a(_T_2380),
        .b(_T_2382)
    );
    wire _T_2384;
    BITWISEOR #(.width(1)) bitwiseor_3003 (
        .y(_T_2384),
        .a(_T_2383),
        .b(reset)
    );
    wire _T_2386;
    EQ_UNSIGNED #(.width(1)) u_eq_3004 (
        .y(_T_2386),
        .a(_T_2384),
        .b(1'h0)
    );
    wire [39:0] _T_2387;
    BITWISENOT #(.width(40)) bitwisenot_3005 (
        .y(_T_2387),
        .in(io_pc)
    );
    wire [39:0] _T_2389;
    wire [39:0] _WTEMP_351;
    PAD_UNSIGNED #(.width(1), .n(40)) u_pad_3006 (
        .y(_WTEMP_351),
        .in(1'h1)
    );
    BITWISEOR #(.width(40)) bitwiseor_3007 (
        .y(_T_2389),
        .a(_T_2387),
        .b(_WTEMP_351)
    );
    wire [39:0] _T_2390;
    BITWISENOT #(.width(40)) bitwisenot_3008 (
        .y(_T_2390),
        .in(_T_2389)
    );
    wire [63:0] _T_2391;
    DSHR_UNSIGNED #(.width_in(64), .width_n(2)) u_dshr_3009 (
        .y(_T_2391),
        .in(read_mstatus),
        .n(_reg_mstatus_prv__q)
    );
    wire _T_2392;
    BITS #(.width(64), .high(0), .low(0)) bits_3010 (
        .y(_T_2392),
        .in(_T_2391)
    );
    wire _T_2400;
    wire [63:0] _WTEMP_352;
    PAD_UNSIGNED #(.width(2), .n(64)) u_pad_3011 (
        .y(_WTEMP_352),
        .in(2'h3)
    );
    EQ_UNSIGNED #(.width(64)) u_eq_3012 (
        .y(_T_2400),
        .a(cause),
        .b(_WTEMP_352)
    );
    wire _T_2401;
    wire [63:0] _WTEMP_353;
    PAD_UNSIGNED #(.width(3), .n(64)) u_pad_3013 (
        .y(_WTEMP_353),
        .in(3'h4)
    );
    EQ_UNSIGNED #(.width(64)) u_eq_3014 (
        .y(_T_2401),
        .a(cause),
        .b(_WTEMP_353)
    );
    wire _T_2402;
    wire [63:0] _WTEMP_354;
    PAD_UNSIGNED #(.width(3), .n(64)) u_pad_3015 (
        .y(_WTEMP_354),
        .in(3'h6)
    );
    EQ_UNSIGNED #(.width(64)) u_eq_3016 (
        .y(_T_2402),
        .a(cause),
        .b(_WTEMP_354)
    );
    wire _T_2403;
    wire [63:0] _WTEMP_355;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3017 (
        .y(_WTEMP_355),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(64)) u_eq_3018 (
        .y(_T_2403),
        .a(cause),
        .b(_WTEMP_355)
    );
    wire _T_2404;
    wire [63:0] _WTEMP_356;
    PAD_UNSIGNED #(.width(3), .n(64)) u_pad_3019 (
        .y(_WTEMP_356),
        .in(3'h5)
    );
    EQ_UNSIGNED #(.width(64)) u_eq_3020 (
        .y(_T_2404),
        .a(cause),
        .b(_WTEMP_356)
    );
    wire _T_2405;
    wire [63:0] _WTEMP_357;
    PAD_UNSIGNED #(.width(3), .n(64)) u_pad_3021 (
        .y(_WTEMP_357),
        .in(3'h7)
    );
    EQ_UNSIGNED #(.width(64)) u_eq_3022 (
        .y(_T_2405),
        .a(cause),
        .b(_WTEMP_357)
    );
    wire _T_2406;
    wire [63:0] _WTEMP_358;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3023 (
        .y(_WTEMP_358),
        .in(1'h1)
    );
    EQ_UNSIGNED #(.width(64)) u_eq_3024 (
        .y(_T_2406),
        .a(cause),
        .b(_WTEMP_358)
    );
    wire _T_2407;
    BITWISEOR #(.width(1)) bitwiseor_3025 (
        .y(_T_2407),
        .a(_T_2400),
        .b(_T_2401)
    );
    wire _T_2408;
    BITWISEOR #(.width(1)) bitwiseor_3026 (
        .y(_T_2408),
        .a(_T_2407),
        .b(_T_2402)
    );
    wire _T_2409;
    BITWISEOR #(.width(1)) bitwiseor_3027 (
        .y(_T_2409),
        .a(_T_2408),
        .b(_T_2403)
    );
    wire _T_2410;
    BITWISEOR #(.width(1)) bitwiseor_3028 (
        .y(_T_2410),
        .a(_T_2409),
        .b(_T_2404)
    );
    wire _T_2411;
    BITWISEOR #(.width(1)) bitwiseor_3029 (
        .y(_T_2411),
        .a(_T_2410),
        .b(_T_2405)
    );
    wire _T_2412;
    BITWISEOR #(.width(1)) bitwiseor_3030 (
        .y(_T_2412),
        .a(_T_2411),
        .b(_T_2406)
    );
    wire [1:0] _T_2418;
    wire [1:0] _WTEMP_359;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_3031 (
        .y(_WTEMP_359),
        .in(1'h1)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_3032 (
        .y(_T_2418),
        .sel(causeIsDebugTrigger),
        .a(2'h2),
        .b(_WTEMP_359)
    );
    wire [1:0] _T_2419;
    MUX_UNSIGNED #(.width(2)) u_mux_3033 (
        .y(_T_2419),
        .sel(causeIsDebugInt),
        .a(2'h3),
        .b(_T_2418)
    );
    wire [2:0] _T_2420;
    wire [2:0] _WTEMP_360;
    PAD_UNSIGNED #(.width(2), .n(3)) u_pad_3034 (
        .y(_WTEMP_360),
        .in(_T_2419)
    );
    MUX_UNSIGNED #(.width(3)) u_mux_3035 (
        .y(_T_2420),
        .sel(_reg_singleStepped__q),
        .a(3'h4),
        .b(_WTEMP_360)
    );
    wire _T_2422;
    EQ_UNSIGNED #(.width(1)) u_eq_3036 (
        .y(_T_2422),
        .a(trapToDebug),
        .b(1'h0)
    );
    wire _T_2423;
    BITWISEAND #(.width(1)) bitwiseand_3037 (
        .y(_T_2423),
        .a(_T_2422),
        .b(delegate)
    );
    wire [39:0] _T_2424;
    BITWISENOT #(.width(40)) bitwisenot_3038 (
        .y(_T_2424),
        .in(_T_2390)
    );
    wire _T_2425;
    BITS #(.width(64), .high(2), .low(2)) bits_3039 (
        .y(_T_2425),
        .in(_reg_misa__q)
    );
    wire _T_2427;
    EQ_UNSIGNED #(.width(1)) u_eq_3040 (
        .y(_T_2427),
        .a(_T_2425),
        .b(1'h0)
    );
    wire [1:0] _T_2429;
    CAT #(.width_a(1), .width_b(1)) cat_3041 (
        .y(_T_2429),
        .a(_T_2427),
        .b(1'h1)
    );
    wire [39:0] _T_2430;
    wire [39:0] _WTEMP_361;
    PAD_UNSIGNED #(.width(2), .n(40)) u_pad_3042 (
        .y(_WTEMP_361),
        .in(_T_2429)
    );
    BITWISEOR #(.width(40)) bitwiseor_3043 (
        .y(_T_2430),
        .a(_T_2424),
        .b(_WTEMP_361)
    );
    wire [39:0] _T_2431;
    BITWISENOT #(.width(40)) bitwisenot_3044 (
        .y(_T_2431),
        .in(_T_2430)
    );
    wire [39:0] _node_10;
    MUX_UNSIGNED #(.width(40)) u_mux_3045 (
        .y(_node_10),
        .sel(_T_2412),
        .a(io_badaddr),
        .b(_reg_sbadaddr__q)
    );
    wire _T_2435;
    EQ_UNSIGNED #(.width(1)) u_eq_3046 (
        .y(_T_2435),
        .a(trapToDebug),
        .b(1'h0)
    );
    wire _T_2437;
    EQ_UNSIGNED #(.width(1)) u_eq_3047 (
        .y(_T_2437),
        .a(delegate),
        .b(1'h0)
    );
    wire _T_2438;
    BITWISEAND #(.width(1)) bitwiseand_3048 (
        .y(_T_2438),
        .a(_T_2435),
        .b(_T_2437)
    );
    wire [39:0] _T_2439;
    BITWISENOT #(.width(40)) bitwisenot_3049 (
        .y(_T_2439),
        .in(_T_2390)
    );
    wire _T_2440;
    BITS #(.width(64), .high(2), .low(2)) bits_3050 (
        .y(_T_2440),
        .in(_reg_misa__q)
    );
    wire _T_2442;
    EQ_UNSIGNED #(.width(1)) u_eq_3051 (
        .y(_T_2442),
        .a(_T_2440),
        .b(1'h0)
    );
    wire [1:0] _T_2444;
    CAT #(.width_a(1), .width_b(1)) cat_3052 (
        .y(_T_2444),
        .a(_T_2442),
        .b(1'h1)
    );
    wire [39:0] _T_2445;
    wire [39:0] _WTEMP_362;
    PAD_UNSIGNED #(.width(2), .n(40)) u_pad_3053 (
        .y(_WTEMP_362),
        .in(_T_2444)
    );
    BITWISEOR #(.width(40)) bitwiseor_3054 (
        .y(_T_2445),
        .a(_T_2439),
        .b(_WTEMP_362)
    );
    wire [39:0] _T_2446;
    BITWISENOT #(.width(40)) bitwisenot_3055 (
        .y(_T_2446),
        .in(_T_2445)
    );
    wire [1:0] _node_11;
    wire [1:0] _WTEMP_363;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_3056 (
        .y(_WTEMP_363),
        .in(1'h1)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_3057 (
        .y(_node_11),
        .sel(_T_2423),
        .a(_WTEMP_363),
        .b(_reg_mstatus_prv__q)
    );
    wire [39:0] _node_12;
    MUX_UNSIGNED #(.width(40)) u_mux_3058 (
        .y(_node_12),
        .sel(_T_2412),
        .a(io_badaddr),
        .b(_reg_mbadaddr__q)
    );
    wire [1:0] _node_13;
    MUX_UNSIGNED #(.width(2)) u_mux_3059 (
        .y(_node_13),
        .sel(_T_2438),
        .a(2'h3),
        .b(_node_11)
    );
    wire [2:0] _node_14;
    MUX_UNSIGNED #(.width(3)) u_mux_3060 (
        .y(_node_14),
        .sel(trapToDebug),
        .a(_T_2420),
        .b(_reg_dcsr_cause__q)
    );
    wire [1:0] _node_15;
    MUX_UNSIGNED #(.width(2)) u_mux_3061 (
        .y(_node_15),
        .sel(trapToDebug),
        .a(_reg_mstatus_prv__q),
        .b(_reg_dcsr_prv__q)
    );
    wire _node_16;
    MUX_UNSIGNED #(.width(1)) u_mux_3062 (
        .y(_node_16),
        .sel(trapToDebug),
        .a(1'h1),
        .b(_reg_debug__q)
    );
    wire [39:0] _node_17;
    MUX_UNSIGNED #(.width(40)) u_mux_3063 (
        .y(_node_17),
        .sel(trapToDebug),
        .a(_T_2390),
        .b(_reg_dpc__q)
    );
    wire [39:0] _node_18;
    MUX_UNSIGNED #(.width(40)) u_mux_3064 (
        .y(_node_18),
        .sel(_T_2438),
        .a(_node_12),
        .b(_reg_mbadaddr__q)
    );
    wire [63:0] _node_19;
    MUX_UNSIGNED #(.width(64)) u_mux_3065 (
        .y(_node_19),
        .sel(_T_2438),
        .a(cause),
        .b(_reg_mcause__q)
    );
    wire [39:0] _node_20;
    MUX_UNSIGNED #(.width(40)) u_mux_3066 (
        .y(_node_20),
        .sel(_T_2438),
        .a(_T_2446),
        .b(_reg_mepc__q)
    );
    wire _node_21;
    MUX_UNSIGNED #(.width(1)) u_mux_3067 (
        .y(_node_21),
        .sel(_T_2438),
        .a(1'h0),
        .b(_reg_mstatus_mie__q)
    );
    wire _node_22;
    MUX_UNSIGNED #(.width(1)) u_mux_3068 (
        .y(_node_22),
        .sel(_T_2438),
        .a(_T_2392),
        .b(_reg_mstatus_mpie__q)
    );
    wire [1:0] _node_23;
    MUX_UNSIGNED #(.width(2)) u_mux_3069 (
        .y(_node_23),
        .sel(_T_2438),
        .a(_reg_mstatus_prv__q),
        .b(_reg_mstatus_mpp__q)
    );
    wire _node_24;
    MUX_UNSIGNED #(.width(1)) u_mux_3070 (
        .y(_node_24),
        .sel(_T_2423),
        .a(1'h0),
        .b(_reg_mstatus_sie__q)
    );
    wire _node_25;
    MUX_UNSIGNED #(.width(1)) u_mux_3071 (
        .y(_node_25),
        .sel(_T_2423),
        .a(_T_2392),
        .b(_reg_mstatus_spie__q)
    );
    wire [1:0] _node_26;
    wire [1:0] _WTEMP_364;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_3072 (
        .y(_WTEMP_364),
        .in(_reg_mstatus_spp__q)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_3073 (
        .y(_node_26),
        .sel(_T_2423),
        .a(_reg_mstatus_prv__q),
        .b(_WTEMP_364)
    );
    wire [39:0] _node_27;
    MUX_UNSIGNED #(.width(40)) u_mux_3074 (
        .y(_node_27),
        .sel(_T_2423),
        .a(_node_10),
        .b(_reg_sbadaddr__q)
    );
    wire [63:0] _node_28;
    MUX_UNSIGNED #(.width(64)) u_mux_3075 (
        .y(_node_28),
        .sel(_T_2423),
        .a(cause),
        .b(_reg_scause__q)
    );
    wire [39:0] _node_29;
    MUX_UNSIGNED #(.width(40)) u_mux_3076 (
        .y(_node_29),
        .sel(_T_2423),
        .a(_T_2431),
        .b(_reg_sepc__q)
    );
    wire _T_2450;
    BITS #(.width(12), .high(9), .low(9)) bits_3077 (
        .y(_T_2450),
        .in(io_rw_addr)
    );
    wire _T_2452;
    EQ_UNSIGNED #(.width(1)) u_eq_3078 (
        .y(_T_2452),
        .a(_T_2450),
        .b(1'h0)
    );
    wire _T_2453;
    BITWISEAND #(.width(1)) bitwiseand_3079 (
        .y(_T_2453),
        .a(1'h1),
        .b(_T_2452)
    );
    wire _T_2454;
    BITS #(.width(1), .high(0), .low(0)) bits_3080 (
        .y(_T_2454),
        .in(_reg_mstatus_spp__q)
    );
    wire _node_30;
    MUX_UNSIGNED #(.width(1)) u_mux_3081 (
        .y(_node_30),
        .sel(exception),
        .a(_node_24),
        .b(_reg_mstatus_sie__q)
    );
    wire [1:0] _node_31;
    MUX_UNSIGNED #(.width(2)) u_mux_3082 (
        .y(_node_31),
        .sel(exception),
        .a(_node_13),
        .b(_reg_mstatus_prv__q)
    );
    wire _node_32;
    MUX_UNSIGNED #(.width(1)) u_mux_3083 (
        .y(_node_32),
        .sel(_T_2454),
        .a(_reg_mstatus_spie__q),
        .b(_node_30)
    );
    wire _node_33;
    MUX_UNSIGNED #(.width(1)) u_mux_3084 (
        .y(_node_33),
        .sel(exception),
        .a(_node_24),
        .b(_reg_mstatus_sie__q)
    );
    wire _node_34;
    MUX_UNSIGNED #(.width(1)) u_mux_3085 (
        .y(_node_34),
        .sel(exception),
        .a(_node_25),
        .b(_reg_mstatus_spie__q)
    );
    wire [1:0] _node_35;
    wire [1:0] _WTEMP_365;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_3086 (
        .y(_WTEMP_365),
        .in(_reg_mstatus_spp__q)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_3087 (
        .y(_node_35),
        .sel(exception),
        .a(_node_26),
        .b(_WTEMP_365)
    );
    wire _T_2458;
    BITS #(.width(12), .high(10), .low(10)) bits_3088 (
        .y(_T_2458),
        .in(io_rw_addr)
    );
    wire _T_2459;
    BITWISEAND #(.width(1)) bitwiseand_3089 (
        .y(_T_2459),
        .a(1'h1),
        .b(_T_2458)
    );
    wire _T_2461;
    EQ_UNSIGNED #(.width(1)) u_eq_3090 (
        .y(_T_2461),
        .a(_T_2453),
        .b(1'h0)
    );
    wire _T_2462;
    BITWISEAND #(.width(1)) bitwiseand_3091 (
        .y(_T_2462),
        .a(_T_2461),
        .b(_T_2459)
    );
    wire [39:0] _node_36;
    MUX_UNSIGNED #(.width(40)) u_mux_3092 (
        .y(_node_36),
        .sel(_T_2453),
        .a(_reg_sepc__q),
        .b(tvec)
    );
    wire [1:0] _node_37;
    wire [1:0] _WTEMP_366;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_3093 (
        .y(_WTEMP_366),
        .in(_reg_mstatus_spp__q)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_3094 (
        .y(_node_37),
        .sel(_T_2453),
        .a(_WTEMP_366),
        .b(_node_31)
    );
    wire _node_38;
    MUX_UNSIGNED #(.width(1)) u_mux_3095 (
        .y(_node_38),
        .sel(exception),
        .a(_node_16),
        .b(_reg_debug__q)
    );
    wire _T_2465;
    EQ_UNSIGNED #(.width(1)) u_eq_3096 (
        .y(_T_2465),
        .a(_T_2453),
        .b(1'h0)
    );
    wire _T_2467;
    EQ_UNSIGNED #(.width(1)) u_eq_3097 (
        .y(_T_2467),
        .a(_T_2459),
        .b(1'h0)
    );
    wire _T_2468;
    BITWISEAND #(.width(1)) bitwiseand_3098 (
        .y(_T_2468),
        .a(_T_2465),
        .b(_T_2467)
    );
    wire _T_2469;
    BITS #(.width(2), .high(1), .low(1)) bits_3099 (
        .y(_T_2469),
        .in(_reg_mstatus_mpp__q)
    );
    wire _node_39;
    MUX_UNSIGNED #(.width(1)) u_mux_3100 (
        .y(_node_39),
        .sel(exception),
        .a(_node_21),
        .b(_reg_mstatus_mie__q)
    );
    wire _T_2471;
    BITS #(.width(2), .high(0), .low(0)) bits_3101 (
        .y(_T_2471),
        .in(_reg_mstatus_mpp__q)
    );
    wire _T_2472;
    BITWISEAND #(.width(1)) bitwiseand_3102 (
        .y(_T_2472),
        .a(1'h1),
        .b(_T_2471)
    );
    wire _T_2474;
    EQ_UNSIGNED #(.width(1)) u_eq_3103 (
        .y(_T_2474),
        .a(_T_2469),
        .b(1'h0)
    );
    wire _T_2475;
    BITWISEAND #(.width(1)) bitwiseand_3104 (
        .y(_T_2475),
        .a(_T_2474),
        .b(_T_2472)
    );
    wire _node_40;
    MUX_UNSIGNED #(.width(1)) u_mux_3105 (
        .y(_node_40),
        .sel(_T_2453),
        .a(_node_32),
        .b(_node_33)
    );
    wire _T_2479;
    assign _T_2479 = 1'h0;
    wire _T_2481;
    assign _T_2481 = 1'h0;
    wire [39:0] _node_41;
    MUX_UNSIGNED #(.width(40)) u_mux_3106 (
        .y(_node_41),
        .sel(_T_2462),
        .a(_reg_dpc__q),
        .b(_node_36)
    );
    wire [1:0] _node_42;
    MUX_UNSIGNED #(.width(2)) u_mux_3107 (
        .y(_node_42),
        .sel(_T_2462),
        .a(_reg_dcsr_prv__q),
        .b(_node_37)
    );
    wire _node_43;
    MUX_UNSIGNED #(.width(1)) u_mux_3108 (
        .y(_node_43),
        .sel(_T_2469),
        .a(_reg_mstatus_mpie__q),
        .b(_node_39)
    );
    wire _node_44;
    MUX_UNSIGNED #(.width(1)) u_mux_3109 (
        .y(_node_44),
        .sel(exception),
        .a(_node_21),
        .b(_reg_mstatus_mie__q)
    );
    wire _node_45;
    MUX_UNSIGNED #(.width(1)) u_mux_3110 (
        .y(_node_45),
        .sel(exception),
        .a(_node_22),
        .b(_reg_mstatus_mpie__q)
    );
    wire [1:0] _node_46;
    MUX_UNSIGNED #(.width(2)) u_mux_3111 (
        .y(_node_46),
        .sel(exception),
        .a(_node_23),
        .b(_reg_mstatus_mpp__q)
    );
    wire _node_47;
    MUX_UNSIGNED #(.width(1)) u_mux_3112 (
        .y(_node_47),
        .sel(_T_2475),
        .a(_reg_mstatus_mpie__q),
        .b(_node_40)
    );
    wire _node_48;
    MUX_UNSIGNED #(.width(1)) u_mux_3113 (
        .y(_node_48),
        .sel(_T_2453),
        .a(_node_32),
        .b(_node_33)
    );
    wire [39:0] _node_49;
    MUX_UNSIGNED #(.width(40)) u_mux_3114 (
        .y(_node_49),
        .sel(_T_2468),
        .a(_reg_mepc__q),
        .b(_node_41)
    );
    wire [1:0] _node_50;
    MUX_UNSIGNED #(.width(2)) u_mux_3115 (
        .y(_node_50),
        .sel(_T_2468),
        .a(_reg_mstatus_mpp__q),
        .b(_node_42)
    );
    wire [1:0] _node_51;
    MUX_UNSIGNED #(.width(2)) u_mux_3116 (
        .y(_node_51),
        .sel(exception),
        .a(_node_13),
        .b(_reg_mstatus_prv__q)
    );
    wire _node_52;
    MUX_UNSIGNED #(.width(1)) u_mux_3117 (
        .y(_node_52),
        .sel(_T_2462),
        .a(1'h0),
        .b(_node_38)
    );
    wire _node_53;
    MUX_UNSIGNED #(.width(1)) u_mux_3118 (
        .y(_node_53),
        .sel(exception),
        .a(_node_16),
        .b(_reg_debug__q)
    );
    wire _node_54;
    MUX_UNSIGNED #(.width(1)) u_mux_3119 (
        .y(_node_54),
        .sel(_T_2468),
        .a(_node_43),
        .b(_node_44)
    );
    wire _node_55;
    MUX_UNSIGNED #(.width(1)) u_mux_3120 (
        .y(_node_55),
        .sel(exception),
        .a(_node_21),
        .b(_reg_mstatus_mie__q)
    );
    wire _node_56;
    MUX_UNSIGNED #(.width(1)) u_mux_3121 (
        .y(_node_56),
        .sel(_T_2468),
        .a(1'h1),
        .b(_node_45)
    );
    wire _node_57;
    MUX_UNSIGNED #(.width(1)) u_mux_3122 (
        .y(_node_57),
        .sel(exception),
        .a(_node_22),
        .b(_reg_mstatus_mpie__q)
    );
    wire [1:0] _node_58;
    wire [1:0] _WTEMP_367;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_3123 (
        .y(_WTEMP_367),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_3124 (
        .y(_node_58),
        .sel(_T_2468),
        .a(_WTEMP_367),
        .b(_node_46)
    );
    wire [1:0] _node_59;
    MUX_UNSIGNED #(.width(2)) u_mux_3125 (
        .y(_node_59),
        .sel(exception),
        .a(_node_23),
        .b(_reg_mstatus_mpp__q)
    );
    wire _node_60;
    MUX_UNSIGNED #(.width(1)) u_mux_3126 (
        .y(_node_60),
        .sel(_T_2468),
        .a(_node_47),
        .b(_node_48)
    );
    wire _node_61;
    MUX_UNSIGNED #(.width(1)) u_mux_3127 (
        .y(_node_61),
        .sel(exception),
        .a(_node_24),
        .b(_reg_mstatus_sie__q)
    );
    wire _node_62;
    MUX_UNSIGNED #(.width(1)) u_mux_3128 (
        .y(_node_62),
        .sel(_T_2453),
        .a(1'h1),
        .b(_node_34)
    );
    wire _node_63;
    MUX_UNSIGNED #(.width(1)) u_mux_3129 (
        .y(_node_63),
        .sel(exception),
        .a(_node_25),
        .b(_reg_mstatus_spie__q)
    );
    wire [1:0] _node_64;
    wire [1:0] _WTEMP_368;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_3130 (
        .y(_WTEMP_368),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_3131 (
        .y(_node_64),
        .sel(_T_2453),
        .a(_WTEMP_368),
        .b(_node_35)
    );
    wire [1:0] _node_65;
    wire [1:0] _WTEMP_369;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_3132 (
        .y(_WTEMP_369),
        .in(_reg_mstatus_spp__q)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_3133 (
        .y(_node_65),
        .sel(exception),
        .a(_node_26),
        .b(_WTEMP_369)
    );
    wire _T_2483;
    assign _T_2483 = 1'h0;
    wire [63:0] _T_2485;
    wire [63:0] _WTEMP_370;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3134 (
        .y(_WTEMP_370),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_3135 (
        .y(_T_2485),
        .sel(_T_1469),
        .a(_T_1304),
        .b(_WTEMP_370)
    );
    wire [63:0] _T_2487;
    wire [63:0] _WTEMP_371;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3136 (
        .y(_WTEMP_371),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_3137 (
        .y(_T_2487),
        .sel(_T_1471),
        .a(_T_1345),
        .b(_WTEMP_371)
    );
    wire _T_2489;
    assign _T_2489 = 1'h0;
    wire _T_2491;
    assign _T_2491 = 1'h0;
    wire _T_2493;
    assign _T_2493 = 1'h0;
    wire [63:0] _T_2495;
    wire [63:0] _WTEMP_372;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3138 (
        .y(_WTEMP_372),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_3139 (
        .y(_T_2495),
        .sel(_T_1479),
        .a(_T_950),
        .b(_WTEMP_372)
    );
    wire [63:0] _T_2497;
    wire [63:0] _WTEMP_373;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3140 (
        .y(_WTEMP_373),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_3141 (
        .y(_T_2497),
        .sel(_T_1481),
        .a(_T_939),
        .b(_WTEMP_373)
    );
    wire [63:0] _T_2499;
    wire [63:0] _WTEMP_374;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3142 (
        .y(_WTEMP_374),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_3143 (
        .y(_T_2499),
        .sel(_T_1483),
        .a(_reg_misa__q),
        .b(_WTEMP_374)
    );
    wire [63:0] _T_2501;
    wire [63:0] _WTEMP_375;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3144 (
        .y(_WTEMP_375),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_3145 (
        .y(_T_2501),
        .sel(_T_1485),
        .a(read_mstatus),
        .b(_WTEMP_375)
    );
    wire [31:0] _T_2503;
    wire [31:0] _WTEMP_376;
    PAD_UNSIGNED #(.width(1), .n(32)) u_pad_3146 (
        .y(_WTEMP_376),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(32)) u_mux_3147 (
        .y(_T_2503),
        .sel(_T_1487),
        .a(_reg_mtvec__q),
        .b(_WTEMP_376)
    );
    wire [12:0] _T_2505;
    wire [12:0] _WTEMP_377;
    PAD_UNSIGNED #(.width(1), .n(13)) u_pad_3148 (
        .y(_WTEMP_377),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(13)) u_mux_3149 (
        .y(_T_2505),
        .sel(_T_1489),
        .a(read_mip),
        .b(_WTEMP_377)
    );
    wire [63:0] _T_2507;
    wire [63:0] _WTEMP_378;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3150 (
        .y(_WTEMP_378),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_3151 (
        .y(_T_2507),
        .sel(_T_1491),
        .a(_reg_mie__q),
        .b(_WTEMP_378)
    );
    wire [63:0] _T_2509;
    wire [63:0] _WTEMP_379;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3152 (
        .y(_WTEMP_379),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_3153 (
        .y(_T_2509),
        .sel(_T_1493),
        .a(_reg_mideleg__q),
        .b(_WTEMP_379)
    );
    wire [63:0] _T_2511;
    wire [63:0] _WTEMP_380;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3154 (
        .y(_WTEMP_380),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_3155 (
        .y(_T_2511),
        .sel(_T_1495),
        .a(_reg_medeleg__q),
        .b(_WTEMP_380)
    );
    wire [63:0] _T_2513;
    wire [63:0] _WTEMP_381;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3156 (
        .y(_WTEMP_381),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_3157 (
        .y(_T_2513),
        .sel(_T_1497),
        .a(_reg_mscratch__q),
        .b(_WTEMP_381)
    );
    wire [63:0] _T_2515;
    wire [63:0] _WTEMP_382;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3158 (
        .y(_WTEMP_382),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_3159 (
        .y(_T_2515),
        .sel(_T_1499),
        .a(_T_1354),
        .b(_WTEMP_382)
    );
    wire [63:0] _T_2517;
    wire [63:0] _WTEMP_383;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3160 (
        .y(_WTEMP_383),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_3161 (
        .y(_T_2517),
        .sel(_T_1501),
        .a(_T_1360),
        .b(_WTEMP_383)
    );
    wire [63:0] _T_2519;
    wire [63:0] _WTEMP_384;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3162 (
        .y(_WTEMP_384),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_3163 (
        .y(_T_2519),
        .sel(_T_1503),
        .a(_reg_mcause__q),
        .b(_WTEMP_384)
    );
    wire [63:0] _T_2521;
    wire [63:0] _WTEMP_385;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3164 (
        .y(_WTEMP_385),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_3165 (
        .y(_T_2521),
        .sel(_T_1505),
        .a(io_hartid),
        .b(_WTEMP_385)
    );
    wire [31:0] _T_2523;
    wire [31:0] _WTEMP_386;
    PAD_UNSIGNED #(.width(1), .n(32)) u_pad_3166 (
        .y(_WTEMP_386),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(32)) u_mux_3167 (
        .y(_T_2523),
        .sel(_T_1507),
        .a(_T_1376),
        .b(_WTEMP_386)
    );
    wire [39:0] _T_2525;
    wire [39:0] _WTEMP_387;
    PAD_UNSIGNED #(.width(1), .n(40)) u_pad_3168 (
        .y(_WTEMP_387),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(40)) u_mux_3169 (
        .y(_T_2525),
        .sel(_T_1509),
        .a(_reg_dpc__q),
        .b(_WTEMP_387)
    );
    wire [63:0] _T_2527;
    wire [63:0] _WTEMP_388;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3170 (
        .y(_WTEMP_388),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_3171 (
        .y(_T_2527),
        .sel(_T_1511),
        .a(_reg_dscratch__q),
        .b(_WTEMP_388)
    );
    wire [4:0] _T_2529;
    wire [4:0] _WTEMP_389;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_3172 (
        .y(_WTEMP_389),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(5)) u_mux_3173 (
        .y(_T_2529),
        .sel(_T_1513),
        .a(_reg_fflags__q),
        .b(_WTEMP_389)
    );
    wire [2:0] _T_2531;
    wire [2:0] _WTEMP_390;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_3174 (
        .y(_WTEMP_390),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(3)) u_mux_3175 (
        .y(_T_2531),
        .sel(_T_1515),
        .a(_reg_frm__q),
        .b(_WTEMP_390)
    );
    wire [7:0] _T_2533;
    wire [7:0] _WTEMP_391;
    PAD_UNSIGNED #(.width(1), .n(8)) u_pad_3176 (
        .y(_WTEMP_391),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(8)) u_mux_3177 (
        .y(_T_2533),
        .sel(_T_1517),
        .a(_T_1377),
        .b(_WTEMP_391)
    );
    wire _T_2535;
    assign _T_2535 = 1'h0;
    wire _T_2537;
    assign _T_2537 = 1'h0;
    wire _T_2539;
    assign _T_2539 = 1'h0;
    wire _T_2541;
    assign _T_2541 = 1'h0;
    wire _T_2543;
    assign _T_2543 = 1'h0;
    wire _T_2545;
    assign _T_2545 = 1'h0;
    wire _T_2547;
    assign _T_2547 = 1'h0;
    wire _T_2549;
    assign _T_2549 = 1'h0;
    wire _T_2551;
    assign _T_2551 = 1'h0;
    wire _T_2553;
    assign _T_2553 = 1'h0;
    wire _T_2555;
    assign _T_2555 = 1'h0;
    wire _T_2557;
    assign _T_2557 = 1'h0;
    wire _T_2559;
    assign _T_2559 = 1'h0;
    wire _T_2561;
    assign _T_2561 = 1'h0;
    wire _T_2563;
    assign _T_2563 = 1'h0;
    wire _T_2565;
    assign _T_2565 = 1'h0;
    wire _T_2567;
    assign _T_2567 = 1'h0;
    wire _T_2569;
    assign _T_2569 = 1'h0;
    wire _T_2571;
    assign _T_2571 = 1'h0;
    wire _T_2573;
    assign _T_2573 = 1'h0;
    wire _T_2575;
    assign _T_2575 = 1'h0;
    wire _T_2577;
    assign _T_2577 = 1'h0;
    wire _T_2579;
    assign _T_2579 = 1'h0;
    wire _T_2581;
    assign _T_2581 = 1'h0;
    wire _T_2583;
    assign _T_2583 = 1'h0;
    wire _T_2585;
    assign _T_2585 = 1'h0;
    wire _T_2587;
    assign _T_2587 = 1'h0;
    wire _T_2589;
    assign _T_2589 = 1'h0;
    wire _T_2591;
    assign _T_2591 = 1'h0;
    wire _T_2593;
    assign _T_2593 = 1'h0;
    wire _T_2595;
    assign _T_2595 = 1'h0;
    wire _T_2597;
    assign _T_2597 = 1'h0;
    wire _T_2599;
    assign _T_2599 = 1'h0;
    wire _T_2601;
    assign _T_2601 = 1'h0;
    wire _T_2603;
    assign _T_2603 = 1'h0;
    wire _T_2605;
    assign _T_2605 = 1'h0;
    wire _T_2607;
    assign _T_2607 = 1'h0;
    wire _T_2609;
    assign _T_2609 = 1'h0;
    wire _T_2611;
    assign _T_2611 = 1'h0;
    wire _T_2613;
    assign _T_2613 = 1'h0;
    wire _T_2615;
    assign _T_2615 = 1'h0;
    wire _T_2617;
    assign _T_2617 = 1'h0;
    wire _T_2619;
    assign _T_2619 = 1'h0;
    wire _T_2621;
    assign _T_2621 = 1'h0;
    wire _T_2623;
    assign _T_2623 = 1'h0;
    wire _T_2625;
    assign _T_2625 = 1'h0;
    wire _T_2627;
    assign _T_2627 = 1'h0;
    wire _T_2629;
    assign _T_2629 = 1'h0;
    wire _T_2631;
    assign _T_2631 = 1'h0;
    wire _T_2633;
    assign _T_2633 = 1'h0;
    wire _T_2635;
    assign _T_2635 = 1'h0;
    wire _T_2637;
    assign _T_2637 = 1'h0;
    wire _T_2639;
    assign _T_2639 = 1'h0;
    wire _T_2641;
    assign _T_2641 = 1'h0;
    wire _T_2643;
    assign _T_2643 = 1'h0;
    wire _T_2645;
    assign _T_2645 = 1'h0;
    wire _T_2647;
    assign _T_2647 = 1'h0;
    wire _T_2649;
    assign _T_2649 = 1'h0;
    wire _T_2651;
    assign _T_2651 = 1'h0;
    wire _T_2653;
    assign _T_2653 = 1'h0;
    wire _T_2655;
    assign _T_2655 = 1'h0;
    wire _T_2657;
    assign _T_2657 = 1'h0;
    wire _T_2659;
    assign _T_2659 = 1'h0;
    wire _T_2661;
    assign _T_2661 = 1'h0;
    wire _T_2663;
    assign _T_2663 = 1'h0;
    wire _T_2665;
    assign _T_2665 = 1'h0;
    wire _T_2667;
    assign _T_2667 = 1'h0;
    wire _T_2669;
    assign _T_2669 = 1'h0;
    wire _T_2671;
    assign _T_2671 = 1'h0;
    wire _T_2673;
    assign _T_2673 = 1'h0;
    wire _T_2675;
    assign _T_2675 = 1'h0;
    wire _T_2677;
    assign _T_2677 = 1'h0;
    wire _T_2679;
    assign _T_2679 = 1'h0;
    wire _T_2681;
    assign _T_2681 = 1'h0;
    wire _T_2683;
    assign _T_2683 = 1'h0;
    wire _T_2685;
    assign _T_2685 = 1'h0;
    wire _T_2687;
    assign _T_2687 = 1'h0;
    wire _T_2689;
    assign _T_2689 = 1'h0;
    wire _T_2691;
    assign _T_2691 = 1'h0;
    wire _T_2693;
    assign _T_2693 = 1'h0;
    wire _T_2695;
    assign _T_2695 = 1'h0;
    wire _T_2697;
    assign _T_2697 = 1'h0;
    wire _T_2699;
    assign _T_2699 = 1'h0;
    wire _T_2701;
    assign _T_2701 = 1'h0;
    wire _T_2703;
    assign _T_2703 = 1'h0;
    wire _T_2705;
    assign _T_2705 = 1'h0;
    wire _T_2707;
    assign _T_2707 = 1'h0;
    wire [63:0] _T_2709;
    wire [63:0] _WTEMP_392;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3178 (
        .y(_WTEMP_392),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_3179 (
        .y(_T_2709),
        .sel(_T_1693),
        .a(_T_1445),
        .b(_WTEMP_392)
    );
    wire [63:0] _T_2711;
    wire [63:0] _WTEMP_393;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3180 (
        .y(_WTEMP_393),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_3181 (
        .y(_T_2711),
        .sel(_T_1695),
        .a(_T_1381),
        .b(_WTEMP_393)
    );
    wire [63:0] _T_2713;
    wire [63:0] _WTEMP_394;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3182 (
        .y(_WTEMP_394),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_3183 (
        .y(_T_2713),
        .sel(_T_1697),
        .a(_T_1380),
        .b(_WTEMP_394)
    );
    wire [63:0] _T_2715;
    wire [63:0] _WTEMP_395;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3184 (
        .y(_WTEMP_395),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_3185 (
        .y(_T_2715),
        .sel(_T_1699),
        .a(_reg_sscratch__q),
        .b(_WTEMP_395)
    );
    wire [63:0] _T_2717;
    wire [63:0] _WTEMP_396;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3186 (
        .y(_WTEMP_396),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_3187 (
        .y(_T_2717),
        .sel(_T_1701),
        .a(_reg_scause__q),
        .b(_WTEMP_396)
    );
    wire [63:0] _T_2719;
    wire [63:0] _WTEMP_397;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3188 (
        .y(_WTEMP_397),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_3189 (
        .y(_T_2719),
        .sel(_T_1703),
        .a(_T_1451),
        .b(_WTEMP_397)
    );
    wire [63:0] _T_2721;
    wire [63:0] _WTEMP_398;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3190 (
        .y(_WTEMP_398),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_3191 (
        .y(_T_2721),
        .sel(_T_1705),
        .a(_T_1453),
        .b(_WTEMP_398)
    );
    wire [63:0] _T_2723;
    wire [63:0] _WTEMP_399;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3192 (
        .y(_WTEMP_399),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_3193 (
        .y(_T_2723),
        .sel(_T_1707),
        .a(_T_1459),
        .b(_WTEMP_399)
    );
    wire [63:0] _T_2725;
    wire [63:0] _WTEMP_400;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3194 (
        .y(_WTEMP_400),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_3195 (
        .y(_T_2725),
        .sel(_T_1709),
        .a(_T_1465),
        .b(_WTEMP_400)
    );
    wire [31:0] _T_2727;
    wire [31:0] _WTEMP_401;
    PAD_UNSIGNED #(.width(1), .n(32)) u_pad_3196 (
        .y(_WTEMP_401),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(32)) u_mux_3197 (
        .y(_T_2727),
        .sel(_T_1711),
        .a(_reg_scounteren__q),
        .b(_WTEMP_401)
    );
    wire [31:0] _T_2729;
    wire [31:0] _WTEMP_402;
    PAD_UNSIGNED #(.width(1), .n(32)) u_pad_3198 (
        .y(_WTEMP_402),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(32)) u_mux_3199 (
        .y(_T_2729),
        .sel(_T_1713),
        .a(_reg_mcounteren__q),
        .b(_WTEMP_402)
    );
    wire [63:0] _T_2731;
    wire [63:0] _WTEMP_403;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3200 (
        .y(_WTEMP_403),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_3201 (
        .y(_T_2731),
        .sel(_T_1715),
        .a(_T_950),
        .b(_WTEMP_403)
    );
    wire [63:0] _T_2733;
    wire [63:0] _WTEMP_404;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3202 (
        .y(_WTEMP_404),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_3203 (
        .y(_T_2733),
        .sel(_T_1717),
        .a(_T_939),
        .b(_WTEMP_404)
    );
    wire [63:0] _T_2735;
    wire [63:0] _WTEMP_405;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3204 (
        .y(_WTEMP_405),
        .in(_T_2483)
    );
    BITWISEOR #(.width(64)) bitwiseor_3205 (
        .y(_T_2735),
        .a(_WTEMP_405),
        .b(_T_2485)
    );
    wire [63:0] _T_2736;
    BITWISEOR #(.width(64)) bitwiseor_3206 (
        .y(_T_2736),
        .a(_T_2735),
        .b(_T_2487)
    );
    wire [63:0] _T_2737;
    wire [63:0] _WTEMP_406;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3207 (
        .y(_WTEMP_406),
        .in(_T_2489)
    );
    BITWISEOR #(.width(64)) bitwiseor_3208 (
        .y(_T_2737),
        .a(_T_2736),
        .b(_WTEMP_406)
    );
    wire [63:0] _T_2738;
    wire [63:0] _WTEMP_407;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3209 (
        .y(_WTEMP_407),
        .in(_T_2491)
    );
    BITWISEOR #(.width(64)) bitwiseor_3210 (
        .y(_T_2738),
        .a(_T_2737),
        .b(_WTEMP_407)
    );
    wire [63:0] _T_2739;
    wire [63:0] _WTEMP_408;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3211 (
        .y(_WTEMP_408),
        .in(_T_2493)
    );
    BITWISEOR #(.width(64)) bitwiseor_3212 (
        .y(_T_2739),
        .a(_T_2738),
        .b(_WTEMP_408)
    );
    wire [63:0] _T_2740;
    BITWISEOR #(.width(64)) bitwiseor_3213 (
        .y(_T_2740),
        .a(_T_2739),
        .b(_T_2495)
    );
    wire [63:0] _T_2741;
    BITWISEOR #(.width(64)) bitwiseor_3214 (
        .y(_T_2741),
        .a(_T_2740),
        .b(_T_2497)
    );
    wire [63:0] _T_2742;
    BITWISEOR #(.width(64)) bitwiseor_3215 (
        .y(_T_2742),
        .a(_T_2741),
        .b(_T_2499)
    );
    wire [63:0] _T_2743;
    BITWISEOR #(.width(64)) bitwiseor_3216 (
        .y(_T_2743),
        .a(_T_2742),
        .b(_T_2501)
    );
    wire [63:0] _T_2744;
    wire [63:0] _WTEMP_409;
    PAD_UNSIGNED #(.width(32), .n(64)) u_pad_3217 (
        .y(_WTEMP_409),
        .in(_T_2503)
    );
    BITWISEOR #(.width(64)) bitwiseor_3218 (
        .y(_T_2744),
        .a(_T_2743),
        .b(_WTEMP_409)
    );
    wire [63:0] _T_2745;
    wire [63:0] _WTEMP_410;
    PAD_UNSIGNED #(.width(13), .n(64)) u_pad_3219 (
        .y(_WTEMP_410),
        .in(_T_2505)
    );
    BITWISEOR #(.width(64)) bitwiseor_3220 (
        .y(_T_2745),
        .a(_T_2744),
        .b(_WTEMP_410)
    );
    wire [63:0] _T_2746;
    BITWISEOR #(.width(64)) bitwiseor_3221 (
        .y(_T_2746),
        .a(_T_2745),
        .b(_T_2507)
    );
    wire [63:0] _T_2747;
    BITWISEOR #(.width(64)) bitwiseor_3222 (
        .y(_T_2747),
        .a(_T_2746),
        .b(_T_2509)
    );
    wire [63:0] _T_2748;
    BITWISEOR #(.width(64)) bitwiseor_3223 (
        .y(_T_2748),
        .a(_T_2747),
        .b(_T_2511)
    );
    wire [63:0] _T_2749;
    BITWISEOR #(.width(64)) bitwiseor_3224 (
        .y(_T_2749),
        .a(_T_2748),
        .b(_T_2513)
    );
    wire [63:0] _T_2750;
    BITWISEOR #(.width(64)) bitwiseor_3225 (
        .y(_T_2750),
        .a(_T_2749),
        .b(_T_2515)
    );
    wire [63:0] _T_2751;
    BITWISEOR #(.width(64)) bitwiseor_3226 (
        .y(_T_2751),
        .a(_T_2750),
        .b(_T_2517)
    );
    wire [63:0] _T_2752;
    BITWISEOR #(.width(64)) bitwiseor_3227 (
        .y(_T_2752),
        .a(_T_2751),
        .b(_T_2519)
    );
    wire [63:0] _T_2753;
    BITWISEOR #(.width(64)) bitwiseor_3228 (
        .y(_T_2753),
        .a(_T_2752),
        .b(_T_2521)
    );
    wire [63:0] _T_2754;
    wire [63:0] _WTEMP_411;
    PAD_UNSIGNED #(.width(32), .n(64)) u_pad_3229 (
        .y(_WTEMP_411),
        .in(_T_2523)
    );
    BITWISEOR #(.width(64)) bitwiseor_3230 (
        .y(_T_2754),
        .a(_T_2753),
        .b(_WTEMP_411)
    );
    wire [63:0] _T_2755;
    wire [63:0] _WTEMP_412;
    PAD_UNSIGNED #(.width(40), .n(64)) u_pad_3231 (
        .y(_WTEMP_412),
        .in(_T_2525)
    );
    BITWISEOR #(.width(64)) bitwiseor_3232 (
        .y(_T_2755),
        .a(_T_2754),
        .b(_WTEMP_412)
    );
    wire [63:0] _T_2756;
    BITWISEOR #(.width(64)) bitwiseor_3233 (
        .y(_T_2756),
        .a(_T_2755),
        .b(_T_2527)
    );
    wire [63:0] _T_2757;
    wire [63:0] _WTEMP_413;
    PAD_UNSIGNED #(.width(5), .n(64)) u_pad_3234 (
        .y(_WTEMP_413),
        .in(_T_2529)
    );
    BITWISEOR #(.width(64)) bitwiseor_3235 (
        .y(_T_2757),
        .a(_T_2756),
        .b(_WTEMP_413)
    );
    wire [63:0] _T_2758;
    wire [63:0] _WTEMP_414;
    PAD_UNSIGNED #(.width(3), .n(64)) u_pad_3236 (
        .y(_WTEMP_414),
        .in(_T_2531)
    );
    BITWISEOR #(.width(64)) bitwiseor_3237 (
        .y(_T_2758),
        .a(_T_2757),
        .b(_WTEMP_414)
    );
    wire [63:0] _T_2759;
    wire [63:0] _WTEMP_415;
    PAD_UNSIGNED #(.width(8), .n(64)) u_pad_3238 (
        .y(_WTEMP_415),
        .in(_T_2533)
    );
    BITWISEOR #(.width(64)) bitwiseor_3239 (
        .y(_T_2759),
        .a(_T_2758),
        .b(_WTEMP_415)
    );
    wire [63:0] _T_2760;
    wire [63:0] _WTEMP_416;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3240 (
        .y(_WTEMP_416),
        .in(_T_2535)
    );
    BITWISEOR #(.width(64)) bitwiseor_3241 (
        .y(_T_2760),
        .a(_T_2759),
        .b(_WTEMP_416)
    );
    wire [63:0] _T_2761;
    wire [63:0] _WTEMP_417;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3242 (
        .y(_WTEMP_417),
        .in(_T_2537)
    );
    BITWISEOR #(.width(64)) bitwiseor_3243 (
        .y(_T_2761),
        .a(_T_2760),
        .b(_WTEMP_417)
    );
    wire [63:0] _T_2762;
    wire [63:0] _WTEMP_418;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3244 (
        .y(_WTEMP_418),
        .in(_T_2539)
    );
    BITWISEOR #(.width(64)) bitwiseor_3245 (
        .y(_T_2762),
        .a(_T_2761),
        .b(_WTEMP_418)
    );
    wire [63:0] _T_2763;
    wire [63:0] _WTEMP_419;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3246 (
        .y(_WTEMP_419),
        .in(_T_2541)
    );
    BITWISEOR #(.width(64)) bitwiseor_3247 (
        .y(_T_2763),
        .a(_T_2762),
        .b(_WTEMP_419)
    );
    wire [63:0] _T_2764;
    wire [63:0] _WTEMP_420;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3248 (
        .y(_WTEMP_420),
        .in(_T_2543)
    );
    BITWISEOR #(.width(64)) bitwiseor_3249 (
        .y(_T_2764),
        .a(_T_2763),
        .b(_WTEMP_420)
    );
    wire [63:0] _T_2765;
    wire [63:0] _WTEMP_421;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3250 (
        .y(_WTEMP_421),
        .in(_T_2545)
    );
    BITWISEOR #(.width(64)) bitwiseor_3251 (
        .y(_T_2765),
        .a(_T_2764),
        .b(_WTEMP_421)
    );
    wire [63:0] _T_2766;
    wire [63:0] _WTEMP_422;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3252 (
        .y(_WTEMP_422),
        .in(_T_2547)
    );
    BITWISEOR #(.width(64)) bitwiseor_3253 (
        .y(_T_2766),
        .a(_T_2765),
        .b(_WTEMP_422)
    );
    wire [63:0] _T_2767;
    wire [63:0] _WTEMP_423;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3254 (
        .y(_WTEMP_423),
        .in(_T_2549)
    );
    BITWISEOR #(.width(64)) bitwiseor_3255 (
        .y(_T_2767),
        .a(_T_2766),
        .b(_WTEMP_423)
    );
    wire [63:0] _T_2768;
    wire [63:0] _WTEMP_424;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3256 (
        .y(_WTEMP_424),
        .in(_T_2551)
    );
    BITWISEOR #(.width(64)) bitwiseor_3257 (
        .y(_T_2768),
        .a(_T_2767),
        .b(_WTEMP_424)
    );
    wire [63:0] _T_2769;
    wire [63:0] _WTEMP_425;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3258 (
        .y(_WTEMP_425),
        .in(_T_2553)
    );
    BITWISEOR #(.width(64)) bitwiseor_3259 (
        .y(_T_2769),
        .a(_T_2768),
        .b(_WTEMP_425)
    );
    wire [63:0] _T_2770;
    wire [63:0] _WTEMP_426;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3260 (
        .y(_WTEMP_426),
        .in(_T_2555)
    );
    BITWISEOR #(.width(64)) bitwiseor_3261 (
        .y(_T_2770),
        .a(_T_2769),
        .b(_WTEMP_426)
    );
    wire [63:0] _T_2771;
    wire [63:0] _WTEMP_427;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3262 (
        .y(_WTEMP_427),
        .in(_T_2557)
    );
    BITWISEOR #(.width(64)) bitwiseor_3263 (
        .y(_T_2771),
        .a(_T_2770),
        .b(_WTEMP_427)
    );
    wire [63:0] _T_2772;
    wire [63:0] _WTEMP_428;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3264 (
        .y(_WTEMP_428),
        .in(_T_2559)
    );
    BITWISEOR #(.width(64)) bitwiseor_3265 (
        .y(_T_2772),
        .a(_T_2771),
        .b(_WTEMP_428)
    );
    wire [63:0] _T_2773;
    wire [63:0] _WTEMP_429;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3266 (
        .y(_WTEMP_429),
        .in(_T_2561)
    );
    BITWISEOR #(.width(64)) bitwiseor_3267 (
        .y(_T_2773),
        .a(_T_2772),
        .b(_WTEMP_429)
    );
    wire [63:0] _T_2774;
    wire [63:0] _WTEMP_430;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3268 (
        .y(_WTEMP_430),
        .in(_T_2563)
    );
    BITWISEOR #(.width(64)) bitwiseor_3269 (
        .y(_T_2774),
        .a(_T_2773),
        .b(_WTEMP_430)
    );
    wire [63:0] _T_2775;
    wire [63:0] _WTEMP_431;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3270 (
        .y(_WTEMP_431),
        .in(_T_2565)
    );
    BITWISEOR #(.width(64)) bitwiseor_3271 (
        .y(_T_2775),
        .a(_T_2774),
        .b(_WTEMP_431)
    );
    wire [63:0] _T_2776;
    wire [63:0] _WTEMP_432;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3272 (
        .y(_WTEMP_432),
        .in(_T_2567)
    );
    BITWISEOR #(.width(64)) bitwiseor_3273 (
        .y(_T_2776),
        .a(_T_2775),
        .b(_WTEMP_432)
    );
    wire [63:0] _T_2777;
    wire [63:0] _WTEMP_433;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3274 (
        .y(_WTEMP_433),
        .in(_T_2569)
    );
    BITWISEOR #(.width(64)) bitwiseor_3275 (
        .y(_T_2777),
        .a(_T_2776),
        .b(_WTEMP_433)
    );
    wire [63:0] _T_2778;
    wire [63:0] _WTEMP_434;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3276 (
        .y(_WTEMP_434),
        .in(_T_2571)
    );
    BITWISEOR #(.width(64)) bitwiseor_3277 (
        .y(_T_2778),
        .a(_T_2777),
        .b(_WTEMP_434)
    );
    wire [63:0] _T_2779;
    wire [63:0] _WTEMP_435;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3278 (
        .y(_WTEMP_435),
        .in(_T_2573)
    );
    BITWISEOR #(.width(64)) bitwiseor_3279 (
        .y(_T_2779),
        .a(_T_2778),
        .b(_WTEMP_435)
    );
    wire [63:0] _T_2780;
    wire [63:0] _WTEMP_436;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3280 (
        .y(_WTEMP_436),
        .in(_T_2575)
    );
    BITWISEOR #(.width(64)) bitwiseor_3281 (
        .y(_T_2780),
        .a(_T_2779),
        .b(_WTEMP_436)
    );
    wire [63:0] _T_2781;
    wire [63:0] _WTEMP_437;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3282 (
        .y(_WTEMP_437),
        .in(_T_2577)
    );
    BITWISEOR #(.width(64)) bitwiseor_3283 (
        .y(_T_2781),
        .a(_T_2780),
        .b(_WTEMP_437)
    );
    wire [63:0] _T_2782;
    wire [63:0] _WTEMP_438;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3284 (
        .y(_WTEMP_438),
        .in(_T_2579)
    );
    BITWISEOR #(.width(64)) bitwiseor_3285 (
        .y(_T_2782),
        .a(_T_2781),
        .b(_WTEMP_438)
    );
    wire [63:0] _T_2783;
    wire [63:0] _WTEMP_439;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3286 (
        .y(_WTEMP_439),
        .in(_T_2581)
    );
    BITWISEOR #(.width(64)) bitwiseor_3287 (
        .y(_T_2783),
        .a(_T_2782),
        .b(_WTEMP_439)
    );
    wire [63:0] _T_2784;
    wire [63:0] _WTEMP_440;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3288 (
        .y(_WTEMP_440),
        .in(_T_2583)
    );
    BITWISEOR #(.width(64)) bitwiseor_3289 (
        .y(_T_2784),
        .a(_T_2783),
        .b(_WTEMP_440)
    );
    wire [63:0] _T_2785;
    wire [63:0] _WTEMP_441;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3290 (
        .y(_WTEMP_441),
        .in(_T_2585)
    );
    BITWISEOR #(.width(64)) bitwiseor_3291 (
        .y(_T_2785),
        .a(_T_2784),
        .b(_WTEMP_441)
    );
    wire [63:0] _T_2786;
    wire [63:0] _WTEMP_442;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3292 (
        .y(_WTEMP_442),
        .in(_T_2587)
    );
    BITWISEOR #(.width(64)) bitwiseor_3293 (
        .y(_T_2786),
        .a(_T_2785),
        .b(_WTEMP_442)
    );
    wire [63:0] _T_2787;
    wire [63:0] _WTEMP_443;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3294 (
        .y(_WTEMP_443),
        .in(_T_2589)
    );
    BITWISEOR #(.width(64)) bitwiseor_3295 (
        .y(_T_2787),
        .a(_T_2786),
        .b(_WTEMP_443)
    );
    wire [63:0] _T_2788;
    wire [63:0] _WTEMP_444;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3296 (
        .y(_WTEMP_444),
        .in(_T_2591)
    );
    BITWISEOR #(.width(64)) bitwiseor_3297 (
        .y(_T_2788),
        .a(_T_2787),
        .b(_WTEMP_444)
    );
    wire [63:0] _T_2789;
    wire [63:0] _WTEMP_445;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3298 (
        .y(_WTEMP_445),
        .in(_T_2593)
    );
    BITWISEOR #(.width(64)) bitwiseor_3299 (
        .y(_T_2789),
        .a(_T_2788),
        .b(_WTEMP_445)
    );
    wire [63:0] _T_2790;
    wire [63:0] _WTEMP_446;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3300 (
        .y(_WTEMP_446),
        .in(_T_2595)
    );
    BITWISEOR #(.width(64)) bitwiseor_3301 (
        .y(_T_2790),
        .a(_T_2789),
        .b(_WTEMP_446)
    );
    wire [63:0] _T_2791;
    wire [63:0] _WTEMP_447;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3302 (
        .y(_WTEMP_447),
        .in(_T_2597)
    );
    BITWISEOR #(.width(64)) bitwiseor_3303 (
        .y(_T_2791),
        .a(_T_2790),
        .b(_WTEMP_447)
    );
    wire [63:0] _T_2792;
    wire [63:0] _WTEMP_448;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3304 (
        .y(_WTEMP_448),
        .in(_T_2599)
    );
    BITWISEOR #(.width(64)) bitwiseor_3305 (
        .y(_T_2792),
        .a(_T_2791),
        .b(_WTEMP_448)
    );
    wire [63:0] _T_2793;
    wire [63:0] _WTEMP_449;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3306 (
        .y(_WTEMP_449),
        .in(_T_2601)
    );
    BITWISEOR #(.width(64)) bitwiseor_3307 (
        .y(_T_2793),
        .a(_T_2792),
        .b(_WTEMP_449)
    );
    wire [63:0] _T_2794;
    wire [63:0] _WTEMP_450;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3308 (
        .y(_WTEMP_450),
        .in(_T_2603)
    );
    BITWISEOR #(.width(64)) bitwiseor_3309 (
        .y(_T_2794),
        .a(_T_2793),
        .b(_WTEMP_450)
    );
    wire [63:0] _T_2795;
    wire [63:0] _WTEMP_451;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3310 (
        .y(_WTEMP_451),
        .in(_T_2605)
    );
    BITWISEOR #(.width(64)) bitwiseor_3311 (
        .y(_T_2795),
        .a(_T_2794),
        .b(_WTEMP_451)
    );
    wire [63:0] _T_2796;
    wire [63:0] _WTEMP_452;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3312 (
        .y(_WTEMP_452),
        .in(_T_2607)
    );
    BITWISEOR #(.width(64)) bitwiseor_3313 (
        .y(_T_2796),
        .a(_T_2795),
        .b(_WTEMP_452)
    );
    wire [63:0] _T_2797;
    wire [63:0] _WTEMP_453;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3314 (
        .y(_WTEMP_453),
        .in(_T_2609)
    );
    BITWISEOR #(.width(64)) bitwiseor_3315 (
        .y(_T_2797),
        .a(_T_2796),
        .b(_WTEMP_453)
    );
    wire [63:0] _T_2798;
    wire [63:0] _WTEMP_454;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3316 (
        .y(_WTEMP_454),
        .in(_T_2611)
    );
    BITWISEOR #(.width(64)) bitwiseor_3317 (
        .y(_T_2798),
        .a(_T_2797),
        .b(_WTEMP_454)
    );
    wire [63:0] _T_2799;
    wire [63:0] _WTEMP_455;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3318 (
        .y(_WTEMP_455),
        .in(_T_2613)
    );
    BITWISEOR #(.width(64)) bitwiseor_3319 (
        .y(_T_2799),
        .a(_T_2798),
        .b(_WTEMP_455)
    );
    wire [63:0] _T_2800;
    wire [63:0] _WTEMP_456;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3320 (
        .y(_WTEMP_456),
        .in(_T_2615)
    );
    BITWISEOR #(.width(64)) bitwiseor_3321 (
        .y(_T_2800),
        .a(_T_2799),
        .b(_WTEMP_456)
    );
    wire [63:0] _T_2801;
    wire [63:0] _WTEMP_457;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3322 (
        .y(_WTEMP_457),
        .in(_T_2617)
    );
    BITWISEOR #(.width(64)) bitwiseor_3323 (
        .y(_T_2801),
        .a(_T_2800),
        .b(_WTEMP_457)
    );
    wire [63:0] _T_2802;
    wire [63:0] _WTEMP_458;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3324 (
        .y(_WTEMP_458),
        .in(_T_2619)
    );
    BITWISEOR #(.width(64)) bitwiseor_3325 (
        .y(_T_2802),
        .a(_T_2801),
        .b(_WTEMP_458)
    );
    wire [63:0] _T_2803;
    wire [63:0] _WTEMP_459;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3326 (
        .y(_WTEMP_459),
        .in(_T_2621)
    );
    BITWISEOR #(.width(64)) bitwiseor_3327 (
        .y(_T_2803),
        .a(_T_2802),
        .b(_WTEMP_459)
    );
    wire [63:0] _T_2804;
    wire [63:0] _WTEMP_460;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3328 (
        .y(_WTEMP_460),
        .in(_T_2623)
    );
    BITWISEOR #(.width(64)) bitwiseor_3329 (
        .y(_T_2804),
        .a(_T_2803),
        .b(_WTEMP_460)
    );
    wire [63:0] _T_2805;
    wire [63:0] _WTEMP_461;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3330 (
        .y(_WTEMP_461),
        .in(_T_2625)
    );
    BITWISEOR #(.width(64)) bitwiseor_3331 (
        .y(_T_2805),
        .a(_T_2804),
        .b(_WTEMP_461)
    );
    wire [63:0] _T_2806;
    wire [63:0] _WTEMP_462;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3332 (
        .y(_WTEMP_462),
        .in(_T_2627)
    );
    BITWISEOR #(.width(64)) bitwiseor_3333 (
        .y(_T_2806),
        .a(_T_2805),
        .b(_WTEMP_462)
    );
    wire [63:0] _T_2807;
    wire [63:0] _WTEMP_463;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3334 (
        .y(_WTEMP_463),
        .in(_T_2629)
    );
    BITWISEOR #(.width(64)) bitwiseor_3335 (
        .y(_T_2807),
        .a(_T_2806),
        .b(_WTEMP_463)
    );
    wire [63:0] _T_2808;
    wire [63:0] _WTEMP_464;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3336 (
        .y(_WTEMP_464),
        .in(_T_2631)
    );
    BITWISEOR #(.width(64)) bitwiseor_3337 (
        .y(_T_2808),
        .a(_T_2807),
        .b(_WTEMP_464)
    );
    wire [63:0] _T_2809;
    wire [63:0] _WTEMP_465;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3338 (
        .y(_WTEMP_465),
        .in(_T_2633)
    );
    BITWISEOR #(.width(64)) bitwiseor_3339 (
        .y(_T_2809),
        .a(_T_2808),
        .b(_WTEMP_465)
    );
    wire [63:0] _T_2810;
    wire [63:0] _WTEMP_466;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3340 (
        .y(_WTEMP_466),
        .in(_T_2635)
    );
    BITWISEOR #(.width(64)) bitwiseor_3341 (
        .y(_T_2810),
        .a(_T_2809),
        .b(_WTEMP_466)
    );
    wire [63:0] _T_2811;
    wire [63:0] _WTEMP_467;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3342 (
        .y(_WTEMP_467),
        .in(_T_2637)
    );
    BITWISEOR #(.width(64)) bitwiseor_3343 (
        .y(_T_2811),
        .a(_T_2810),
        .b(_WTEMP_467)
    );
    wire [63:0] _T_2812;
    wire [63:0] _WTEMP_468;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3344 (
        .y(_WTEMP_468),
        .in(_T_2639)
    );
    BITWISEOR #(.width(64)) bitwiseor_3345 (
        .y(_T_2812),
        .a(_T_2811),
        .b(_WTEMP_468)
    );
    wire [63:0] _T_2813;
    wire [63:0] _WTEMP_469;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3346 (
        .y(_WTEMP_469),
        .in(_T_2641)
    );
    BITWISEOR #(.width(64)) bitwiseor_3347 (
        .y(_T_2813),
        .a(_T_2812),
        .b(_WTEMP_469)
    );
    wire [63:0] _T_2814;
    wire [63:0] _WTEMP_470;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3348 (
        .y(_WTEMP_470),
        .in(_T_2643)
    );
    BITWISEOR #(.width(64)) bitwiseor_3349 (
        .y(_T_2814),
        .a(_T_2813),
        .b(_WTEMP_470)
    );
    wire [63:0] _T_2815;
    wire [63:0] _WTEMP_471;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3350 (
        .y(_WTEMP_471),
        .in(_T_2645)
    );
    BITWISEOR #(.width(64)) bitwiseor_3351 (
        .y(_T_2815),
        .a(_T_2814),
        .b(_WTEMP_471)
    );
    wire [63:0] _T_2816;
    wire [63:0] _WTEMP_472;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3352 (
        .y(_WTEMP_472),
        .in(_T_2647)
    );
    BITWISEOR #(.width(64)) bitwiseor_3353 (
        .y(_T_2816),
        .a(_T_2815),
        .b(_WTEMP_472)
    );
    wire [63:0] _T_2817;
    wire [63:0] _WTEMP_473;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3354 (
        .y(_WTEMP_473),
        .in(_T_2649)
    );
    BITWISEOR #(.width(64)) bitwiseor_3355 (
        .y(_T_2817),
        .a(_T_2816),
        .b(_WTEMP_473)
    );
    wire [63:0] _T_2818;
    wire [63:0] _WTEMP_474;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3356 (
        .y(_WTEMP_474),
        .in(_T_2651)
    );
    BITWISEOR #(.width(64)) bitwiseor_3357 (
        .y(_T_2818),
        .a(_T_2817),
        .b(_WTEMP_474)
    );
    wire [63:0] _T_2819;
    wire [63:0] _WTEMP_475;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3358 (
        .y(_WTEMP_475),
        .in(_T_2653)
    );
    BITWISEOR #(.width(64)) bitwiseor_3359 (
        .y(_T_2819),
        .a(_T_2818),
        .b(_WTEMP_475)
    );
    wire [63:0] _T_2820;
    wire [63:0] _WTEMP_476;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3360 (
        .y(_WTEMP_476),
        .in(_T_2655)
    );
    BITWISEOR #(.width(64)) bitwiseor_3361 (
        .y(_T_2820),
        .a(_T_2819),
        .b(_WTEMP_476)
    );
    wire [63:0] _T_2821;
    wire [63:0] _WTEMP_477;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3362 (
        .y(_WTEMP_477),
        .in(_T_2657)
    );
    BITWISEOR #(.width(64)) bitwiseor_3363 (
        .y(_T_2821),
        .a(_T_2820),
        .b(_WTEMP_477)
    );
    wire [63:0] _T_2822;
    wire [63:0] _WTEMP_478;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3364 (
        .y(_WTEMP_478),
        .in(_T_2659)
    );
    BITWISEOR #(.width(64)) bitwiseor_3365 (
        .y(_T_2822),
        .a(_T_2821),
        .b(_WTEMP_478)
    );
    wire [63:0] _T_2823;
    wire [63:0] _WTEMP_479;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3366 (
        .y(_WTEMP_479),
        .in(_T_2661)
    );
    BITWISEOR #(.width(64)) bitwiseor_3367 (
        .y(_T_2823),
        .a(_T_2822),
        .b(_WTEMP_479)
    );
    wire [63:0] _T_2824;
    wire [63:0] _WTEMP_480;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3368 (
        .y(_WTEMP_480),
        .in(_T_2663)
    );
    BITWISEOR #(.width(64)) bitwiseor_3369 (
        .y(_T_2824),
        .a(_T_2823),
        .b(_WTEMP_480)
    );
    wire [63:0] _T_2825;
    wire [63:0] _WTEMP_481;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3370 (
        .y(_WTEMP_481),
        .in(_T_2665)
    );
    BITWISEOR #(.width(64)) bitwiseor_3371 (
        .y(_T_2825),
        .a(_T_2824),
        .b(_WTEMP_481)
    );
    wire [63:0] _T_2826;
    wire [63:0] _WTEMP_482;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3372 (
        .y(_WTEMP_482),
        .in(_T_2667)
    );
    BITWISEOR #(.width(64)) bitwiseor_3373 (
        .y(_T_2826),
        .a(_T_2825),
        .b(_WTEMP_482)
    );
    wire [63:0] _T_2827;
    wire [63:0] _WTEMP_483;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3374 (
        .y(_WTEMP_483),
        .in(_T_2669)
    );
    BITWISEOR #(.width(64)) bitwiseor_3375 (
        .y(_T_2827),
        .a(_T_2826),
        .b(_WTEMP_483)
    );
    wire [63:0] _T_2828;
    wire [63:0] _WTEMP_484;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3376 (
        .y(_WTEMP_484),
        .in(_T_2671)
    );
    BITWISEOR #(.width(64)) bitwiseor_3377 (
        .y(_T_2828),
        .a(_T_2827),
        .b(_WTEMP_484)
    );
    wire [63:0] _T_2829;
    wire [63:0] _WTEMP_485;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3378 (
        .y(_WTEMP_485),
        .in(_T_2673)
    );
    BITWISEOR #(.width(64)) bitwiseor_3379 (
        .y(_T_2829),
        .a(_T_2828),
        .b(_WTEMP_485)
    );
    wire [63:0] _T_2830;
    wire [63:0] _WTEMP_486;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3380 (
        .y(_WTEMP_486),
        .in(_T_2675)
    );
    BITWISEOR #(.width(64)) bitwiseor_3381 (
        .y(_T_2830),
        .a(_T_2829),
        .b(_WTEMP_486)
    );
    wire [63:0] _T_2831;
    wire [63:0] _WTEMP_487;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3382 (
        .y(_WTEMP_487),
        .in(_T_2677)
    );
    BITWISEOR #(.width(64)) bitwiseor_3383 (
        .y(_T_2831),
        .a(_T_2830),
        .b(_WTEMP_487)
    );
    wire [63:0] _T_2832;
    wire [63:0] _WTEMP_488;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3384 (
        .y(_WTEMP_488),
        .in(_T_2679)
    );
    BITWISEOR #(.width(64)) bitwiseor_3385 (
        .y(_T_2832),
        .a(_T_2831),
        .b(_WTEMP_488)
    );
    wire [63:0] _T_2833;
    wire [63:0] _WTEMP_489;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3386 (
        .y(_WTEMP_489),
        .in(_T_2681)
    );
    BITWISEOR #(.width(64)) bitwiseor_3387 (
        .y(_T_2833),
        .a(_T_2832),
        .b(_WTEMP_489)
    );
    wire [63:0] _T_2834;
    wire [63:0] _WTEMP_490;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3388 (
        .y(_WTEMP_490),
        .in(_T_2683)
    );
    BITWISEOR #(.width(64)) bitwiseor_3389 (
        .y(_T_2834),
        .a(_T_2833),
        .b(_WTEMP_490)
    );
    wire [63:0] _T_2835;
    wire [63:0] _WTEMP_491;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3390 (
        .y(_WTEMP_491),
        .in(_T_2685)
    );
    BITWISEOR #(.width(64)) bitwiseor_3391 (
        .y(_T_2835),
        .a(_T_2834),
        .b(_WTEMP_491)
    );
    wire [63:0] _T_2836;
    wire [63:0] _WTEMP_492;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3392 (
        .y(_WTEMP_492),
        .in(_T_2687)
    );
    BITWISEOR #(.width(64)) bitwiseor_3393 (
        .y(_T_2836),
        .a(_T_2835),
        .b(_WTEMP_492)
    );
    wire [63:0] _T_2837;
    wire [63:0] _WTEMP_493;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3394 (
        .y(_WTEMP_493),
        .in(_T_2689)
    );
    BITWISEOR #(.width(64)) bitwiseor_3395 (
        .y(_T_2837),
        .a(_T_2836),
        .b(_WTEMP_493)
    );
    wire [63:0] _T_2838;
    wire [63:0] _WTEMP_494;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3396 (
        .y(_WTEMP_494),
        .in(_T_2691)
    );
    BITWISEOR #(.width(64)) bitwiseor_3397 (
        .y(_T_2838),
        .a(_T_2837),
        .b(_WTEMP_494)
    );
    wire [63:0] _T_2839;
    wire [63:0] _WTEMP_495;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3398 (
        .y(_WTEMP_495),
        .in(_T_2693)
    );
    BITWISEOR #(.width(64)) bitwiseor_3399 (
        .y(_T_2839),
        .a(_T_2838),
        .b(_WTEMP_495)
    );
    wire [63:0] _T_2840;
    wire [63:0] _WTEMP_496;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3400 (
        .y(_WTEMP_496),
        .in(_T_2695)
    );
    BITWISEOR #(.width(64)) bitwiseor_3401 (
        .y(_T_2840),
        .a(_T_2839),
        .b(_WTEMP_496)
    );
    wire [63:0] _T_2841;
    wire [63:0] _WTEMP_497;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3402 (
        .y(_WTEMP_497),
        .in(_T_2697)
    );
    BITWISEOR #(.width(64)) bitwiseor_3403 (
        .y(_T_2841),
        .a(_T_2840),
        .b(_WTEMP_497)
    );
    wire [63:0] _T_2842;
    wire [63:0] _WTEMP_498;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3404 (
        .y(_WTEMP_498),
        .in(_T_2699)
    );
    BITWISEOR #(.width(64)) bitwiseor_3405 (
        .y(_T_2842),
        .a(_T_2841),
        .b(_WTEMP_498)
    );
    wire [63:0] _T_2843;
    wire [63:0] _WTEMP_499;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3406 (
        .y(_WTEMP_499),
        .in(_T_2701)
    );
    BITWISEOR #(.width(64)) bitwiseor_3407 (
        .y(_T_2843),
        .a(_T_2842),
        .b(_WTEMP_499)
    );
    wire [63:0] _T_2844;
    wire [63:0] _WTEMP_500;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3408 (
        .y(_WTEMP_500),
        .in(_T_2703)
    );
    BITWISEOR #(.width(64)) bitwiseor_3409 (
        .y(_T_2844),
        .a(_T_2843),
        .b(_WTEMP_500)
    );
    wire [63:0] _T_2845;
    wire [63:0] _WTEMP_501;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3410 (
        .y(_WTEMP_501),
        .in(_T_2705)
    );
    BITWISEOR #(.width(64)) bitwiseor_3411 (
        .y(_T_2845),
        .a(_T_2844),
        .b(_WTEMP_501)
    );
    wire [63:0] _T_2846;
    wire [63:0] _WTEMP_502;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3412 (
        .y(_WTEMP_502),
        .in(_T_2707)
    );
    BITWISEOR #(.width(64)) bitwiseor_3413 (
        .y(_T_2846),
        .a(_T_2845),
        .b(_WTEMP_502)
    );
    wire [63:0] _T_2847;
    BITWISEOR #(.width(64)) bitwiseor_3414 (
        .y(_T_2847),
        .a(_T_2846),
        .b(_T_2709)
    );
    wire [63:0] _T_2848;
    BITWISEOR #(.width(64)) bitwiseor_3415 (
        .y(_T_2848),
        .a(_T_2847),
        .b(_T_2711)
    );
    wire [63:0] _T_2849;
    BITWISEOR #(.width(64)) bitwiseor_3416 (
        .y(_T_2849),
        .a(_T_2848),
        .b(_T_2713)
    );
    wire [63:0] _T_2850;
    BITWISEOR #(.width(64)) bitwiseor_3417 (
        .y(_T_2850),
        .a(_T_2849),
        .b(_T_2715)
    );
    wire [63:0] _T_2851;
    BITWISEOR #(.width(64)) bitwiseor_3418 (
        .y(_T_2851),
        .a(_T_2850),
        .b(_T_2717)
    );
    wire [63:0] _T_2852;
    BITWISEOR #(.width(64)) bitwiseor_3419 (
        .y(_T_2852),
        .a(_T_2851),
        .b(_T_2719)
    );
    wire [63:0] _T_2853;
    BITWISEOR #(.width(64)) bitwiseor_3420 (
        .y(_T_2853),
        .a(_T_2852),
        .b(_T_2721)
    );
    wire [63:0] _T_2854;
    BITWISEOR #(.width(64)) bitwiseor_3421 (
        .y(_T_2854),
        .a(_T_2853),
        .b(_T_2723)
    );
    wire [63:0] _T_2855;
    BITWISEOR #(.width(64)) bitwiseor_3422 (
        .y(_T_2855),
        .a(_T_2854),
        .b(_T_2725)
    );
    wire [63:0] _T_2856;
    wire [63:0] _WTEMP_503;
    PAD_UNSIGNED #(.width(32), .n(64)) u_pad_3423 (
        .y(_WTEMP_503),
        .in(_T_2727)
    );
    BITWISEOR #(.width(64)) bitwiseor_3424 (
        .y(_T_2856),
        .a(_T_2855),
        .b(_WTEMP_503)
    );
    wire [63:0] _T_2857;
    wire [63:0] _WTEMP_504;
    PAD_UNSIGNED #(.width(32), .n(64)) u_pad_3425 (
        .y(_WTEMP_504),
        .in(_T_2729)
    );
    BITWISEOR #(.width(64)) bitwiseor_3426 (
        .y(_T_2857),
        .a(_T_2856),
        .b(_WTEMP_504)
    );
    wire [63:0] _T_2858;
    BITWISEOR #(.width(64)) bitwiseor_3427 (
        .y(_T_2858),
        .a(_T_2857),
        .b(_T_2731)
    );
    wire [63:0] _T_2859;
    BITWISEOR #(.width(64)) bitwiseor_3428 (
        .y(_T_2859),
        .a(_T_2858),
        .b(_T_2733)
    );
    wire [63:0] _T_2861;
    wire [4:0] _T_2862;
    BITWISEOR #(.width(5)) bitwiseor_3429 (
        .y(_T_2862),
        .a(_reg_fflags__q),
        .b(io_fcsr_flags_bits)
    );
    wire _T_2866;
    EQ_UNSIGNED #(.width(3)) u_eq_3430 (
        .y(_T_2866),
        .a(io_rw_cmd),
        .b(3'h2)
    );
    wire _T_2867;
    EQ_UNSIGNED #(.width(3)) u_eq_3431 (
        .y(_T_2867),
        .a(io_rw_cmd),
        .b(3'h3)
    );
    wire _T_2868;
    EQ_UNSIGNED #(.width(3)) u_eq_3432 (
        .y(_T_2868),
        .a(io_rw_cmd),
        .b(3'h1)
    );
    wire _T_2869;
    BITWISEOR #(.width(1)) bitwiseor_3433 (
        .y(_T_2869),
        .a(_T_2866),
        .b(_T_2867)
    );
    wire _T_2870;
    BITWISEOR #(.width(1)) bitwiseor_3434 (
        .y(_T_2870),
        .a(_T_2869),
        .b(_T_2868)
    );
    wire _T_2929_debug;
    wire [31:0] _T_2929_isa;
    wire [1:0] _T_2929_prv;
    wire _T_2929_sd;
    wire [26:0] _T_2929_zero2;
    wire [1:0] _T_2929_sxl;
    wire [1:0] _T_2929_uxl;
    wire _T_2929_sd_rv32;
    wire [7:0] _T_2929_zero1;
    wire _T_2929_tsr;
    wire _T_2929_tw;
    wire _T_2929_tvm;
    wire _T_2929_mxr;
    wire _T_2929_pum;
    wire _T_2929_mprv;
    wire [1:0] _T_2929_xs;
    wire [1:0] _T_2929_fs;
    wire [1:0] _T_2929_mpp;
    wire [1:0] _T_2929_hpp;
    wire _T_2929_spp;
    wire _T_2929_mpie;
    wire _T_2929_hpie;
    wire _T_2929_spie;
    wire _T_2929_upie;
    wire _T_2929_mie;
    wire _T_2929_hie;
    wire _T_2929_sie;
    wire _T_2929_uie;
    wire [98:0] _T_2959;
    wire _T_2960;
    BITS #(.width(99), .high(0), .low(0)) bits_3435 (
        .y(_T_2960),
        .in(_T_2959)
    );
    wire _T_2961;
    BITS #(.width(99), .high(1), .low(1)) bits_3436 (
        .y(_T_2961),
        .in(_T_2959)
    );
    wire _T_2962;
    BITS #(.width(99), .high(2), .low(2)) bits_3437 (
        .y(_T_2962),
        .in(_T_2959)
    );
    wire _T_2963;
    BITS #(.width(99), .high(3), .low(3)) bits_3438 (
        .y(_T_2963),
        .in(_T_2959)
    );
    wire _T_2964;
    BITS #(.width(99), .high(4), .low(4)) bits_3439 (
        .y(_T_2964),
        .in(_T_2959)
    );
    wire _T_2965;
    BITS #(.width(99), .high(5), .low(5)) bits_3440 (
        .y(_T_2965),
        .in(_T_2959)
    );
    wire _T_2966;
    BITS #(.width(99), .high(6), .low(6)) bits_3441 (
        .y(_T_2966),
        .in(_T_2959)
    );
    wire _T_2967;
    BITS #(.width(99), .high(7), .low(7)) bits_3442 (
        .y(_T_2967),
        .in(_T_2959)
    );
    wire _T_2968;
    BITS #(.width(99), .high(8), .low(8)) bits_3443 (
        .y(_T_2968),
        .in(_T_2959)
    );
    wire [1:0] _T_2969;
    BITS #(.width(99), .high(10), .low(9)) bits_3444 (
        .y(_T_2969),
        .in(_T_2959)
    );
    wire [1:0] _T_2970;
    BITS #(.width(99), .high(12), .low(11)) bits_3445 (
        .y(_T_2970),
        .in(_T_2959)
    );
    wire [1:0] _T_2971;
    BITS #(.width(99), .high(14), .low(13)) bits_3446 (
        .y(_T_2971),
        .in(_T_2959)
    );
    wire [1:0] _T_2972;
    BITS #(.width(99), .high(16), .low(15)) bits_3447 (
        .y(_T_2972),
        .in(_T_2959)
    );
    wire _T_2973;
    BITS #(.width(99), .high(17), .low(17)) bits_3448 (
        .y(_T_2973),
        .in(_T_2959)
    );
    wire _T_2974;
    BITS #(.width(99), .high(18), .low(18)) bits_3449 (
        .y(_T_2974),
        .in(_T_2959)
    );
    wire _T_2975;
    BITS #(.width(99), .high(19), .low(19)) bits_3450 (
        .y(_T_2975),
        .in(_T_2959)
    );
    wire _T_2976;
    BITS #(.width(99), .high(20), .low(20)) bits_3451 (
        .y(_T_2976),
        .in(_T_2959)
    );
    wire _T_2977;
    BITS #(.width(99), .high(21), .low(21)) bits_3452 (
        .y(_T_2977),
        .in(_T_2959)
    );
    wire _T_2978;
    BITS #(.width(99), .high(22), .low(22)) bits_3453 (
        .y(_T_2978),
        .in(_T_2959)
    );
    wire [7:0] _T_2979;
    BITS #(.width(99), .high(30), .low(23)) bits_3454 (
        .y(_T_2979),
        .in(_T_2959)
    );
    wire _T_2980;
    BITS #(.width(99), .high(31), .low(31)) bits_3455 (
        .y(_T_2980),
        .in(_T_2959)
    );
    wire [1:0] _T_2981;
    BITS #(.width(99), .high(33), .low(32)) bits_3456 (
        .y(_T_2981),
        .in(_T_2959)
    );
    wire [1:0] _T_2982;
    BITS #(.width(99), .high(35), .low(34)) bits_3457 (
        .y(_T_2982),
        .in(_T_2959)
    );
    wire [26:0] _T_2983;
    BITS #(.width(99), .high(62), .low(36)) bits_3458 (
        .y(_T_2983),
        .in(_T_2959)
    );
    wire _T_2984;
    BITS #(.width(99), .high(63), .low(63)) bits_3459 (
        .y(_T_2984),
        .in(_T_2959)
    );
    wire [1:0] _T_2985;
    BITS #(.width(99), .high(65), .low(64)) bits_3460 (
        .y(_T_2985),
        .in(_T_2959)
    );
    wire [31:0] _T_2986;
    BITS #(.width(99), .high(97), .low(66)) bits_3461 (
        .y(_T_2986),
        .in(_T_2959)
    );
    wire _T_2987;
    BITS #(.width(99), .high(98), .low(98)) bits_3462 (
        .y(_T_2987),
        .in(_T_2959)
    );
    wire _T_2989;
    wire [1:0] _WTEMP_505;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_3463 (
        .y(_WTEMP_505),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(2)) u_neq_3464 (
        .y(_T_2989),
        .a(_T_2929_fs),
        .b(_WTEMP_505)
    );
    wire _T_2990;
    BITS #(.width(1), .high(0), .low(0)) bits_3465 (
        .y(_T_2990),
        .in(_T_2989)
    );
    wire [1:0] _T_2993;
    MUX_UNSIGNED #(.width(2)) u_mux_3466 (
        .y(_T_2993),
        .sel(_T_2990),
        .a(2'h3),
        .b(2'h0)
    );
    wire _node_66;
    MUX_UNSIGNED #(.width(1)) u_mux_3467 (
        .y(_node_66),
        .sel(insn_ret),
        .a(_node_54),
        .b(_node_55)
    );
    wire _node_67;
    MUX_UNSIGNED #(.width(1)) u_mux_3468 (
        .y(_node_67),
        .sel(insn_ret),
        .a(_node_56),
        .b(_node_57)
    );
    wire [1:0] _node_68;
    MUX_UNSIGNED #(.width(2)) u_mux_3469 (
        .y(_node_68),
        .sel(insn_ret),
        .a(_node_58),
        .b(_node_59)
    );
    wire _node_69;
    MUX_UNSIGNED #(.width(1)) u_mux_3470 (
        .y(_node_69),
        .sel(insn_ret),
        .a(_node_60),
        .b(_node_61)
    );
    wire _node_70;
    MUX_UNSIGNED #(.width(1)) u_mux_3471 (
        .y(_node_70),
        .sel(insn_ret),
        .a(_node_62),
        .b(_node_63)
    );
    wire [1:0] _node_71;
    MUX_UNSIGNED #(.width(2)) u_mux_3472 (
        .y(_node_71),
        .sel(insn_ret),
        .a(_node_64),
        .b(_node_65)
    );
    wire _T_2995;
    BITS #(.width(64), .high(5), .low(5)) bits_3473 (
        .y(_T_2995),
        .in(wdata)
    );
    wire [63:0] _T_2996;
    BITWISENOT #(.width(64)) bitwisenot_3474 (
        .y(_T_2996),
        .in(wdata)
    );
    wire _T_2998;
    EQ_UNSIGNED #(.width(1)) u_eq_3475 (
        .y(_T_2998),
        .a(_T_2995),
        .b(1'h0)
    );
    wire [3:0] _T_2999;
    SHL_UNSIGNED #(.width(1), .n(3)) u_shl_3476 (
        .y(_T_2999),
        .in(_T_2998)
    );
    wire [63:0] _T_3000;
    wire [63:0] _WTEMP_506;
    PAD_UNSIGNED #(.width(4), .n(64)) u_pad_3477 (
        .y(_WTEMP_506),
        .in(_T_2999)
    );
    BITWISEOR #(.width(64)) bitwiseor_3478 (
        .y(_T_3000),
        .a(_T_2996),
        .b(_WTEMP_506)
    );
    wire [63:0] _T_3001;
    BITWISENOT #(.width(64)) bitwisenot_3479 (
        .y(_T_3001),
        .in(_T_3000)
    );
    wire [63:0] _T_3002;
    wire [63:0] _WTEMP_507;
    PAD_UNSIGNED #(.width(13), .n(64)) u_pad_3480 (
        .y(_WTEMP_507),
        .in(13'h102D)
    );
    BITWISEAND #(.width(64)) bitwiseand_3481 (
        .y(_T_3002),
        .a(_T_3001),
        .b(_WTEMP_507)
    );
    wire [12:0] _T_3003;
    assign _T_3003 = 13'hFD2;
    wire [63:0] _T_3004;
    wire [63:0] _WTEMP_508;
    PAD_UNSIGNED #(.width(13), .n(64)) u_pad_3482 (
        .y(_WTEMP_508),
        .in(_T_3003)
    );
    BITWISEAND #(.width(64)) bitwiseand_3483 (
        .y(_T_3004),
        .a(_reg_misa__q),
        .b(_WTEMP_508)
    );
    wire [63:0] _T_3005;
    BITWISEOR #(.width(64)) bitwiseor_3484 (
        .y(_T_3005),
        .a(_T_3002),
        .b(_T_3004)
    );
    wire _T_3034_rocc;
    wire _T_3034_meip;
    wire _T_3034_heip;
    wire _T_3034_seip;
    wire _T_3034_ueip;
    wire _T_3034_mtip;
    wire _T_3034_htip;
    wire _T_3034_stip;
    wire _T_3034_utip;
    wire _T_3034_msip;
    wire _T_3034_hsip;
    wire _T_3034_ssip;
    wire _T_3034_usip;
    wire [12:0] _T_3049;
    wire _T_3050;
    BITS #(.width(13), .high(0), .low(0)) bits_3485 (
        .y(_T_3050),
        .in(_T_3049)
    );
    wire _T_3051;
    BITS #(.width(13), .high(1), .low(1)) bits_3486 (
        .y(_T_3051),
        .in(_T_3049)
    );
    wire _T_3052;
    BITS #(.width(13), .high(2), .low(2)) bits_3487 (
        .y(_T_3052),
        .in(_T_3049)
    );
    wire _T_3053;
    BITS #(.width(13), .high(3), .low(3)) bits_3488 (
        .y(_T_3053),
        .in(_T_3049)
    );
    wire _T_3054;
    BITS #(.width(13), .high(4), .low(4)) bits_3489 (
        .y(_T_3054),
        .in(_T_3049)
    );
    wire _T_3055;
    BITS #(.width(13), .high(5), .low(5)) bits_3490 (
        .y(_T_3055),
        .in(_T_3049)
    );
    wire _T_3056;
    BITS #(.width(13), .high(6), .low(6)) bits_3491 (
        .y(_T_3056),
        .in(_T_3049)
    );
    wire _T_3057;
    BITS #(.width(13), .high(7), .low(7)) bits_3492 (
        .y(_T_3057),
        .in(_T_3049)
    );
    wire _T_3058;
    BITS #(.width(13), .high(8), .low(8)) bits_3493 (
        .y(_T_3058),
        .in(_T_3049)
    );
    wire _T_3059;
    BITS #(.width(13), .high(9), .low(9)) bits_3494 (
        .y(_T_3059),
        .in(_T_3049)
    );
    wire _T_3060;
    BITS #(.width(13), .high(10), .low(10)) bits_3495 (
        .y(_T_3060),
        .in(_T_3049)
    );
    wire _T_3061;
    BITS #(.width(13), .high(11), .low(11)) bits_3496 (
        .y(_T_3061),
        .in(_T_3049)
    );
    wire _T_3062;
    BITS #(.width(13), .high(12), .low(12)) bits_3497 (
        .y(_T_3062),
        .in(_T_3049)
    );
    wire [63:0] _T_3063;
    wire [63:0] _WTEMP_509;
    PAD_UNSIGNED #(.width(13), .n(64)) u_pad_3498 (
        .y(_WTEMP_509),
        .in(supported_interrupts)
    );
    BITWISEAND #(.width(64)) bitwiseand_3499 (
        .y(_T_3063),
        .a(wdata),
        .b(_WTEMP_509)
    );
    wire [63:0] _T_3064;
    BITWISENOT #(.width(64)) bitwisenot_3500 (
        .y(_T_3064),
        .in(wdata)
    );
    wire _T_3065;
    BITS #(.width(64), .high(2), .low(2)) bits_3501 (
        .y(_T_3065),
        .in(_reg_misa__q)
    );
    wire _T_3067;
    EQ_UNSIGNED #(.width(1)) u_eq_3502 (
        .y(_T_3067),
        .a(_T_3065),
        .b(1'h0)
    );
    wire [1:0] _T_3069;
    CAT #(.width_a(1), .width_b(1)) cat_3503 (
        .y(_T_3069),
        .a(_T_3067),
        .b(1'h1)
    );
    wire [63:0] _T_3070;
    wire [63:0] _WTEMP_510;
    PAD_UNSIGNED #(.width(2), .n(64)) u_pad_3504 (
        .y(_WTEMP_510),
        .in(_T_3069)
    );
    BITWISEOR #(.width(64)) bitwiseor_3505 (
        .y(_T_3070),
        .a(_T_3064),
        .b(_WTEMP_510)
    );
    wire [63:0] _T_3071;
    BITWISENOT #(.width(64)) bitwisenot_3506 (
        .y(_T_3071),
        .in(_T_3070)
    );
    wire [39:0] _node_72;
    MUX_UNSIGNED #(.width(40)) u_mux_3507 (
        .y(_node_72),
        .sel(exception),
        .a(_node_20),
        .b(_reg_mepc__q)
    );
    wire [61:0] _T_3072;
    SHR_UNSIGNED #(.width(64), .n(2)) u_shr_3508 (
        .y(_T_3072),
        .in(wdata)
    );
    wire [63:0] _T_3073;
    SHL_UNSIGNED #(.width(62), .n(2)) u_shl_3509 (
        .y(_T_3073),
        .in(_T_3072)
    );
    wire [63:0] _T_3075;
    BITWISEAND #(.width(64)) bitwiseand_3510 (
        .y(_T_3075),
        .a(wdata),
        .b(64'h800000000000001F)
    );
    wire [63:0] _node_73;
    MUX_UNSIGNED #(.width(64)) u_mux_3511 (
        .y(_node_73),
        .sel(exception),
        .a(_node_19),
        .b(_reg_mcause__q)
    );
    wire [39:0] _T_3076;
    BITS #(.width(64), .high(39), .low(0)) bits_3512 (
        .y(_T_3076),
        .in(wdata)
    );
    wire [39:0] _node_74;
    MUX_UNSIGNED #(.width(40)) u_mux_3513 (
        .y(_node_74),
        .sel(exception),
        .a(_node_18),
        .b(_reg_mbadaddr__q)
    );
    wire [63:0] _T_3077;
    BITS #(.width(64), .high(63), .low(0)) bits_3514 (
        .y(_T_3077),
        .in(wdata)
    );
    wire [57:0] _T_3078;
    SHR_UNSIGNED #(.width(64), .n(6)) u_shr_3515 (
        .y(_T_3078),
        .in(_T_3077)
    );
    wire [57:0] _node_75;
    MUX_UNSIGNED #(.width(58)) u_mux_3516 (
        .y(_node_75),
        .sel(_T_946),
        .a(_T_949),
        .b(__T_945__q)
    );
    wire [63:0] _T_3079;
    BITS #(.width(64), .high(63), .low(0)) bits_3517 (
        .y(_T_3079),
        .in(wdata)
    );
    wire [57:0] _T_3080;
    SHR_UNSIGNED #(.width(64), .n(6)) u_shr_3518 (
        .y(_T_3080),
        .in(_T_3079)
    );
    wire [57:0] _node_76;
    MUX_UNSIGNED #(.width(58)) u_mux_3519 (
        .y(_node_76),
        .sel(_T_935),
        .a(_T_938),
        .b(__T_934__q)
    );
    wire [4:0] _node_77;
    MUX_UNSIGNED #(.width(5)) u_mux_3520 (
        .y(_node_77),
        .sel(io_fcsr_flags_valid),
        .a(_T_2862),
        .b(_reg_fflags__q)
    );
    wire [58:0] _T_3081;
    SHR_UNSIGNED #(.width(64), .n(5)) u_shr_3521 (
        .y(_T_3081),
        .in(wdata)
    );
    wire [63:0] _node_78;
    wire [63:0] _WTEMP_511;
    PAD_UNSIGNED #(.width(5), .n(64)) u_pad_3522 (
        .y(_WTEMP_511),
        .in(_node_77)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_3523 (
        .y(_node_78),
        .sel(_T_1513),
        .a(wdata),
        .b(_WTEMP_511)
    );
    wire [63:0] _node_79;
    wire [63:0] _WTEMP_512;
    PAD_UNSIGNED #(.width(3), .n(64)) u_pad_3524 (
        .y(_WTEMP_512),
        .in(_reg_frm__q)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_3525 (
        .y(_node_79),
        .sel(_T_1515),
        .a(wdata),
        .b(_WTEMP_512)
    );
    wire [1:0] _T_3118_xdebugver;
    wire _T_3118_ndreset;
    wire _T_3118_fullreset;
    wire [11:0] _T_3118_zero3;
    wire _T_3118_ebreakm;
    wire _T_3118_ebreakh;
    wire _T_3118_ebreaks;
    wire _T_3118_ebreaku;
    wire _T_3118_zero2;
    wire _T_3118_stopcycle;
    wire _T_3118_stoptime;
    wire [2:0] _T_3118_cause;
    wire _T_3118_debugint;
    wire _T_3118_zero1;
    wire _T_3118_halt;
    wire _T_3118_step;
    wire [1:0] _T_3118_prv;
    wire [31:0] _T_3137;
    wire [1:0] _T_3138;
    BITS #(.width(32), .high(1), .low(0)) bits_3526 (
        .y(_T_3138),
        .in(_T_3137)
    );
    wire _T_3139;
    BITS #(.width(32), .high(2), .low(2)) bits_3527 (
        .y(_T_3139),
        .in(_T_3137)
    );
    wire _T_3140;
    BITS #(.width(32), .high(3), .low(3)) bits_3528 (
        .y(_T_3140),
        .in(_T_3137)
    );
    wire _T_3141;
    BITS #(.width(32), .high(4), .low(4)) bits_3529 (
        .y(_T_3141),
        .in(_T_3137)
    );
    wire _T_3142;
    BITS #(.width(32), .high(5), .low(5)) bits_3530 (
        .y(_T_3142),
        .in(_T_3137)
    );
    wire [2:0] _T_3143;
    BITS #(.width(32), .high(8), .low(6)) bits_3531 (
        .y(_T_3143),
        .in(_T_3137)
    );
    wire _T_3144;
    BITS #(.width(32), .high(9), .low(9)) bits_3532 (
        .y(_T_3144),
        .in(_T_3137)
    );
    wire _T_3145;
    BITS #(.width(32), .high(10), .low(10)) bits_3533 (
        .y(_T_3145),
        .in(_T_3137)
    );
    wire _T_3146;
    BITS #(.width(32), .high(11), .low(11)) bits_3534 (
        .y(_T_3146),
        .in(_T_3137)
    );
    wire _T_3147;
    BITS #(.width(32), .high(12), .low(12)) bits_3535 (
        .y(_T_3147),
        .in(_T_3137)
    );
    wire _T_3148;
    BITS #(.width(32), .high(13), .low(13)) bits_3536 (
        .y(_T_3148),
        .in(_T_3137)
    );
    wire _T_3149;
    BITS #(.width(32), .high(14), .low(14)) bits_3537 (
        .y(_T_3149),
        .in(_T_3137)
    );
    wire _T_3150;
    BITS #(.width(32), .high(15), .low(15)) bits_3538 (
        .y(_T_3150),
        .in(_T_3137)
    );
    wire [11:0] _T_3151;
    BITS #(.width(32), .high(27), .low(16)) bits_3539 (
        .y(_T_3151),
        .in(_T_3137)
    );
    wire _T_3152;
    BITS #(.width(32), .high(28), .low(28)) bits_3540 (
        .y(_T_3152),
        .in(_T_3137)
    );
    wire _T_3153;
    BITS #(.width(32), .high(29), .low(29)) bits_3541 (
        .y(_T_3153),
        .in(_T_3137)
    );
    wire [1:0] _T_3154;
    BITS #(.width(32), .high(31), .low(30)) bits_3542 (
        .y(_T_3154),
        .in(_T_3137)
    );
    wire [1:0] _node_80;
    MUX_UNSIGNED #(.width(2)) u_mux_3543 (
        .y(_node_80),
        .sel(exception),
        .a(_node_15),
        .b(_reg_dcsr_prv__q)
    );
    wire [63:0] _T_3155;
    BITWISENOT #(.width(64)) bitwisenot_3544 (
        .y(_T_3155),
        .in(wdata)
    );
    wire [63:0] _T_3157;
    wire [63:0] _WTEMP_513;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_3545 (
        .y(_WTEMP_513),
        .in(1'h1)
    );
    BITWISEOR #(.width(64)) bitwiseor_3546 (
        .y(_T_3157),
        .a(_T_3155),
        .b(_WTEMP_513)
    );
    wire [63:0] _T_3158;
    BITWISENOT #(.width(64)) bitwisenot_3547 (
        .y(_T_3158),
        .in(_T_3157)
    );
    wire [39:0] _node_81;
    MUX_UNSIGNED #(.width(40)) u_mux_3548 (
        .y(_node_81),
        .sel(exception),
        .a(_node_17),
        .b(_reg_dpc__q)
    );
    wire _T_3217_debug;
    wire [31:0] _T_3217_isa;
    wire [1:0] _T_3217_prv;
    wire _T_3217_sd;
    wire [26:0] _T_3217_zero2;
    wire [1:0] _T_3217_sxl;
    wire [1:0] _T_3217_uxl;
    wire _T_3217_sd_rv32;
    wire [7:0] _T_3217_zero1;
    wire _T_3217_tsr;
    wire _T_3217_tw;
    wire _T_3217_tvm;
    wire _T_3217_mxr;
    wire _T_3217_pum;
    wire _T_3217_mprv;
    wire [1:0] _T_3217_xs;
    wire [1:0] _T_3217_fs;
    wire [1:0] _T_3217_mpp;
    wire [1:0] _T_3217_hpp;
    wire _T_3217_spp;
    wire _T_3217_mpie;
    wire _T_3217_hpie;
    wire _T_3217_spie;
    wire _T_3217_upie;
    wire _T_3217_mie;
    wire _T_3217_hie;
    wire _T_3217_sie;
    wire _T_3217_uie;
    wire [98:0] _T_3247;
    wire _T_3248;
    BITS #(.width(99), .high(0), .low(0)) bits_3549 (
        .y(_T_3248),
        .in(_T_3247)
    );
    wire _T_3249;
    BITS #(.width(99), .high(1), .low(1)) bits_3550 (
        .y(_T_3249),
        .in(_T_3247)
    );
    wire _T_3250;
    BITS #(.width(99), .high(2), .low(2)) bits_3551 (
        .y(_T_3250),
        .in(_T_3247)
    );
    wire _T_3251;
    BITS #(.width(99), .high(3), .low(3)) bits_3552 (
        .y(_T_3251),
        .in(_T_3247)
    );
    wire _T_3252;
    BITS #(.width(99), .high(4), .low(4)) bits_3553 (
        .y(_T_3252),
        .in(_T_3247)
    );
    wire _T_3253;
    BITS #(.width(99), .high(5), .low(5)) bits_3554 (
        .y(_T_3253),
        .in(_T_3247)
    );
    wire _T_3254;
    BITS #(.width(99), .high(6), .low(6)) bits_3555 (
        .y(_T_3254),
        .in(_T_3247)
    );
    wire _T_3255;
    BITS #(.width(99), .high(7), .low(7)) bits_3556 (
        .y(_T_3255),
        .in(_T_3247)
    );
    wire _T_3256;
    BITS #(.width(99), .high(8), .low(8)) bits_3557 (
        .y(_T_3256),
        .in(_T_3247)
    );
    wire [1:0] _T_3257;
    BITS #(.width(99), .high(10), .low(9)) bits_3558 (
        .y(_T_3257),
        .in(_T_3247)
    );
    wire [1:0] _T_3258;
    BITS #(.width(99), .high(12), .low(11)) bits_3559 (
        .y(_T_3258),
        .in(_T_3247)
    );
    wire [1:0] _T_3259;
    BITS #(.width(99), .high(14), .low(13)) bits_3560 (
        .y(_T_3259),
        .in(_T_3247)
    );
    wire [1:0] _T_3260;
    BITS #(.width(99), .high(16), .low(15)) bits_3561 (
        .y(_T_3260),
        .in(_T_3247)
    );
    wire _T_3261;
    BITS #(.width(99), .high(17), .low(17)) bits_3562 (
        .y(_T_3261),
        .in(_T_3247)
    );
    wire _T_3262;
    BITS #(.width(99), .high(18), .low(18)) bits_3563 (
        .y(_T_3262),
        .in(_T_3247)
    );
    wire _T_3263;
    BITS #(.width(99), .high(19), .low(19)) bits_3564 (
        .y(_T_3263),
        .in(_T_3247)
    );
    wire _T_3264;
    BITS #(.width(99), .high(20), .low(20)) bits_3565 (
        .y(_T_3264),
        .in(_T_3247)
    );
    wire _T_3265;
    BITS #(.width(99), .high(21), .low(21)) bits_3566 (
        .y(_T_3265),
        .in(_T_3247)
    );
    wire _T_3266;
    BITS #(.width(99), .high(22), .low(22)) bits_3567 (
        .y(_T_3266),
        .in(_T_3247)
    );
    wire [7:0] _T_3267;
    BITS #(.width(99), .high(30), .low(23)) bits_3568 (
        .y(_T_3267),
        .in(_T_3247)
    );
    wire _T_3268;
    BITS #(.width(99), .high(31), .low(31)) bits_3569 (
        .y(_T_3268),
        .in(_T_3247)
    );
    wire [1:0] _T_3269;
    BITS #(.width(99), .high(33), .low(32)) bits_3570 (
        .y(_T_3269),
        .in(_T_3247)
    );
    wire [1:0] _T_3270;
    BITS #(.width(99), .high(35), .low(34)) bits_3571 (
        .y(_T_3270),
        .in(_T_3247)
    );
    wire [26:0] _T_3271;
    BITS #(.width(99), .high(62), .low(36)) bits_3572 (
        .y(_T_3271),
        .in(_T_3247)
    );
    wire _T_3272;
    BITS #(.width(99), .high(63), .low(63)) bits_3573 (
        .y(_T_3272),
        .in(_T_3247)
    );
    wire [1:0] _T_3273;
    BITS #(.width(99), .high(65), .low(64)) bits_3574 (
        .y(_T_3273),
        .in(_T_3247)
    );
    wire [31:0] _T_3274;
    BITS #(.width(99), .high(97), .low(66)) bits_3575 (
        .y(_T_3274),
        .in(_T_3247)
    );
    wire _T_3275;
    BITS #(.width(99), .high(98), .low(98)) bits_3576 (
        .y(_T_3275),
        .in(_T_3247)
    );
    wire _T_3277;
    wire [1:0] _WTEMP_514;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_3577 (
        .y(_WTEMP_514),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(2)) u_neq_3578 (
        .y(_T_3277),
        .a(_T_3217_fs),
        .b(_WTEMP_514)
    );
    wire _T_3278;
    BITS #(.width(1), .high(0), .low(0)) bits_3579 (
        .y(_T_3278),
        .in(_T_3277)
    );
    wire [1:0] _T_3281;
    MUX_UNSIGNED #(.width(2)) u_mux_3580 (
        .y(_T_3281),
        .sel(_T_3278),
        .a(2'h3),
        .b(2'h0)
    );
    wire [1:0] _node_82;
    MUX_UNSIGNED #(.width(2)) u_mux_3581 (
        .y(_node_82),
        .sel(_T_1485),
        .a(_T_2993),
        .b(_reg_mstatus_fs__q)
    );
    wire _node_83;
    MUX_UNSIGNED #(.width(1)) u_mux_3582 (
        .y(_node_83),
        .sel(_T_1485),
        .a(_T_2929_pum),
        .b(_reg_mstatus_pum__q)
    );
    wire _node_84;
    MUX_UNSIGNED #(.width(1)) u_mux_3583 (
        .y(_node_84),
        .sel(_T_1485),
        .a(_T_2929_sie),
        .b(_node_69)
    );
    wire _node_85;
    MUX_UNSIGNED #(.width(1)) u_mux_3584 (
        .y(_node_85),
        .sel(_T_1485),
        .a(_T_2929_spie),
        .b(_node_70)
    );
    wire [1:0] _node_86;
    wire [1:0] _WTEMP_515;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_3585 (
        .y(_WTEMP_515),
        .in(_T_2929_spp)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_3586 (
        .y(_node_86),
        .sel(_T_1485),
        .a(_WTEMP_515),
        .b(_node_71)
    );
    wire _T_3310_rocc;
    wire _T_3310_meip;
    wire _T_3310_heip;
    wire _T_3310_seip;
    wire _T_3310_ueip;
    wire _T_3310_mtip;
    wire _T_3310_htip;
    wire _T_3310_stip;
    wire _T_3310_utip;
    wire _T_3310_msip;
    wire _T_3310_hsip;
    wire _T_3310_ssip;
    wire _T_3310_usip;
    wire [12:0] _T_3325;
    wire _T_3326;
    BITS #(.width(13), .high(0), .low(0)) bits_3587 (
        .y(_T_3326),
        .in(_T_3325)
    );
    wire _T_3327;
    BITS #(.width(13), .high(1), .low(1)) bits_3588 (
        .y(_T_3327),
        .in(_T_3325)
    );
    wire _T_3328;
    BITS #(.width(13), .high(2), .low(2)) bits_3589 (
        .y(_T_3328),
        .in(_T_3325)
    );
    wire _T_3329;
    BITS #(.width(13), .high(3), .low(3)) bits_3590 (
        .y(_T_3329),
        .in(_T_3325)
    );
    wire _T_3330;
    BITS #(.width(13), .high(4), .low(4)) bits_3591 (
        .y(_T_3330),
        .in(_T_3325)
    );
    wire _T_3331;
    BITS #(.width(13), .high(5), .low(5)) bits_3592 (
        .y(_T_3331),
        .in(_T_3325)
    );
    wire _T_3332;
    BITS #(.width(13), .high(6), .low(6)) bits_3593 (
        .y(_T_3332),
        .in(_T_3325)
    );
    wire _T_3333;
    BITS #(.width(13), .high(7), .low(7)) bits_3594 (
        .y(_T_3333),
        .in(_T_3325)
    );
    wire _T_3334;
    BITS #(.width(13), .high(8), .low(8)) bits_3595 (
        .y(_T_3334),
        .in(_T_3325)
    );
    wire _T_3335;
    BITS #(.width(13), .high(9), .low(9)) bits_3596 (
        .y(_T_3335),
        .in(_T_3325)
    );
    wire _T_3336;
    BITS #(.width(13), .high(10), .low(10)) bits_3597 (
        .y(_T_3336),
        .in(_T_3325)
    );
    wire _T_3337;
    BITS #(.width(13), .high(11), .low(11)) bits_3598 (
        .y(_T_3337),
        .in(_T_3325)
    );
    wire _T_3338;
    BITS #(.width(13), .high(12), .low(12)) bits_3599 (
        .y(_T_3338),
        .in(_T_3325)
    );
    wire _node_87;
    MUX_UNSIGNED #(.width(1)) u_mux_3600 (
        .y(_node_87),
        .sel(_T_1489),
        .a(_T_3034_ssip),
        .b(_reg_mip_ssip__q)
    );
    wire [3:0] _T_3347_mode;
    wire [15:0] _T_3347_asid;
    wire [43:0] _T_3347_ppn;
    wire [63:0] _T_3352;
    wire [43:0] _T_3353;
    BITS #(.width(64), .high(43), .low(0)) bits_3601 (
        .y(_T_3353),
        .in(_T_3352)
    );
    wire [15:0] _T_3354;
    BITS #(.width(64), .high(59), .low(44)) bits_3602 (
        .y(_T_3354),
        .in(_T_3352)
    );
    wire [3:0] _T_3355;
    BITS #(.width(64), .high(63), .low(60)) bits_3603 (
        .y(_T_3355),
        .in(_T_3352)
    );
    wire _T_3357;
    wire [3:0] _WTEMP_516;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_3604 (
        .y(_WTEMP_516),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(4)) u_eq_3605 (
        .y(_T_3357),
        .a(_T_3347_mode),
        .b(_WTEMP_516)
    );
    wire _T_3360;
    EQ_UNSIGNED #(.width(4)) u_eq_3606 (
        .y(_T_3360),
        .a(_T_3347_mode),
        .b(4'h8)
    );
    wire [3:0] _node_88;
    wire [3:0] _WTEMP_517;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_3607 (
        .y(_WTEMP_517),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(4)) u_mux_3608 (
        .y(_node_88),
        .sel(_T_3357),
        .a(_WTEMP_517),
        .b(_reg_sptbr_mode__q)
    );
    wire _T_3363;
    wire [3:0] _WTEMP_518;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_3609 (
        .y(_WTEMP_518),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(4)) u_eq_3610 (
        .y(_T_3363),
        .a(_T_3347_mode),
        .b(_WTEMP_518)
    );
    wire _T_3365;
    EQ_UNSIGNED #(.width(4)) u_eq_3611 (
        .y(_T_3365),
        .a(_T_3347_mode),
        .b(4'h8)
    );
    wire _T_3366;
    BITWISEOR #(.width(1)) bitwiseor_3612 (
        .y(_T_3366),
        .a(_T_3363),
        .b(_T_3365)
    );
    wire [19:0] _T_3367;
    BITS #(.width(44), .high(19), .low(0)) bits_3613 (
        .y(_T_3367),
        .in(_T_3347_ppn)
    );
    wire [3:0] _node_89;
    MUX_UNSIGNED #(.width(4)) u_mux_3614 (
        .y(_node_89),
        .sel(_T_3360),
        .a(4'h8),
        .b(_node_88)
    );
    wire [43:0] _node_90;
    wire [43:0] _WTEMP_519;
    PAD_UNSIGNED #(.width(20), .n(44)) u_pad_3615 (
        .y(_WTEMP_519),
        .in(_T_3367)
    );
    MUX_UNSIGNED #(.width(44)) u_mux_3616 (
        .y(_node_90),
        .sel(_T_3366),
        .a(_WTEMP_519),
        .b(_reg_sptbr_ppn__q)
    );
    wire [63:0] _T_3368;
    BITWISENOT #(.width(64)) bitwisenot_3617 (
        .y(_T_3368),
        .in(_reg_mideleg__q)
    );
    wire [63:0] _T_3369;
    BITWISEAND #(.width(64)) bitwiseand_3618 (
        .y(_T_3369),
        .a(_reg_mie__q),
        .b(_T_3368)
    );
    wire [63:0] _T_3370;
    BITWISEAND #(.width(64)) bitwiseand_3619 (
        .y(_T_3370),
        .a(wdata),
        .b(_reg_mideleg__q)
    );
    wire [63:0] _T_3371;
    BITWISEOR #(.width(64)) bitwiseor_3620 (
        .y(_T_3371),
        .a(_T_3369),
        .b(_T_3370)
    );
    wire [63:0] _node_91;
    MUX_UNSIGNED #(.width(64)) u_mux_3621 (
        .y(_node_91),
        .sel(_T_1491),
        .a(_T_3063),
        .b(_reg_mie__q)
    );
    wire [63:0] _T_3372;
    BITWISENOT #(.width(64)) bitwisenot_3622 (
        .y(_T_3372),
        .in(wdata)
    );
    wire _T_3373;
    BITS #(.width(64), .high(2), .low(2)) bits_3623 (
        .y(_T_3373),
        .in(_reg_misa__q)
    );
    wire _T_3375;
    EQ_UNSIGNED #(.width(1)) u_eq_3624 (
        .y(_T_3375),
        .a(_T_3373),
        .b(1'h0)
    );
    wire [1:0] _T_3377;
    CAT #(.width_a(1), .width_b(1)) cat_3625 (
        .y(_T_3377),
        .a(_T_3375),
        .b(1'h1)
    );
    wire [63:0] _T_3378;
    wire [63:0] _WTEMP_520;
    PAD_UNSIGNED #(.width(2), .n(64)) u_pad_3626 (
        .y(_WTEMP_520),
        .in(_T_3377)
    );
    BITWISEOR #(.width(64)) bitwiseor_3627 (
        .y(_T_3378),
        .a(_T_3372),
        .b(_WTEMP_520)
    );
    wire [63:0] _T_3379;
    BITWISENOT #(.width(64)) bitwisenot_3628 (
        .y(_T_3379),
        .in(_T_3378)
    );
    wire [39:0] _node_92;
    MUX_UNSIGNED #(.width(40)) u_mux_3629 (
        .y(_node_92),
        .sel(exception),
        .a(_node_29),
        .b(_reg_sepc__q)
    );
    wire [61:0] _T_3380;
    SHR_UNSIGNED #(.width(64), .n(2)) u_shr_3630 (
        .y(_T_3380),
        .in(wdata)
    );
    wire [63:0] _T_3381;
    SHL_UNSIGNED #(.width(62), .n(2)) u_shl_3631 (
        .y(_T_3381),
        .in(_T_3380)
    );
    wire [63:0] _T_3383;
    BITWISEAND #(.width(64)) bitwiseand_3632 (
        .y(_T_3383),
        .a(wdata),
        .b(64'h800000000000001F)
    );
    wire [63:0] _node_93;
    MUX_UNSIGNED #(.width(64)) u_mux_3633 (
        .y(_node_93),
        .sel(exception),
        .a(_node_28),
        .b(_reg_scause__q)
    );
    wire [39:0] _T_3384;
    BITS #(.width(64), .high(39), .low(0)) bits_3634 (
        .y(_T_3384),
        .in(wdata)
    );
    wire [39:0] _node_94;
    MUX_UNSIGNED #(.width(40)) u_mux_3635 (
        .y(_node_94),
        .sel(exception),
        .a(_node_27),
        .b(_reg_sbadaddr__q)
    );
    wire [63:0] _T_3385;
    wire [63:0] _WTEMP_521;
    PAD_UNSIGNED #(.width(13), .n(64)) u_pad_3636 (
        .y(_WTEMP_521),
        .in(delegable_interrupts)
    );
    BITWISEAND #(.width(64)) bitwiseand_3637 (
        .y(_T_3385),
        .a(wdata),
        .b(_WTEMP_521)
    );
    wire [63:0] _T_3386;
    wire [63:0] _WTEMP_522;
    PAD_UNSIGNED #(.width(9), .n(64)) u_pad_3638 (
        .y(_WTEMP_522),
        .in(9'h1AB)
    );
    BITWISEAND #(.width(64)) bitwiseand_3639 (
        .y(_T_3386),
        .a(wdata),
        .b(_WTEMP_522)
    );
    wire [63:0] _T_3388;
    wire [63:0] _WTEMP_523;
    PAD_UNSIGNED #(.width(3), .n(64)) u_pad_3640 (
        .y(_WTEMP_523),
        .in(3'h7)
    );
    BITWISEAND #(.width(64)) bitwiseand_3641 (
        .y(_T_3388),
        .a(wdata),
        .b(_WTEMP_523)
    );
    wire [63:0] _T_3390;
    wire [63:0] _WTEMP_524;
    PAD_UNSIGNED #(.width(3), .n(64)) u_pad_3642 (
        .y(_WTEMP_524),
        .in(3'h7)
    );
    BITWISEAND #(.width(64)) bitwiseand_3643 (
        .y(_T_3390),
        .a(wdata),
        .b(_WTEMP_524)
    );
    wire _T_3427;
    EQ_UNSIGNED #(.width(1)) u_eq_3644 (
        .y(_T_3427),
        .a(_reg_bp_0_control_dmode__q),
        .b(1'h0)
    );
    wire _T_3428;
    BITWISEOR #(.width(1)) bitwiseor_3645 (
        .y(_T_3428),
        .a(_T_3427),
        .b(_reg_debug__q)
    );
    wire [3:0] _T_3461_ttype;
    wire _T_3461_dmode;
    wire [5:0] _T_3461_maskmax;
    wire [39:0] _T_3461_reserved;
    wire _T_3461_action;
    wire _T_3461_chain;
    wire [1:0] _T_3461_zero;
    wire [1:0] _T_3461_tmatch;
    wire _T_3461_m;
    wire _T_3461_h;
    wire _T_3461_s;
    wire _T_3461_u;
    wire _T_3461_x;
    wire _T_3461_w;
    wire _T_3461_r;
    wire [63:0] _T_3478;
    wire _T_3479;
    BITS #(.width(64), .high(0), .low(0)) bits_3646 (
        .y(_T_3479),
        .in(_T_3478)
    );
    wire _T_3480;
    BITS #(.width(64), .high(1), .low(1)) bits_3647 (
        .y(_T_3480),
        .in(_T_3478)
    );
    wire _T_3481;
    BITS #(.width(64), .high(2), .low(2)) bits_3648 (
        .y(_T_3481),
        .in(_T_3478)
    );
    wire _T_3482;
    BITS #(.width(64), .high(3), .low(3)) bits_3649 (
        .y(_T_3482),
        .in(_T_3478)
    );
    wire _T_3483;
    BITS #(.width(64), .high(4), .low(4)) bits_3650 (
        .y(_T_3483),
        .in(_T_3478)
    );
    wire _T_3484;
    BITS #(.width(64), .high(5), .low(5)) bits_3651 (
        .y(_T_3484),
        .in(_T_3478)
    );
    wire _T_3485;
    BITS #(.width(64), .high(6), .low(6)) bits_3652 (
        .y(_T_3485),
        .in(_T_3478)
    );
    wire [1:0] _T_3486;
    BITS #(.width(64), .high(8), .low(7)) bits_3653 (
        .y(_T_3486),
        .in(_T_3478)
    );
    wire [1:0] _T_3487;
    BITS #(.width(64), .high(10), .low(9)) bits_3654 (
        .y(_T_3487),
        .in(_T_3478)
    );
    wire _T_3488;
    BITS #(.width(64), .high(11), .low(11)) bits_3655 (
        .y(_T_3488),
        .in(_T_3478)
    );
    wire _T_3489;
    BITS #(.width(64), .high(12), .low(12)) bits_3656 (
        .y(_T_3489),
        .in(_T_3478)
    );
    wire [39:0] _T_3490;
    BITS #(.width(64), .high(52), .low(13)) bits_3657 (
        .y(_T_3490),
        .in(_T_3478)
    );
    wire [5:0] _T_3491;
    BITS #(.width(64), .high(58), .low(53)) bits_3658 (
        .y(_T_3491),
        .in(_T_3478)
    );
    wire _T_3492;
    BITS #(.width(64), .high(59), .low(59)) bits_3659 (
        .y(_T_3492),
        .in(_T_3478)
    );
    wire [3:0] _T_3493;
    BITS #(.width(64), .high(63), .low(60)) bits_3660 (
        .y(_T_3493),
        .in(_T_3478)
    );
    wire _T_3494;
    BITWISEAND #(.width(1)) bitwiseand_3661 (
        .y(_T_3494),
        .a(_T_3461_dmode),
        .b(_reg_debug__q)
    );
    wire _T_3495;
    BITWISEAND #(.width(1)) bitwiseand_3662 (
        .y(_T_3495),
        .a(_T_3494),
        .b(_T_3461_action)
    );
    wire _node_95;
    assign _node_95 = _T_3489;
    wire _node_96;
    assign _node_96 = _T_3488;
    wire _node_97;
    assign _node_97 = _T_3492;
    wire _node_98;
    assign _node_98 = _T_3484;
    wire _node_99;
    assign _node_99 = _T_3485;
    wire [5:0] _node_100;
    assign _node_100 = _T_3491;
    wire _node_101;
    assign _node_101 = _T_3479;
    wire [39:0] _node_102;
    assign _node_102 = _T_3490;
    wire _node_103;
    assign _node_103 = _T_3483;
    wire [1:0] _node_104;
    assign _node_104 = _T_3486;
    wire [3:0] _node_105;
    assign _node_105 = _T_3493;
    wire _node_106;
    assign _node_106 = _T_3482;
    wire _node_107;
    assign _node_107 = _T_3480;
    wire _node_108;
    assign _node_108 = _T_3481;
    wire [1:0] _node_109;
    assign _node_109 = _T_3487;
    wire [63:0] _node_110;
    assign _node_110 = wdata;
    wire [63:0] _node_111;
    wire [63:0] _WTEMP_525;
    PAD_UNSIGNED #(.width(39), .n(64)) u_pad_3663 (
        .y(_WTEMP_525),
        .in(_reg_bp_0_address__q)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_3664 (
        .y(_node_111),
        .sel(_T_1471),
        .a(wdata),
        .b(_WTEMP_525)
    );
    wire _node_112;
    MUX_UNSIGNED #(.width(1)) u_mux_3665 (
        .y(_node_112),
        .sel(_T_1469),
        .a(_T_3495),
        .b(_reg_bp_0_control_action__q)
    );
    wire _node_113;
    MUX_UNSIGNED #(.width(1)) u_mux_3666 (
        .y(_node_113),
        .sel(_T_1469),
        .a(_T_3494),
        .b(_reg_bp_0_control_dmode__q)
    );
    wire _node_114;
    MUX_UNSIGNED #(.width(1)) u_mux_3667 (
        .y(_node_114),
        .sel(_T_1469),
        .a(_T_3461_m),
        .b(_reg_bp_0_control_m__q)
    );
    wire _node_115;
    MUX_UNSIGNED #(.width(1)) u_mux_3668 (
        .y(_node_115),
        .sel(_T_1469),
        .a(_T_3461_r),
        .b(_reg_bp_0_control_r__q)
    );
    wire _node_116;
    MUX_UNSIGNED #(.width(1)) u_mux_3669 (
        .y(_node_116),
        .sel(_T_1469),
        .a(_T_3461_s),
        .b(_reg_bp_0_control_s__q)
    );
    wire [1:0] _node_117;
    MUX_UNSIGNED #(.width(2)) u_mux_3670 (
        .y(_node_117),
        .sel(_T_1469),
        .a(_T_3461_tmatch),
        .b(_reg_bp_0_control_tmatch__q)
    );
    wire _node_118;
    MUX_UNSIGNED #(.width(1)) u_mux_3671 (
        .y(_node_118),
        .sel(_T_1469),
        .a(_T_3461_u),
        .b(_reg_bp_0_control_u__q)
    );
    wire _node_119;
    MUX_UNSIGNED #(.width(1)) u_mux_3672 (
        .y(_node_119),
        .sel(_T_1469),
        .a(_T_3461_w),
        .b(_reg_bp_0_control_w__q)
    );
    wire _node_120;
    MUX_UNSIGNED #(.width(1)) u_mux_3673 (
        .y(_node_120),
        .sel(_T_1469),
        .a(_T_3461_x),
        .b(_reg_bp_0_control_x__q)
    );
    wire _node_121;
    assign _node_121 = _T_2987;
    wire [1:0] _node_122;
    assign _node_122 = _T_2971;
    wire _node_123;
    assign _node_123 = _T_2962;
    wire _node_124;
    assign _node_124 = _T_2966;
    wire [1:0] _node_125;
    assign _node_125 = _T_2969;
    wire [31:0] _node_126;
    assign _node_126 = _T_2986;
    wire _node_127;
    assign _node_127 = _T_2963;
    wire _node_128;
    assign _node_128 = _T_2967;
    wire [1:0] _node_129;
    assign _node_129 = _T_2970;
    wire _node_130;
    assign _node_130 = _T_2973;
    wire _node_131;
    assign _node_131 = _T_2975;
    wire [1:0] _node_132;
    assign _node_132 = _T_2985;
    wire _node_133;
    assign _node_133 = _T_2974;
    wire _node_134;
    assign _node_134 = _T_2984;
    wire _node_135;
    assign _node_135 = _T_2980;
    wire _node_136;
    assign _node_136 = _T_2961;
    wire _node_137;
    assign _node_137 = _T_2965;
    wire _node_138;
    assign _node_138 = _T_2968;
    wire [1:0] _node_139;
    assign _node_139 = _T_2982;
    wire _node_140;
    assign _node_140 = _T_2978;
    wire _node_141;
    assign _node_141 = _T_2976;
    wire _node_142;
    assign _node_142 = _T_2977;
    wire _node_143;
    assign _node_143 = _T_2960;
    wire _node_144;
    assign _node_144 = _T_2964;
    wire [1:0] _node_145;
    assign _node_145 = _T_2981;
    wire [1:0] _node_146;
    assign _node_146 = _T_2972;
    wire [7:0] _node_147;
    assign _node_147 = _T_2979;
    wire [26:0] _node_148;
    assign _node_148 = _T_2983;
    wire [63:0] _node_149;
    assign _node_149 = wdata;
    wire _node_150;
    assign _node_150 = _T_3060;
    wire _node_151;
    assign _node_151 = _T_3052;
    wire _node_152;
    assign _node_152 = _T_3056;
    wire _node_153;
    assign _node_153 = _T_3061;
    wire _node_154;
    assign _node_154 = _T_3053;
    wire _node_155;
    assign _node_155 = _T_3057;
    wire _node_156;
    assign _node_156 = _T_3062;
    wire _node_157;
    assign _node_157 = _T_3059;
    wire _node_158;
    assign _node_158 = _T_3051;
    wire _node_159;
    assign _node_159 = _T_3055;
    wire _node_160;
    assign _node_160 = _T_3058;
    wire _node_161;
    assign _node_161 = _T_3050;
    wire _node_162;
    assign _node_162 = _T_3054;
    wire [63:0] _node_163;
    assign _node_163 = wdata;
    wire [2:0] _node_164;
    assign _node_164 = _T_3143;
    wire _node_165;
    assign _node_165 = _T_3142;
    wire _node_166;
    assign _node_166 = _T_3149;
    wire _node_167;
    assign _node_167 = _T_3150;
    wire _node_168;
    assign _node_168 = _T_3148;
    wire _node_169;
    assign _node_169 = _T_3147;
    wire _node_170;
    assign _node_170 = _T_3152;
    wire _node_171;
    assign _node_171 = _T_3140;
    wire _node_172;
    assign _node_172 = _T_3153;
    wire [1:0] _node_173;
    assign _node_173 = _T_3138;
    wire _node_174;
    assign _node_174 = _T_3139;
    wire _node_175;
    assign _node_175 = _T_3145;
    wire _node_176;
    assign _node_176 = _T_3144;
    wire [1:0] _node_177;
    assign _node_177 = _T_3154;
    wire _node_178;
    assign _node_178 = _T_3141;
    wire _node_179;
    assign _node_179 = _T_3146;
    wire [11:0] _node_180;
    assign _node_180 = _T_3151;
    wire [63:0] _node_181;
    assign _node_181 = wdata;
    wire _node_182;
    assign _node_182 = _T_3275;
    wire [1:0] _node_183;
    assign _node_183 = _T_3259;
    wire _node_184;
    assign _node_184 = _T_3250;
    wire _node_185;
    assign _node_185 = _T_3254;
    wire [1:0] _node_186;
    assign _node_186 = _T_3257;
    wire [31:0] _node_187;
    assign _node_187 = _T_3274;
    wire _node_188;
    assign _node_188 = _T_3251;
    wire _node_189;
    assign _node_189 = _T_3255;
    wire [1:0] _node_190;
    assign _node_190 = _T_3258;
    wire _node_191;
    assign _node_191 = _T_3261;
    wire _node_192;
    assign _node_192 = _T_3263;
    wire [1:0] _node_193;
    assign _node_193 = _T_3273;
    wire _node_194;
    assign _node_194 = _T_3262;
    wire _node_195;
    assign _node_195 = _T_3272;
    wire _node_196;
    assign _node_196 = _T_3268;
    wire _node_197;
    assign _node_197 = _T_3249;
    wire _node_198;
    assign _node_198 = _T_3253;
    wire _node_199;
    assign _node_199 = _T_3256;
    wire [1:0] _node_200;
    assign _node_200 = _T_3270;
    wire _node_201;
    assign _node_201 = _T_3266;
    wire _node_202;
    assign _node_202 = _T_3264;
    wire _node_203;
    assign _node_203 = _T_3265;
    wire _node_204;
    assign _node_204 = _T_3248;
    wire _node_205;
    assign _node_205 = _T_3252;
    wire [1:0] _node_206;
    assign _node_206 = _T_3269;
    wire [1:0] _node_207;
    assign _node_207 = _T_3260;
    wire [7:0] _node_208;
    assign _node_208 = _T_3267;
    wire [26:0] _node_209;
    assign _node_209 = _T_3271;
    wire [63:0] _node_210;
    assign _node_210 = wdata;
    wire _node_211;
    assign _node_211 = _T_3336;
    wire _node_212;
    assign _node_212 = _T_3328;
    wire _node_213;
    assign _node_213 = _T_3332;
    wire _node_214;
    assign _node_214 = _T_3337;
    wire _node_215;
    assign _node_215 = _T_3329;
    wire _node_216;
    assign _node_216 = _T_3333;
    wire _node_217;
    assign _node_217 = _T_3338;
    wire _node_218;
    assign _node_218 = _T_3335;
    wire _node_219;
    assign _node_219 = _T_3327;
    wire _node_220;
    assign _node_220 = _T_3331;
    wire _node_221;
    assign _node_221 = _T_3334;
    wire _node_222;
    assign _node_222 = _T_3326;
    wire _node_223;
    assign _node_223 = _T_3330;
    wire [63:0] _node_224;
    assign _node_224 = wdata;
    wire [15:0] _node_225;
    assign _node_225 = _T_3354;
    wire [3:0] _node_226;
    assign _node_226 = _T_3355;
    wire [43:0] _node_227;
    assign _node_227 = _T_3353;
    wire [63:0] _node_228;
    assign _node_228 = wdata;
    wire _node_229;
    assign _node_229 = _node_95;
    wire _node_230;
    assign _node_230 = _node_96;
    wire _node_231;
    assign _node_231 = _node_97;
    wire _node_232;
    assign _node_232 = _node_98;
    wire _node_233;
    assign _node_233 = _node_99;
    wire [5:0] _node_234;
    assign _node_234 = _node_100;
    wire _node_235;
    assign _node_235 = _node_101;
    wire [39:0] _node_236;
    assign _node_236 = _node_102;
    wire _node_237;
    assign _node_237 = _node_103;
    wire [1:0] _node_238;
    assign _node_238 = _node_104;
    wire [3:0] _node_239;
    assign _node_239 = _node_105;
    wire _node_240;
    assign _node_240 = _node_106;
    wire _node_241;
    assign _node_241 = _node_107;
    wire _node_242;
    assign _node_242 = _node_108;
    wire [1:0] _node_243;
    assign _node_243 = _node_109;
    wire [63:0] _node_244;
    assign _node_244 = _node_110;
    wire [63:0] _node_245;
    wire [63:0] _WTEMP_526;
    PAD_UNSIGNED #(.width(7), .n(64)) u_pad_3674 (
        .y(_WTEMP_526),
        .in(_T_932)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_3675 (
        .y(_node_245),
        .sel(_T_1481),
        .a(_T_3079),
        .b(_WTEMP_526)
    );
    wire [57:0] _node_246;
    MUX_UNSIGNED #(.width(58)) u_mux_3676 (
        .y(_node_246),
        .sel(_T_1481),
        .a(_T_3080),
        .b(_node_76)
    );
    wire [57:0] _node_247;
    MUX_UNSIGNED #(.width(58)) u_mux_3677 (
        .y(_node_247),
        .sel(_T_935),
        .a(_T_938),
        .b(__T_934__q)
    );
    wire [63:0] _node_248;
    wire [63:0] _WTEMP_527;
    PAD_UNSIGNED #(.width(7), .n(64)) u_pad_3678 (
        .y(_WTEMP_527),
        .in(_T_943)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_3679 (
        .y(_node_248),
        .sel(_T_1479),
        .a(_T_3077),
        .b(_WTEMP_527)
    );
    wire [57:0] _node_249;
    MUX_UNSIGNED #(.width(58)) u_mux_3680 (
        .y(_node_249),
        .sel(_T_1479),
        .a(_T_3078),
        .b(_node_75)
    );
    wire [57:0] _node_250;
    MUX_UNSIGNED #(.width(58)) u_mux_3681 (
        .y(_node_250),
        .sel(_T_946),
        .a(_T_949),
        .b(__T_945__q)
    );
    wire [63:0] _node_251;
    wire [63:0] _WTEMP_528;
    PAD_UNSIGNED #(.width(39), .n(64)) u_pad_3682 (
        .y(_WTEMP_528),
        .in(_reg_bp_0_address__q)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_3683 (
        .y(_node_251),
        .sel(_T_3428),
        .a(_node_111),
        .b(_WTEMP_528)
    );
    wire _node_252;
    MUX_UNSIGNED #(.width(1)) u_mux_3684 (
        .y(_node_252),
        .sel(_T_3428),
        .a(_node_112),
        .b(_reg_bp_0_control_action__q)
    );
    wire _node_253;
    MUX_UNSIGNED #(.width(1)) u_mux_3685 (
        .y(_node_253),
        .sel(_T_3428),
        .a(_node_113),
        .b(_reg_bp_0_control_dmode__q)
    );
    wire _node_254;
    MUX_UNSIGNED #(.width(1)) u_mux_3686 (
        .y(_node_254),
        .sel(_T_3428),
        .a(_node_114),
        .b(_reg_bp_0_control_m__q)
    );
    wire _node_255;
    MUX_UNSIGNED #(.width(1)) u_mux_3687 (
        .y(_node_255),
        .sel(_T_3428),
        .a(_node_115),
        .b(_reg_bp_0_control_r__q)
    );
    wire _node_256;
    MUX_UNSIGNED #(.width(1)) u_mux_3688 (
        .y(_node_256),
        .sel(_T_3428),
        .a(_node_116),
        .b(_reg_bp_0_control_s__q)
    );
    wire [1:0] _node_257;
    MUX_UNSIGNED #(.width(2)) u_mux_3689 (
        .y(_node_257),
        .sel(_T_3428),
        .a(_node_117),
        .b(_reg_bp_0_control_tmatch__q)
    );
    wire _node_258;
    MUX_UNSIGNED #(.width(1)) u_mux_3690 (
        .y(_node_258),
        .sel(_T_3428),
        .a(_node_118),
        .b(_reg_bp_0_control_u__q)
    );
    wire _node_259;
    MUX_UNSIGNED #(.width(1)) u_mux_3691 (
        .y(_node_259),
        .sel(_T_3428),
        .a(_node_119),
        .b(_reg_bp_0_control_w__q)
    );
    wire _node_260;
    MUX_UNSIGNED #(.width(1)) u_mux_3692 (
        .y(_node_260),
        .sel(_T_3428),
        .a(_node_120),
        .b(_reg_bp_0_control_x__q)
    );
    wire _node_261;
    MUX_UNSIGNED #(.width(1)) u_mux_3693 (
        .y(_node_261),
        .sel(_T_1507),
        .a(_T_3118_ebreakm),
        .b(_reg_dcsr_ebreakm__q)
    );
    wire _node_262;
    MUX_UNSIGNED #(.width(1)) u_mux_3694 (
        .y(_node_262),
        .sel(_T_1507),
        .a(_T_3118_ebreaks),
        .b(_reg_dcsr_ebreaks__q)
    );
    wire _node_263;
    MUX_UNSIGNED #(.width(1)) u_mux_3695 (
        .y(_node_263),
        .sel(_T_1507),
        .a(_T_3118_ebreaku),
        .b(_reg_dcsr_ebreaku__q)
    );
    wire _node_264;
    MUX_UNSIGNED #(.width(1)) u_mux_3696 (
        .y(_node_264),
        .sel(_T_1507),
        .a(_T_3118_halt),
        .b(_reg_dcsr_halt__q)
    );
    wire [1:0] _node_265;
    MUX_UNSIGNED #(.width(2)) u_mux_3697 (
        .y(_node_265),
        .sel(_T_1507),
        .a(_T_3118_prv),
        .b(_node_80)
    );
    wire [1:0] _node_266;
    MUX_UNSIGNED #(.width(2)) u_mux_3698 (
        .y(_node_266),
        .sel(exception),
        .a(_node_15),
        .b(_reg_dcsr_prv__q)
    );
    wire _node_267;
    MUX_UNSIGNED #(.width(1)) u_mux_3699 (
        .y(_node_267),
        .sel(_T_1507),
        .a(_T_3118_step),
        .b(_reg_dcsr_step__q)
    );
    wire [63:0] _node_268;
    wire [63:0] _WTEMP_529;
    PAD_UNSIGNED #(.width(40), .n(64)) u_pad_3700 (
        .y(_WTEMP_529),
        .in(_node_81)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_3701 (
        .y(_node_268),
        .sel(_T_1509),
        .a(_T_3158),
        .b(_WTEMP_529)
    );
    wire [39:0] _node_269;
    MUX_UNSIGNED #(.width(40)) u_mux_3702 (
        .y(_node_269),
        .sel(exception),
        .a(_node_17),
        .b(_reg_dpc__q)
    );
    wire [63:0] _node_270;
    MUX_UNSIGNED #(.width(64)) u_mux_3703 (
        .y(_node_270),
        .sel(_T_1511),
        .a(wdata),
        .b(_reg_dscratch__q)
    );
    wire [63:0] _node_271;
    MUX_UNSIGNED #(.width(64)) u_mux_3704 (
        .y(_node_271),
        .sel(_T_1517),
        .a(wdata),
        .b(_node_78)
    );
    wire [4:0] _node_272;
    MUX_UNSIGNED #(.width(5)) u_mux_3705 (
        .y(_node_272),
        .sel(io_fcsr_flags_valid),
        .a(_T_2862),
        .b(_reg_fflags__q)
    );
    wire [63:0] _node_273;
    wire [63:0] _WTEMP_530;
    PAD_UNSIGNED #(.width(59), .n(64)) u_pad_3706 (
        .y(_WTEMP_530),
        .in(_T_3081)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_3707 (
        .y(_node_273),
        .sel(_T_1517),
        .a(_WTEMP_530),
        .b(_node_79)
    );
    wire [39:0] _node_274;
    MUX_UNSIGNED #(.width(40)) u_mux_3708 (
        .y(_node_274),
        .sel(_T_1501),
        .a(_T_3076),
        .b(_node_74)
    );
    wire [39:0] _node_275;
    MUX_UNSIGNED #(.width(40)) u_mux_3709 (
        .y(_node_275),
        .sel(exception),
        .a(_node_18),
        .b(_reg_mbadaddr__q)
    );
    wire [63:0] _node_276;
    MUX_UNSIGNED #(.width(64)) u_mux_3710 (
        .y(_node_276),
        .sel(_T_1503),
        .a(_T_3075),
        .b(_node_73)
    );
    wire [63:0] _node_277;
    MUX_UNSIGNED #(.width(64)) u_mux_3711 (
        .y(_node_277),
        .sel(exception),
        .a(_node_19),
        .b(_reg_mcause__q)
    );
    wire [63:0] _node_278;
    wire [63:0] _WTEMP_531;
    PAD_UNSIGNED #(.width(32), .n(64)) u_pad_3712 (
        .y(_WTEMP_531),
        .in(_reg_mcounteren__q)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_3713 (
        .y(_node_278),
        .sel(_T_1713),
        .a(_T_3390),
        .b(_WTEMP_531)
    );
    wire [63:0] _node_279;
    MUX_UNSIGNED #(.width(64)) u_mux_3714 (
        .y(_node_279),
        .sel(_T_1495),
        .a(_T_3386),
        .b(_reg_medeleg__q)
    );
    wire [63:0] _node_280;
    wire [63:0] _WTEMP_532;
    PAD_UNSIGNED #(.width(40), .n(64)) u_pad_3715 (
        .y(_WTEMP_532),
        .in(_node_72)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_3716 (
        .y(_node_280),
        .sel(_T_1499),
        .a(_T_3071),
        .b(_WTEMP_532)
    );
    wire [39:0] _node_281;
    MUX_UNSIGNED #(.width(40)) u_mux_3717 (
        .y(_node_281),
        .sel(exception),
        .a(_node_20),
        .b(_reg_mepc__q)
    );
    wire [63:0] _node_282;
    MUX_UNSIGNED #(.width(64)) u_mux_3718 (
        .y(_node_282),
        .sel(_T_1493),
        .a(_T_3385),
        .b(_reg_mideleg__q)
    );
    wire [63:0] _node_283;
    MUX_UNSIGNED #(.width(64)) u_mux_3719 (
        .y(_node_283),
        .sel(_T_1697),
        .a(_T_3371),
        .b(_node_91)
    );
    wire _node_284;
    MUX_UNSIGNED #(.width(1)) u_mux_3720 (
        .y(_node_284),
        .sel(_T_1695),
        .a(_T_3310_ssip),
        .b(_node_87)
    );
    wire _node_285;
    MUX_UNSIGNED #(.width(1)) u_mux_3721 (
        .y(_node_285),
        .sel(_T_1489),
        .a(_T_3034_stip),
        .b(_reg_mip_stip__q)
    );
    wire [63:0] _node_286;
    MUX_UNSIGNED #(.width(64)) u_mux_3722 (
        .y(_node_286),
        .sel(_T_1483),
        .a(_T_3005),
        .b(_reg_misa__q)
    );
    wire [63:0] _node_287;
    MUX_UNSIGNED #(.width(64)) u_mux_3723 (
        .y(_node_287),
        .sel(_T_1497),
        .a(wdata),
        .b(_reg_mscratch__q)
    );
    wire [1:0] _node_288;
    MUX_UNSIGNED #(.width(2)) u_mux_3724 (
        .y(_node_288),
        .sel(_T_1693),
        .a(_T_3281),
        .b(_node_82)
    );
    wire _node_289;
    MUX_UNSIGNED #(.width(1)) u_mux_3725 (
        .y(_node_289),
        .sel(_T_1485),
        .a(_T_2929_mie),
        .b(_node_66)
    );
    wire _node_290;
    MUX_UNSIGNED #(.width(1)) u_mux_3726 (
        .y(_node_290),
        .sel(insn_ret),
        .a(_node_54),
        .b(_node_55)
    );
    wire _node_291;
    MUX_UNSIGNED #(.width(1)) u_mux_3727 (
        .y(_node_291),
        .sel(_T_1485),
        .a(_T_2929_mpie),
        .b(_node_67)
    );
    wire _node_292;
    MUX_UNSIGNED #(.width(1)) u_mux_3728 (
        .y(_node_292),
        .sel(insn_ret),
        .a(_node_56),
        .b(_node_57)
    );
    wire [1:0] _node_293;
    MUX_UNSIGNED #(.width(2)) u_mux_3729 (
        .y(_node_293),
        .sel(_T_1485),
        .a(_T_2929_mpp),
        .b(_node_68)
    );
    wire [1:0] _node_294;
    MUX_UNSIGNED #(.width(2)) u_mux_3730 (
        .y(_node_294),
        .sel(insn_ret),
        .a(_node_58),
        .b(_node_59)
    );
    wire _node_295;
    MUX_UNSIGNED #(.width(1)) u_mux_3731 (
        .y(_node_295),
        .sel(_T_1485),
        .a(_T_2929_mprv),
        .b(_reg_mstatus_mprv__q)
    );
    wire _node_296;
    MUX_UNSIGNED #(.width(1)) u_mux_3732 (
        .y(_node_296),
        .sel(_T_1485),
        .a(_T_2929_mxr),
        .b(_reg_mstatus_mxr__q)
    );
    wire _node_297;
    MUX_UNSIGNED #(.width(1)) u_mux_3733 (
        .y(_node_297),
        .sel(_T_1693),
        .a(_T_3217_pum),
        .b(_node_83)
    );
    wire _node_298;
    MUX_UNSIGNED #(.width(1)) u_mux_3734 (
        .y(_node_298),
        .sel(_T_1693),
        .a(_T_3217_sie),
        .b(_node_84)
    );
    wire _node_299;
    MUX_UNSIGNED #(.width(1)) u_mux_3735 (
        .y(_node_299),
        .sel(insn_ret),
        .a(_node_60),
        .b(_node_61)
    );
    wire _node_300;
    MUX_UNSIGNED #(.width(1)) u_mux_3736 (
        .y(_node_300),
        .sel(_T_1693),
        .a(_T_3217_spie),
        .b(_node_85)
    );
    wire _node_301;
    MUX_UNSIGNED #(.width(1)) u_mux_3737 (
        .y(_node_301),
        .sel(insn_ret),
        .a(_node_62),
        .b(_node_63)
    );
    wire [1:0] _node_302;
    wire [1:0] _WTEMP_533;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_3738 (
        .y(_WTEMP_533),
        .in(_T_3217_spp)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_3739 (
        .y(_node_302),
        .sel(_T_1693),
        .a(_WTEMP_533),
        .b(_node_86)
    );
    wire [1:0] _node_303;
    MUX_UNSIGNED #(.width(2)) u_mux_3740 (
        .y(_node_303),
        .sel(insn_ret),
        .a(_node_64),
        .b(_node_65)
    );
    wire _node_304;
    MUX_UNSIGNED #(.width(1)) u_mux_3741 (
        .y(_node_304),
        .sel(_T_1485),
        .a(_T_2929_tsr),
        .b(_reg_mstatus_tsr__q)
    );
    wire _node_305;
    MUX_UNSIGNED #(.width(1)) u_mux_3742 (
        .y(_node_305),
        .sel(_T_1485),
        .a(_T_2929_tvm),
        .b(_reg_mstatus_tvm__q)
    );
    wire _node_306;
    MUX_UNSIGNED #(.width(1)) u_mux_3743 (
        .y(_node_306),
        .sel(_T_1485),
        .a(_T_2929_tw),
        .b(_reg_mstatus_tw__q)
    );
    wire [63:0] _node_307;
    wire [63:0] _WTEMP_534;
    PAD_UNSIGNED #(.width(32), .n(64)) u_pad_3744 (
        .y(_WTEMP_534),
        .in(_reg_mtvec__q)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_3745 (
        .y(_node_307),
        .sel(_T_1487),
        .a(_T_3073),
        .b(_WTEMP_534)
    );
    wire [39:0] _node_308;
    MUX_UNSIGNED #(.width(40)) u_mux_3746 (
        .y(_node_308),
        .sel(_T_1703),
        .a(_T_3384),
        .b(_node_94)
    );
    wire [39:0] _node_309;
    MUX_UNSIGNED #(.width(40)) u_mux_3747 (
        .y(_node_309),
        .sel(exception),
        .a(_node_27),
        .b(_reg_sbadaddr__q)
    );
    wire [63:0] _node_310;
    MUX_UNSIGNED #(.width(64)) u_mux_3748 (
        .y(_node_310),
        .sel(_T_1701),
        .a(_T_3383),
        .b(_node_93)
    );
    wire [63:0] _node_311;
    MUX_UNSIGNED #(.width(64)) u_mux_3749 (
        .y(_node_311),
        .sel(exception),
        .a(_node_28),
        .b(_reg_scause__q)
    );
    wire [63:0] _node_312;
    wire [63:0] _WTEMP_535;
    PAD_UNSIGNED #(.width(32), .n(64)) u_pad_3750 (
        .y(_WTEMP_535),
        .in(_reg_scounteren__q)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_3751 (
        .y(_node_312),
        .sel(_T_1711),
        .a(_T_3388),
        .b(_WTEMP_535)
    );
    wire [63:0] _node_313;
    wire [63:0] _WTEMP_536;
    PAD_UNSIGNED #(.width(40), .n(64)) u_pad_3752 (
        .y(_WTEMP_536),
        .in(_node_92)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_3753 (
        .y(_node_313),
        .sel(_T_1707),
        .a(_T_3379),
        .b(_WTEMP_536)
    );
    wire [39:0] _node_314;
    MUX_UNSIGNED #(.width(40)) u_mux_3754 (
        .y(_node_314),
        .sel(exception),
        .a(_node_29),
        .b(_reg_sepc__q)
    );
    wire [3:0] _node_315;
    MUX_UNSIGNED #(.width(4)) u_mux_3755 (
        .y(_node_315),
        .sel(_T_1705),
        .a(_node_89),
        .b(_reg_sptbr_mode__q)
    );
    wire [43:0] _node_316;
    MUX_UNSIGNED #(.width(44)) u_mux_3756 (
        .y(_node_316),
        .sel(_T_1705),
        .a(_node_90),
        .b(_reg_sptbr_ppn__q)
    );
    wire [63:0] _node_317;
    MUX_UNSIGNED #(.width(64)) u_mux_3757 (
        .y(_node_317),
        .sel(_T_1699),
        .a(wdata),
        .b(_reg_sscratch__q)
    );
    wire [63:0] _node_318;
    wire [63:0] _WTEMP_537;
    PAD_UNSIGNED #(.width(39), .n(64)) u_pad_3758 (
        .y(_WTEMP_537),
        .in(_reg_stvec__q)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_3759 (
        .y(_node_318),
        .sel(_T_1709),
        .a(_T_3381),
        .b(_WTEMP_537)
    );
    wire _node_319;
    MUX_UNSIGNED #(.width(1)) u_mux_3760 (
        .y(_node_319),
        .sel(_T_2870),
        .a(_node_252),
        .b(_reg_bp_0_control_action__q)
    );
    wire _node_320;
    MUX_UNSIGNED #(.width(1)) u_mux_3761 (
        .y(_node_320),
        .sel(_T_2870),
        .a(_node_253),
        .b(_reg_bp_0_control_dmode__q)
    );
    wire _node_321;
    MUX_UNSIGNED #(.width(1)) u_mux_3762 (
        .y(_node_321),
        .sel(_T_2870),
        .a(_node_255),
        .b(_reg_bp_0_control_r__q)
    );
    wire _node_322;
    MUX_UNSIGNED #(.width(1)) u_mux_3763 (
        .y(_node_322),
        .sel(_T_2870),
        .a(_node_259),
        .b(_reg_bp_0_control_w__q)
    );
    wire _node_323;
    MUX_UNSIGNED #(.width(1)) u_mux_3764 (
        .y(_node_323),
        .sel(_T_2870),
        .a(_node_260),
        .b(_reg_bp_0_control_x__q)
    );
    wire [3:0] _T_3556_control_ttype;
    wire _T_3556_control_dmode;
    wire [5:0] _T_3556_control_maskmax;
    wire [39:0] _T_3556_control_reserved;
    wire _T_3556_control_action;
    wire _T_3556_control_chain;
    wire [1:0] _T_3556_control_zero;
    wire [1:0] _T_3556_control_tmatch;
    wire _T_3556_control_m;
    wire _T_3556_control_h;
    wire _T_3556_control_s;
    wire _T_3556_control_u;
    wire _T_3556_control_x;
    wire _T_3556_control_w;
    wire _T_3556_control_r;
    wire [38:0] _T_3556_address;
    wire [102:0] _T_3575;
    wire [38:0] _T_3576;
    BITS #(.width(103), .high(38), .low(0)) bits_3765 (
        .y(_T_3576),
        .in(_T_3575)
    );
    wire [63:0] _T_3577;
    BITS #(.width(103), .high(102), .low(39)) bits_3766 (
        .y(_T_3577),
        .in(_T_3575)
    );
    wire [63:0] _T_3579;
    wire _T_3580;
    BITS #(.width(64), .high(0), .low(0)) bits_3767 (
        .y(_T_3580),
        .in(_T_3579)
    );
    wire _T_3581;
    BITS #(.width(64), .high(1), .low(1)) bits_3768 (
        .y(_T_3581),
        .in(_T_3579)
    );
    wire _T_3582;
    BITS #(.width(64), .high(2), .low(2)) bits_3769 (
        .y(_T_3582),
        .in(_T_3579)
    );
    wire _T_3583;
    BITS #(.width(64), .high(3), .low(3)) bits_3770 (
        .y(_T_3583),
        .in(_T_3579)
    );
    wire _T_3584;
    BITS #(.width(64), .high(4), .low(4)) bits_3771 (
        .y(_T_3584),
        .in(_T_3579)
    );
    wire _T_3585;
    BITS #(.width(64), .high(5), .low(5)) bits_3772 (
        .y(_T_3585),
        .in(_T_3579)
    );
    wire _T_3586;
    BITS #(.width(64), .high(6), .low(6)) bits_3773 (
        .y(_T_3586),
        .in(_T_3579)
    );
    wire [1:0] _T_3587;
    BITS #(.width(64), .high(8), .low(7)) bits_3774 (
        .y(_T_3587),
        .in(_T_3579)
    );
    wire [1:0] _T_3588;
    BITS #(.width(64), .high(10), .low(9)) bits_3775 (
        .y(_T_3588),
        .in(_T_3579)
    );
    wire _T_3589;
    BITS #(.width(64), .high(11), .low(11)) bits_3776 (
        .y(_T_3589),
        .in(_T_3579)
    );
    wire _T_3590;
    BITS #(.width(64), .high(12), .low(12)) bits_3777 (
        .y(_T_3590),
        .in(_T_3579)
    );
    wire [39:0] _T_3591;
    BITS #(.width(64), .high(52), .low(13)) bits_3778 (
        .y(_T_3591),
        .in(_T_3579)
    );
    wire [5:0] _T_3592;
    BITS #(.width(64), .high(58), .low(53)) bits_3779 (
        .y(_T_3592),
        .in(_T_3579)
    );
    wire _T_3593;
    BITS #(.width(64), .high(59), .low(59)) bits_3780 (
        .y(_T_3593),
        .in(_T_3579)
    );
    wire [3:0] _T_3594;
    BITS #(.width(64), .high(63), .low(60)) bits_3781 (
        .y(_T_3594),
        .in(_T_3579)
    );
    assign _T_1382_debug = io_status_debug;
    assign _T_1382_fs = io_status_fs;
    assign _T_1382_hie = 1'h0;
    assign _T_1382_hpie = 1'h0;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_3782 (
        .y(_T_1382_hpp),
        .in(1'h0)
    );
    assign _T_1382_isa = io_status_isa;
    assign _T_1382_mie = 1'h0;
    assign _T_1382_mpie = 1'h0;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_3783 (
        .y(_T_1382_mpp),
        .in(1'h0)
    );
    assign _T_1382_mprv = 1'h0;
    assign _T_1382_mxr = io_status_mxr;
    assign _T_1382_prv = io_status_prv;
    assign _T_1382_pum = io_status_pum;
    assign _T_1382_sd = io_status_sd;
    assign _T_1382_sd_rv32 = io_status_sd_rv32;
    assign _T_1382_sie = io_status_sie;
    assign _T_1382_spie = io_status_spie;
    assign _T_1382_spp = io_status_spp;
    assign _T_1382_sxl = io_status_sxl;
    assign _T_1382_tsr = io_status_tsr;
    assign _T_1382_tvm = io_status_tvm;
    assign _T_1382_tw = io_status_tw;
    assign _T_1382_uie = io_status_uie;
    assign _T_1382_upie = io_status_upie;
    assign _T_1382_uxl = io_status_uxl;
    assign _T_1382_xs = io_status_xs;
    assign _T_1382_zero1 = io_status_zero1;
    assign _T_1382_zero2 = io_status_zero2;
    assign _T_2861 = _T_2859;
    assign _T_2929_debug = _node_121;
    assign _T_2929_fs = _node_122;
    assign _T_2929_hie = _node_123;
    assign _T_2929_hpie = _node_124;
    assign _T_2929_hpp = _node_125;
    assign _T_2929_isa = _node_126;
    assign _T_2929_mie = _node_127;
    assign _T_2929_mpie = _node_128;
    assign _T_2929_mpp = _node_129;
    assign _T_2929_mprv = _node_130;
    assign _T_2929_mxr = _node_131;
    assign _T_2929_prv = _node_132;
    assign _T_2929_pum = _node_133;
    assign _T_2929_sd = _node_134;
    assign _T_2929_sd_rv32 = _node_135;
    assign _T_2929_sie = _node_136;
    assign _T_2929_spie = _node_137;
    assign _T_2929_spp = _node_138;
    assign _T_2929_sxl = _node_139;
    assign _T_2929_tsr = _node_140;
    assign _T_2929_tvm = _node_141;
    assign _T_2929_tw = _node_142;
    assign _T_2929_uie = _node_143;
    assign _T_2929_upie = _node_144;
    assign _T_2929_uxl = _node_145;
    assign _T_2929_xs = _node_146;
    assign _T_2929_zero1 = _node_147;
    assign _T_2929_zero2 = _node_148;
    PAD_UNSIGNED #(.width(64), .n(99)) u_pad_3784 (
        .y(_T_2959),
        .in(_node_149)
    );
    assign _T_3034_heip = _node_150;
    assign _T_3034_hsip = _node_151;
    assign _T_3034_htip = _node_152;
    assign _T_3034_meip = _node_153;
    assign _T_3034_msip = _node_154;
    assign _T_3034_mtip = _node_155;
    assign _T_3034_rocc = _node_156;
    assign _T_3034_seip = _node_157;
    assign _T_3034_ssip = _node_158;
    assign _T_3034_stip = _node_159;
    assign _T_3034_ueip = _node_160;
    assign _T_3034_usip = _node_161;
    assign _T_3034_utip = _node_162;
    BITS #(.width(64), .high(12), .low(0)) bits_3785 (
        .y(_T_3049),
        .in(_node_163)
    );
    assign _T_3118_cause = _node_164;
    assign _T_3118_debugint = _node_165;
    assign _T_3118_ebreakh = _node_166;
    assign _T_3118_ebreakm = _node_167;
    assign _T_3118_ebreaks = _node_168;
    assign _T_3118_ebreaku = _node_169;
    assign _T_3118_fullreset = _node_170;
    assign _T_3118_halt = _node_171;
    assign _T_3118_ndreset = _node_172;
    assign _T_3118_prv = _node_173;
    assign _T_3118_step = _node_174;
    assign _T_3118_stopcycle = _node_175;
    assign _T_3118_stoptime = _node_176;
    assign _T_3118_xdebugver = _node_177;
    assign _T_3118_zero1 = _node_178;
    assign _T_3118_zero2 = _node_179;
    assign _T_3118_zero3 = _node_180;
    BITS #(.width(64), .high(31), .low(0)) bits_3786 (
        .y(_T_3137),
        .in(_node_181)
    );
    assign _T_3217_debug = _node_182;
    assign _T_3217_fs = _node_183;
    assign _T_3217_hie = _node_184;
    assign _T_3217_hpie = _node_185;
    assign _T_3217_hpp = _node_186;
    assign _T_3217_isa = _node_187;
    assign _T_3217_mie = _node_188;
    assign _T_3217_mpie = _node_189;
    assign _T_3217_mpp = _node_190;
    assign _T_3217_mprv = _node_191;
    assign _T_3217_mxr = _node_192;
    assign _T_3217_prv = _node_193;
    assign _T_3217_pum = _node_194;
    assign _T_3217_sd = _node_195;
    assign _T_3217_sd_rv32 = _node_196;
    assign _T_3217_sie = _node_197;
    assign _T_3217_spie = _node_198;
    assign _T_3217_spp = _node_199;
    assign _T_3217_sxl = _node_200;
    assign _T_3217_tsr = _node_201;
    assign _T_3217_tvm = _node_202;
    assign _T_3217_tw = _node_203;
    assign _T_3217_uie = _node_204;
    assign _T_3217_upie = _node_205;
    assign _T_3217_uxl = _node_206;
    assign _T_3217_xs = _node_207;
    assign _T_3217_zero1 = _node_208;
    assign _T_3217_zero2 = _node_209;
    PAD_UNSIGNED #(.width(64), .n(99)) u_pad_3787 (
        .y(_T_3247),
        .in(_node_210)
    );
    assign _T_3310_heip = _node_211;
    assign _T_3310_hsip = _node_212;
    assign _T_3310_htip = _node_213;
    assign _T_3310_meip = _node_214;
    assign _T_3310_msip = _node_215;
    assign _T_3310_mtip = _node_216;
    assign _T_3310_rocc = _node_217;
    assign _T_3310_seip = _node_218;
    assign _T_3310_ssip = _node_219;
    assign _T_3310_stip = _node_220;
    assign _T_3310_ueip = _node_221;
    assign _T_3310_usip = _node_222;
    assign _T_3310_utip = _node_223;
    BITS #(.width(64), .high(12), .low(0)) bits_3788 (
        .y(_T_3325),
        .in(_node_224)
    );
    assign _T_3347_asid = _node_225;
    assign _T_3347_mode = _node_226;
    assign _T_3347_ppn = _node_227;
    assign _T_3352 = _node_228;
    assign _T_3461_action = _node_229;
    assign _T_3461_chain = _node_230;
    assign _T_3461_dmode = _node_231;
    assign _T_3461_h = _node_232;
    assign _T_3461_m = _node_233;
    assign _T_3461_maskmax = _node_234;
    assign _T_3461_r = _node_235;
    assign _T_3461_reserved = _node_236;
    assign _T_3461_s = _node_237;
    assign _T_3461_tmatch = _node_238;
    assign _T_3461_ttype = _node_239;
    assign _T_3461_u = _node_240;
    assign _T_3461_w = _node_241;
    assign _T_3461_x = _node_242;
    assign _T_3461_zero = _node_243;
    assign _T_347_debug = _T_405;
    assign _T_347_fs = _T_389;
    assign _T_347_hie = _T_380;
    assign _T_347_hpie = _T_384;
    assign _T_347_hpp = _T_387;
    assign _T_347_isa = _T_404;
    assign _T_347_mie = _T_381;
    assign _T_347_mpie = _T_385;
    assign _T_347_mpp = _T_388;
    assign _T_347_mprv = _T_391;
    assign _T_347_mxr = _T_393;
    assign _T_347_prv = _T_403;
    assign _T_347_pum = _T_392;
    assign _T_347_sd = _T_402;
    assign _T_347_sd_rv32 = _T_398;
    assign _T_347_sie = _T_379;
    assign _T_347_spie = _T_383;
    assign _T_347_spp = _T_386;
    assign _T_347_sxl = _T_400;
    assign _T_347_tsr = _T_396;
    assign _T_347_tvm = _T_394;
    assign _T_347_tw = _T_395;
    assign _T_347_uie = _T_378;
    assign _T_347_upie = _T_382;
    assign _T_347_uxl = _T_399;
    assign _T_347_xs = _T_390;
    assign _T_347_zero1 = _T_397;
    assign _T_347_zero2 = _T_401;
    assign _T_3478 = _node_244;
    assign _T_3556_address = _T_3576;
    assign _T_3556_control_action = _T_3590;
    assign _T_3556_control_chain = _T_3589;
    assign _T_3556_control_dmode = _T_3593;
    assign _T_3556_control_h = _T_3585;
    assign _T_3556_control_m = _T_3586;
    assign _T_3556_control_maskmax = _T_3592;
    assign _T_3556_control_r = _T_3580;
    assign _T_3556_control_reserved = _T_3591;
    assign _T_3556_control_s = _T_3584;
    assign _T_3556_control_tmatch = _T_3587;
    assign _T_3556_control_ttype = _T_3594;
    assign _T_3556_control_u = _T_3583;
    assign _T_3556_control_w = _T_3581;
    assign _T_3556_control_x = _T_3582;
    assign _T_3556_control_zero = _T_3588;
    PAD_UNSIGNED #(.width(1), .n(103)) u_pad_3789 (
        .y(_T_3575),
        .in(1'h0)
    );
    assign _T_3579 = _T_3577;
    PAD_UNSIGNED #(.width(1), .n(99)) u_pad_3790 (
        .y(_T_377),
        .in(1'h0)
    );
    assign _T_505_cause = _T_530;
    assign _T_505_debugint = _T_529;
    assign _T_505_ebreakh = _T_536;
    assign _T_505_ebreakm = _T_537;
    assign _T_505_ebreaks = _T_535;
    assign _T_505_ebreaku = _T_534;
    assign _T_505_fullreset = _T_539;
    assign _T_505_halt = _T_527;
    assign _T_505_ndreset = _T_540;
    assign _T_505_prv = _T_525;
    assign _T_505_step = _T_526;
    assign _T_505_stopcycle = _T_532;
    assign _T_505_stoptime = _T_531;
    assign _T_505_xdebugver = _T_541;
    assign _T_505_zero1 = _T_528;
    assign _T_505_zero2 = _T_533;
    assign _T_505_zero3 = _T_538;
    PAD_UNSIGNED #(.width(1), .n(32)) u_pad_3791 (
        .y(_T_524),
        .in(1'h0)
    );
    assign _T_607_heip = _T_633;
    assign _T_607_hsip = _T_625;
    assign _T_607_htip = _T_629;
    assign _T_607_meip = _T_634;
    assign _T_607_msip = _T_626;
    assign _T_607_mtip = _T_630;
    assign _T_607_rocc = _T_635;
    assign _T_607_seip = _T_632;
    assign _T_607_ssip = _T_624;
    assign _T_607_stip = _T_628;
    assign _T_607_ueip = _T_631;
    assign _T_607_usip = _T_623;
    assign _T_607_utip = _T_627;
    PAD_UNSIGNED #(.width(1), .n(13)) u_pad_3792 (
        .y(_T_622),
        .in(1'h0)
    );
    assign _T_636_heip = _T_607_heip;
    assign _T_636_hsip = _T_607_hsip;
    assign _T_636_htip = _T_607_htip;
    assign _T_636_meip = 1'h1;
    assign _T_636_msip = 1'h1;
    assign _T_636_mtip = 1'h1;
    assign _T_636_rocc = 1'h0;
    assign _T_636_seip = 1'h1;
    assign _T_636_ssip = 1'h1;
    assign _T_636_stip = 1'h1;
    assign _T_636_ueip = _T_607_ueip;
    assign _T_636_usip = _T_607_usip;
    assign _T_636_utip = _T_607_utip;
    assign _T_657_heip = _T_636_heip;
    assign _T_657_hsip = _T_636_hsip;
    assign _T_657_htip = _T_636_htip;
    assign _T_657_meip = 1'h0;
    assign _T_657_msip = 1'h0;
    assign _T_657_mtip = 1'h0;
    assign _T_657_rocc = _T_636_rocc;
    assign _T_657_seip = _T_636_seip;
    assign _T_657_ssip = _T_636_ssip;
    assign _T_657_stip = _T_636_stip;
    assign _T_657_ueip = _T_636_ueip;
    assign _T_657_usip = _T_636_usip;
    assign _T_657_utip = _T_636_utip;
    wire [63:0] _WTEMP_538;
    wire [63:0] _WTEMP_539;
    PAD_UNSIGNED #(.width(7), .n(64)) u_pad_3793 (
        .y(_WTEMP_539),
        .in(_T_932)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_3794 (
        .y(_WTEMP_538),
        .sel(_T_2870),
        .a(_node_245),
        .b(_WTEMP_539)
    );
    BITS #(.width(64), .high(5), .low(0)) bits_3795 (
        .y(_WTEMP_144),
        .in(_WTEMP_538)
    );
    MUX_UNSIGNED #(.width(58)) u_mux_3796 (
        .y(_WTEMP_146),
        .sel(_T_2870),
        .a(_node_246),
        .b(_node_247)
    );
    wire [63:0] _WTEMP_540;
    wire [63:0] _WTEMP_541;
    PAD_UNSIGNED #(.width(7), .n(64)) u_pad_3797 (
        .y(_WTEMP_541),
        .in(_T_943)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_3798 (
        .y(_WTEMP_540),
        .sel(_T_2870),
        .a(_node_248),
        .b(_WTEMP_541)
    );
    BITS #(.width(64), .high(5), .low(0)) bits_3799 (
        .y(_WTEMP_148),
        .in(_WTEMP_540)
    );
    MUX_UNSIGNED #(.width(58)) u_mux_3800 (
        .y(_WTEMP_150),
        .sel(_T_2870),
        .a(_node_249),
        .b(_node_250)
    );
    assign io_bp_0_address = _reg_bp_0_address__q;
    assign io_bp_0_control_action = _reg_bp_0_control_action__q;
    assign io_bp_0_control_chain = 1'h0;
    assign io_bp_0_control_dmode = _reg_bp_0_control_dmode__q;
    assign io_bp_0_control_h = 1'h0;
    assign io_bp_0_control_m = _reg_bp_0_control_m__q;
    assign io_bp_0_control_maskmax = 6'h4;
    assign io_bp_0_control_r = _reg_bp_0_control_r__q;
    assign io_bp_0_control_reserved = 40'h0;
    assign io_bp_0_control_s = _reg_bp_0_control_s__q;
    assign io_bp_0_control_tmatch = _reg_bp_0_control_tmatch__q;
    assign io_bp_0_control_ttype = 4'h2;
    assign io_bp_0_control_u = _reg_bp_0_control_u__q;
    assign io_bp_0_control_w = _reg_bp_0_control_w__q;
    assign io_bp_0_control_x = _reg_bp_0_control_x__q;
    assign io_bp_0_control_zero = 2'h0;
    assign io_csr_stall = _reg_wfi__q;
    assign io_decode_fp_illegal = _T_1764;
    assign io_decode_read_illegal = _T_2203;
    assign io_decode_rocc_illegal = _T_1770;
    assign io_decode_system_illegal = _T_2245;
    assign io_decode_write_flush = _T_2220;
    assign io_decode_write_illegal = _T_2207;
    assign io_eret = _T_2331;
    MUX_UNSIGNED #(.width(40)) u_mux_3801 (
        .y(io_evec),
        .sel(insn_ret),
        .a(_node_49),
        .b(tvec)
    );
    assign io_fatc = insn_sfence_vma;
    assign io_fcsr_rm = _reg_frm__q;
    MUX_UNSIGNED #(.width(1)) u_mux_3802 (
        .y(io_interrupt),
        .sel(_T_1208),
        .a(1'h1),
        .b(_T_1203)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_3803 (
        .y(io_interrupt_cause),
        .sel(_T_1208),
        .a(64'h800000000000000D),
        .b(interruptCause)
    );
    assign io_ptbr_asid = 16'h0;
    assign io_ptbr_mode = _reg_sptbr_mode__q;
    assign io_ptbr_ppn = _reg_sptbr_ppn__q;
    assign io_rw_rdata = _T_2861;
    assign io_singleStep = _T_2334;
    assign io_status_debug = _reg_debug__q;
    assign io_status_fs = _reg_mstatus_fs__q;
    assign io_status_hie = 1'h0;
    assign io_status_hpie = 1'h0;
    assign io_status_hpp = 2'h0;
    BITS #(.width(64), .high(31), .low(0)) bits_3804 (
        .y(io_status_isa),
        .in(_reg_misa__q)
    );
    assign io_status_mie = _reg_mstatus_mie__q;
    assign io_status_mpie = _reg_mstatus_mpie__q;
    assign io_status_mpp = _reg_mstatus_mpp__q;
    assign io_status_mprv = _reg_mstatus_mprv__q;
    assign io_status_mxr = _reg_mstatus_mxr__q;
    assign io_status_prv = _reg_mstatus_prv__q;
    assign io_status_pum = _reg_mstatus_pum__q;
    assign io_status_sd = _T_2341;
    assign io_status_sd_rv32 = 1'h0;
    assign io_status_sie = _reg_mstatus_sie__q;
    assign io_status_spie = _reg_mstatus_spie__q;
    assign io_status_spp = _reg_mstatus_spp__q;
    assign io_status_sxl = 2'h2;
    assign io_status_tsr = _reg_mstatus_tsr__q;
    assign io_status_tvm = _reg_mstatus_tvm__q;
    assign io_status_tw = _reg_mstatus_tw__q;
    assign io_status_uie = 1'h0;
    assign io_status_upie = 1'h0;
    assign io_status_uxl = 2'h2;
    assign io_status_xs = 2'h0;
    assign io_status_zero1 = 8'h0;
    assign io_status_zero2 = 27'h0;
    assign io_time = _T_950;
    assign mip_heip = _reg_mip_heip__q;
    assign mip_hsip = _reg_mip_hsip__q;
    assign mip_htip = _reg_mip_htip__q;
    assign mip_meip = _reg_mip_meip__q;
    assign mip_msip = _reg_mip_msip__q;
    assign mip_mtip = _reg_mip_mtip__q;
    assign mip_rocc = io_rocc_interrupt;
    assign mip_seip = _reg_mip_seip__q;
    assign mip_ssip = _reg_mip_ssip__q;
    assign mip_stip = _reg_mip_stip__q;
    assign mip_ueip = _reg_mip_ueip__q;
    assign mip_usip = _reg_mip_usip__q;
    assign mip_utip = _reg_mip_utip__q;
    MUX_UNSIGNED #(.width(2)) u_mux_3805 (
        .y(new_prv),
        .sel(insn_ret),
        .a(_node_50),
        .b(_node_51)
    );
    wire [63:0] _WTEMP_542;
    BITS #(.width(64), .high(38), .low(0)) bits_3806 (
        .y(_reg_bp_0_address__d),
        .in(_WTEMP_542)
    );
    wire [63:0] _WTEMP_543;
    PAD_UNSIGNED #(.width(39), .n(64)) u_pad_3807 (
        .y(_WTEMP_543),
        .in(_reg_bp_0_address__q)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_3808 (
        .y(_WTEMP_542),
        .sel(_T_2870),
        .a(_node_251),
        .b(_WTEMP_543)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_3809 (
        .y(_reg_bp_0_control_action__d),
        .sel(reset),
        .a(1'h0),
        .b(_node_319)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_3810 (
        .y(_reg_bp_0_control_dmode__d),
        .sel(reset),
        .a(1'h0),
        .b(_node_320)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_3811 (
        .y(_reg_bp_0_control_m__d),
        .sel(_T_2870),
        .a(_node_254),
        .b(_reg_bp_0_control_m__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_3812 (
        .y(_reg_bp_0_control_r__d),
        .sel(reset),
        .a(1'h0),
        .b(_node_321)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_3813 (
        .y(_reg_bp_0_control_s__d),
        .sel(_T_2870),
        .a(_node_256),
        .b(_reg_bp_0_control_s__q)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_3814 (
        .y(_reg_bp_0_control_tmatch__d),
        .sel(_T_2870),
        .a(_node_257),
        .b(_reg_bp_0_control_tmatch__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_3815 (
        .y(_reg_bp_0_control_u__d),
        .sel(_T_2870),
        .a(_node_258),
        .b(_reg_bp_0_control_u__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_3816 (
        .y(_reg_bp_0_control_w__d),
        .sel(reset),
        .a(1'h0),
        .b(_node_322)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_3817 (
        .y(_reg_bp_0_control_x__d),
        .sel(reset),
        .a(1'h0),
        .b(_node_323)
    );
    assign _reg_bp_1_address__d = _T_3556_address;
    assign _reg_bp_1_control_action__d = _T_3556_control_action;
    assign _reg_bp_1_control_dmode__d = _T_3556_control_dmode;
    assign _reg_bp_1_control_m__d = _T_3556_control_m;
    assign _reg_bp_1_control_r__d = _T_3556_control_r;
    assign _reg_bp_1_control_s__d = _T_3556_control_s;
    assign _reg_bp_1_control_tmatch__d = _T_3556_control_tmatch;
    assign _reg_bp_1_control_u__d = _T_3556_control_u;
    assign _reg_bp_1_control_w__d = _T_3556_control_w;
    assign _reg_bp_1_control_x__d = _T_3556_control_x;
    MUX_UNSIGNED #(.width(3)) u_mux_3818 (
        .y(_WTEMP_136),
        .sel(exception),
        .a(_node_14),
        .b(_reg_dcsr_cause__q)
    );
    assign _WTEMP_137 = io_interrupts_debug;
    MUX_UNSIGNED #(.width(1)) u_mux_3819 (
        .y(_WTEMP_133),
        .sel(_T_2870),
        .a(_node_261),
        .b(_reg_dcsr_ebreakm__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_3820 (
        .y(_WTEMP_134),
        .sel(_T_2870),
        .a(_node_262),
        .b(_reg_dcsr_ebreaks__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_3821 (
        .y(_WTEMP_135),
        .sel(_T_2870),
        .a(_node_263),
        .b(_reg_dcsr_ebreaku__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_3822 (
        .y(_WTEMP_138),
        .sel(_T_2870),
        .a(_node_264),
        .b(_reg_dcsr_halt__q)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_3823 (
        .y(_WTEMP_140),
        .sel(_T_2870),
        .a(_node_265),
        .b(_node_266)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_3824 (
        .y(_WTEMP_139),
        .sel(_T_2870),
        .a(_node_267),
        .b(_reg_dcsr_step__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_3825 (
        .y(_WTEMP_141),
        .sel(insn_ret),
        .a(_node_52),
        .b(_node_53)
    );
    wire [63:0] _WTEMP_544;
    BITS #(.width(64), .high(39), .low(0)) bits_3826 (
        .y(_reg_dpc__d),
        .in(_WTEMP_544)
    );
    wire [63:0] _WTEMP_545;
    PAD_UNSIGNED #(.width(40), .n(64)) u_pad_3827 (
        .y(_WTEMP_545),
        .in(_node_269)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_3828 (
        .y(_WTEMP_544),
        .sel(_T_2870),
        .a(_node_268),
        .b(_WTEMP_545)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_3829 (
        .y(_reg_dscratch__d),
        .sel(_T_2870),
        .a(_node_270),
        .b(_reg_dscratch__q)
    );
    wire [63:0] _WTEMP_546;
    BITS #(.width(64), .high(4), .low(0)) bits_3830 (
        .y(_reg_fflags__d),
        .in(_WTEMP_546)
    );
    wire [63:0] _WTEMP_547;
    PAD_UNSIGNED #(.width(5), .n(64)) u_pad_3831 (
        .y(_WTEMP_547),
        .in(_node_272)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_3832 (
        .y(_WTEMP_546),
        .sel(_T_2870),
        .a(_node_271),
        .b(_WTEMP_547)
    );
    wire [63:0] _WTEMP_548;
    BITS #(.width(64), .high(2), .low(0)) bits_3833 (
        .y(_reg_frm__d),
        .in(_WTEMP_548)
    );
    wire [63:0] _WTEMP_549;
    PAD_UNSIGNED #(.width(3), .n(64)) u_pad_3834 (
        .y(_WTEMP_549),
        .in(_reg_frm__q)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_3835 (
        .y(_WTEMP_548),
        .sel(_T_2870),
        .a(_node_273),
        .b(_WTEMP_549)
    );
    MUX_UNSIGNED #(.width(40)) u_mux_3836 (
        .y(_reg_mbadaddr__d),
        .sel(_T_2870),
        .a(_node_274),
        .b(_node_275)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_3837 (
        .y(_reg_mcause__d),
        .sel(_T_2870),
        .a(_node_276),
        .b(_node_277)
    );
    wire [63:0] _WTEMP_550;
    BITS #(.width(64), .high(31), .low(0)) bits_3838 (
        .y(_reg_mcounteren__d),
        .in(_WTEMP_550)
    );
    wire [63:0] _WTEMP_551;
    PAD_UNSIGNED #(.width(32), .n(64)) u_pad_3839 (
        .y(_WTEMP_551),
        .in(_reg_mcounteren__q)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_3840 (
        .y(_WTEMP_550),
        .sel(_T_2870),
        .a(_node_278),
        .b(_WTEMP_551)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_3841 (
        .y(_reg_medeleg__d),
        .sel(_T_2870),
        .a(_node_279),
        .b(_reg_medeleg__q)
    );
    wire [63:0] _WTEMP_552;
    BITS #(.width(64), .high(39), .low(0)) bits_3842 (
        .y(_reg_mepc__d),
        .in(_WTEMP_552)
    );
    wire [63:0] _WTEMP_553;
    PAD_UNSIGNED #(.width(40), .n(64)) u_pad_3843 (
        .y(_WTEMP_553),
        .in(_node_281)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_3844 (
        .y(_WTEMP_552),
        .sel(_T_2870),
        .a(_node_280),
        .b(_WTEMP_553)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_3845 (
        .y(_reg_mideleg__d),
        .sel(_T_2870),
        .a(_node_282),
        .b(_reg_mideleg__q)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_3846 (
        .y(_reg_mie__d),
        .sel(_T_2870),
        .a(_node_283),
        .b(_reg_mie__q)
    );
    assign _reg_mip_meip__d = io_interrupts_meip;
    assign _reg_mip_msip__d = io_interrupts_msip;
    assign _reg_mip_mtip__d = io_interrupts_mtip;
    assign _reg_mip_seip__d = io_interrupts_seip;
    MUX_UNSIGNED #(.width(1)) u_mux_3847 (
        .y(_reg_mip_ssip__d),
        .sel(_T_2870),
        .a(_node_284),
        .b(_reg_mip_ssip__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_3848 (
        .y(_reg_mip_stip__d),
        .sel(_T_2870),
        .a(_node_285),
        .b(_reg_mip_stip__q)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_3849 (
        .y(_WTEMP_195),
        .sel(_T_2870),
        .a(_node_286),
        .b(_reg_misa__q)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_3850 (
        .y(_reg_mscratch__d),
        .sel(_T_2870),
        .a(_node_287),
        .b(_reg_mscratch__q)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_3851 (
        .y(_WTEMP_125),
        .sel(_T_2870),
        .a(_node_288),
        .b(_reg_mstatus_fs__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_3852 (
        .y(_WTEMP_130),
        .sel(_T_2870),
        .a(_node_289),
        .b(_node_290)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_3853 (
        .y(_WTEMP_128),
        .sel(_T_2870),
        .a(_node_291),
        .b(_node_292)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_3854 (
        .y(_WTEMP_126),
        .sel(_T_2870),
        .a(_node_293),
        .b(_node_294)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_3855 (
        .y(_WTEMP_124),
        .sel(_T_2870),
        .a(_node_295),
        .b(_reg_mstatus_mprv__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_3856 (
        .y(_WTEMP_122),
        .sel(_T_2870),
        .a(_node_296),
        .b(_reg_mstatus_mxr__q)
    );
    assign _WTEMP_118 = _T_467;
    MUX_UNSIGNED #(.width(1)) u_mux_3857 (
        .y(_WTEMP_123),
        .sel(_T_2870),
        .a(_node_297),
        .b(_reg_mstatus_pum__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_3858 (
        .y(_WTEMP_131),
        .sel(_T_2870),
        .a(_node_298),
        .b(_node_299)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_3859 (
        .y(_WTEMP_129),
        .sel(_T_2870),
        .a(_node_300),
        .b(_node_301)
    );
    wire [1:0] _WTEMP_554;
    MUX_UNSIGNED #(.width(2)) u_mux_3860 (
        .y(_WTEMP_554),
        .sel(_T_2870),
        .a(_node_302),
        .b(_node_303)
    );
    BITS #(.width(2), .high(0), .low(0)) bits_3861 (
        .y(_WTEMP_127),
        .in(_WTEMP_554)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_3862 (
        .y(_WTEMP_119),
        .sel(_T_2870),
        .a(_node_304),
        .b(_reg_mstatus_tsr__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_3863 (
        .y(_WTEMP_121),
        .sel(_T_2870),
        .a(_node_305),
        .b(_reg_mstatus_tvm__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_3864 (
        .y(_WTEMP_120),
        .sel(_T_2870),
        .a(_node_306),
        .b(_reg_mstatus_tw__q)
    );
    wire [63:0] _WTEMP_555;
    wire [63:0] _WTEMP_556;
    PAD_UNSIGNED #(.width(32), .n(64)) u_pad_3865 (
        .y(_WTEMP_556),
        .in(_reg_mtvec__q)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_3866 (
        .y(_WTEMP_555),
        .sel(_T_2870),
        .a(_node_307),
        .b(_WTEMP_556)
    );
    BITS #(.width(64), .high(31), .low(0)) bits_3867 (
        .y(_WTEMP_142),
        .in(_WTEMP_555)
    );
    MUX_UNSIGNED #(.width(40)) u_mux_3868 (
        .y(_reg_sbadaddr__d),
        .sel(_T_2870),
        .a(_node_308),
        .b(_node_309)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_3869 (
        .y(_reg_scause__d),
        .sel(_T_2870),
        .a(_node_310),
        .b(_node_311)
    );
    wire [63:0] _WTEMP_557;
    BITS #(.width(64), .high(31), .low(0)) bits_3870 (
        .y(_reg_scounteren__d),
        .in(_WTEMP_557)
    );
    wire [63:0] _WTEMP_558;
    PAD_UNSIGNED #(.width(32), .n(64)) u_pad_3871 (
        .y(_WTEMP_558),
        .in(_reg_scounteren__q)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_3872 (
        .y(_WTEMP_557),
        .sel(_T_2870),
        .a(_node_312),
        .b(_WTEMP_558)
    );
    wire [63:0] _WTEMP_559;
    BITS #(.width(64), .high(39), .low(0)) bits_3873 (
        .y(_reg_sepc__d),
        .in(_WTEMP_559)
    );
    wire [63:0] _WTEMP_560;
    PAD_UNSIGNED #(.width(40), .n(64)) u_pad_3874 (
        .y(_WTEMP_560),
        .in(_node_314)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_3875 (
        .y(_WTEMP_559),
        .sel(_T_2870),
        .a(_node_313),
        .b(_WTEMP_560)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_3876 (
        .y(_reg_singleStepped__d),
        .sel(_T_2369),
        .a(1'h0),
        .b(_node_9)
    );
    MUX_UNSIGNED #(.width(4)) u_mux_3877 (
        .y(_reg_sptbr_mode__d),
        .sel(_T_2870),
        .a(_node_315),
        .b(_reg_sptbr_mode__q)
    );
    MUX_UNSIGNED #(.width(44)) u_mux_3878 (
        .y(_reg_sptbr_ppn__d),
        .sel(_T_2870),
        .a(_node_316),
        .b(_reg_sptbr_ppn__q)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_3879 (
        .y(_reg_sscratch__d),
        .sel(_T_2870),
        .a(_node_317),
        .b(_reg_sscratch__q)
    );
    wire [63:0] _WTEMP_561;
    BITS #(.width(64), .high(38), .low(0)) bits_3880 (
        .y(_reg_stvec__d),
        .in(_WTEMP_561)
    );
    wire [63:0] _WTEMP_562;
    PAD_UNSIGNED #(.width(39), .n(64)) u_pad_3881 (
        .y(_WTEMP_562),
        .in(_reg_stvec__q)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_3882 (
        .y(_WTEMP_561),
        .sel(_T_2870),
        .a(_node_318),
        .b(_WTEMP_562)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_3883 (
        .y(_WTEMP_143),
        .sel(_T_2356),
        .a(1'h0),
        .b(_node_8)
    );
    assign reset_dcsr_cause = _T_505_cause;
    assign reset_dcsr_debugint = _T_505_debugint;
    assign reset_dcsr_ebreakm = _T_505_ebreakm;
    assign reset_dcsr_ebreaks = _T_505_ebreaks;
    assign reset_dcsr_ebreaku = _T_505_ebreaku;
    assign reset_dcsr_halt = _T_505_halt;
    assign reset_dcsr_prv = 2'h3;
    assign reset_dcsr_step = _T_505_step;
    assign reset_mstatus_fs = _T_347_fs;
    assign reset_mstatus_mie = _T_347_mie;
    assign reset_mstatus_mpie = _T_347_mpie;
    assign reset_mstatus_mpp = 2'h3;
    assign reset_mstatus_mprv = _T_347_mprv;
    assign reset_mstatus_mxr = _T_347_mxr;
    assign reset_mstatus_prv = 2'h3;
    assign reset_mstatus_pum = _T_347_pum;
    assign reset_mstatus_sie = _T_347_sie;
    assign reset_mstatus_spie = _T_347_spie;
    assign reset_mstatus_spp = _T_347_spp;
    assign reset_mstatus_tsr = _T_347_tsr;
    assign reset_mstatus_tvm = _T_347_tvm;
    assign reset_mstatus_tw = _T_347_tw;
endmodule //CSRFile
module LEQ_UNSIGNED(y, a, b);
    parameter width = 4;
    output y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a <= b;
endmodule // LEQ_UNSIGNED
module BreakpointUnit(
    input clock,
    input reset,
    input io_status_debug,
    input [31:0] io_status_isa,
    input [1:0] io_status_prv,
    input io_status_sd,
    input [26:0] io_status_zero2,
    input [1:0] io_status_sxl,
    input [1:0] io_status_uxl,
    input io_status_sd_rv32,
    input [7:0] io_status_zero1,
    input io_status_tsr,
    input io_status_tw,
    input io_status_tvm,
    input io_status_mxr,
    input io_status_pum,
    input io_status_mprv,
    input [1:0] io_status_xs,
    input [1:0] io_status_fs,
    input [1:0] io_status_mpp,
    input [1:0] io_status_hpp,
    input io_status_spp,
    input io_status_mpie,
    input io_status_hpie,
    input io_status_spie,
    input io_status_upie,
    input io_status_mie,
    input io_status_hie,
    input io_status_sie,
    input io_status_uie,
    input [3:0] io_bp_0_control_ttype,
    input io_bp_0_control_dmode,
    input [5:0] io_bp_0_control_maskmax,
    input [39:0] io_bp_0_control_reserved,
    input io_bp_0_control_action,
    input io_bp_0_control_chain,
    input [1:0] io_bp_0_control_zero,
    input [1:0] io_bp_0_control_tmatch,
    input io_bp_0_control_m,
    input io_bp_0_control_h,
    input io_bp_0_control_s,
    input io_bp_0_control_u,
    input io_bp_0_control_x,
    input io_bp_0_control_w,
    input io_bp_0_control_r,
    input [38:0] io_bp_0_address,
    input [38:0] io_pc,
    input [38:0] io_ea,
    output io_xcpt_if,
    output io_xcpt_ld,
    output io_xcpt_st,
    output io_debug_if,
    output io_debug_ld,
    output io_debug_st
);
    wire _T_212;
    EQ_UNSIGNED #(.width(1)) u_eq_3948 (
        .y(_T_212),
        .a(io_status_debug),
        .b(1'h0)
    );
    wire [1:0] _T_213;
    CAT #(.width_a(1), .width_b(1)) cat_3949 (
        .y(_T_213),
        .a(io_bp_0_control_s),
        .b(io_bp_0_control_u)
    );
    wire [1:0] _T_214;
    CAT #(.width_a(1), .width_b(1)) cat_3950 (
        .y(_T_214),
        .a(io_bp_0_control_m),
        .b(io_bp_0_control_h)
    );
    wire [3:0] _T_215;
    CAT #(.width_a(2), .width_b(2)) cat_3951 (
        .y(_T_215),
        .a(_T_214),
        .b(_T_213)
    );
    wire [3:0] _T_216;
    DSHR_UNSIGNED #(.width_in(4), .width_n(2)) u_dshr_3952 (
        .y(_T_216),
        .in(_T_215),
        .n(io_status_prv)
    );
    wire _T_217;
    BITS #(.width(4), .high(0), .low(0)) bits_3953 (
        .y(_T_217),
        .in(_T_216)
    );
    wire _T_218;
    BITWISEAND #(.width(1)) bitwiseand_3954 (
        .y(_T_218),
        .a(_T_212),
        .b(_T_217)
    );
    wire _T_219;
    BITWISEAND #(.width(1)) bitwiseand_3955 (
        .y(_T_219),
        .a(_T_218),
        .b(1'h1)
    );
    wire _T_220;
    BITWISEAND #(.width(1)) bitwiseand_3956 (
        .y(_T_220),
        .a(_T_219),
        .b(io_bp_0_control_r)
    );
    wire _T_221;
    BITS #(.width(2), .high(1), .low(1)) bits_3957 (
        .y(_T_221),
        .in(io_bp_0_control_tmatch)
    );
    wire _T_222;
    GEQ_UNSIGNED #(.width(39)) u_geq_3958 (
        .y(_T_222),
        .a(io_ea),
        .b(io_bp_0_address)
    );
    wire _T_223;
    BITS #(.width(2), .high(0), .low(0)) bits_3959 (
        .y(_T_223),
        .in(io_bp_0_control_tmatch)
    );
    wire _T_224;
    BITWISEXOR #(.width(1)) bitwisexor_3960 (
        .y(_T_224),
        .a(_T_222),
        .b(_T_223)
    );
    wire [38:0] _T_225;
    BITWISENOT #(.width(39)) bitwisenot_3961 (
        .y(_T_225),
        .in(io_ea)
    );
    wire _T_226;
    BITS #(.width(2), .high(0), .low(0)) bits_3962 (
        .y(_T_226),
        .in(io_bp_0_control_tmatch)
    );
    wire _T_227;
    BITS #(.width(39), .high(0), .low(0)) bits_3963 (
        .y(_T_227),
        .in(io_bp_0_address)
    );
    wire _T_228;
    BITWISEAND #(.width(1)) bitwiseand_3964 (
        .y(_T_228),
        .a(_T_226),
        .b(_T_227)
    );
    wire _T_229;
    BITS #(.width(39), .high(1), .low(1)) bits_3965 (
        .y(_T_229),
        .in(io_bp_0_address)
    );
    wire _T_230;
    BITWISEAND #(.width(1)) bitwiseand_3966 (
        .y(_T_230),
        .a(_T_228),
        .b(_T_229)
    );
    wire _T_231;
    BITS #(.width(39), .high(2), .low(2)) bits_3967 (
        .y(_T_231),
        .in(io_bp_0_address)
    );
    wire _T_232;
    BITWISEAND #(.width(1)) bitwiseand_3968 (
        .y(_T_232),
        .a(_T_230),
        .b(_T_231)
    );
    wire [1:0] _T_233;
    CAT #(.width_a(1), .width_b(1)) cat_3969 (
        .y(_T_233),
        .a(_T_228),
        .b(_T_226)
    );
    wire [1:0] _T_234;
    CAT #(.width_a(1), .width_b(1)) cat_3970 (
        .y(_T_234),
        .a(_T_232),
        .b(_T_230)
    );
    wire [3:0] _T_235;
    CAT #(.width_a(2), .width_b(2)) cat_3971 (
        .y(_T_235),
        .a(_T_234),
        .b(_T_233)
    );
    wire [38:0] _T_236;
    wire [38:0] _WTEMP_564;
    PAD_UNSIGNED #(.width(4), .n(39)) u_pad_3972 (
        .y(_WTEMP_564),
        .in(_T_235)
    );
    BITWISEOR #(.width(39)) bitwiseor_3973 (
        .y(_T_236),
        .a(_T_225),
        .b(_WTEMP_564)
    );
    wire [38:0] _T_237;
    BITWISENOT #(.width(39)) bitwisenot_3974 (
        .y(_T_237),
        .in(io_bp_0_address)
    );
    wire _T_238;
    BITS #(.width(2), .high(0), .low(0)) bits_3975 (
        .y(_T_238),
        .in(io_bp_0_control_tmatch)
    );
    wire _T_239;
    BITS #(.width(39), .high(0), .low(0)) bits_3976 (
        .y(_T_239),
        .in(io_bp_0_address)
    );
    wire _T_240;
    BITWISEAND #(.width(1)) bitwiseand_3977 (
        .y(_T_240),
        .a(_T_238),
        .b(_T_239)
    );
    wire _T_241;
    BITS #(.width(39), .high(1), .low(1)) bits_3978 (
        .y(_T_241),
        .in(io_bp_0_address)
    );
    wire _T_242;
    BITWISEAND #(.width(1)) bitwiseand_3979 (
        .y(_T_242),
        .a(_T_240),
        .b(_T_241)
    );
    wire _T_243;
    BITS #(.width(39), .high(2), .low(2)) bits_3980 (
        .y(_T_243),
        .in(io_bp_0_address)
    );
    wire _T_244;
    BITWISEAND #(.width(1)) bitwiseand_3981 (
        .y(_T_244),
        .a(_T_242),
        .b(_T_243)
    );
    wire [1:0] _T_245;
    CAT #(.width_a(1), .width_b(1)) cat_3982 (
        .y(_T_245),
        .a(_T_240),
        .b(_T_238)
    );
    wire [1:0] _T_246;
    CAT #(.width_a(1), .width_b(1)) cat_3983 (
        .y(_T_246),
        .a(_T_244),
        .b(_T_242)
    );
    wire [3:0] _T_247;
    CAT #(.width_a(2), .width_b(2)) cat_3984 (
        .y(_T_247),
        .a(_T_246),
        .b(_T_245)
    );
    wire [38:0] _T_248;
    wire [38:0] _WTEMP_565;
    PAD_UNSIGNED #(.width(4), .n(39)) u_pad_3985 (
        .y(_WTEMP_565),
        .in(_T_247)
    );
    BITWISEOR #(.width(39)) bitwiseor_3986 (
        .y(_T_248),
        .a(_T_237),
        .b(_WTEMP_565)
    );
    wire _T_249;
    EQ_UNSIGNED #(.width(39)) u_eq_3987 (
        .y(_T_249),
        .a(_T_236),
        .b(_T_248)
    );
    wire _T_250;
    MUX_UNSIGNED #(.width(1)) u_mux_3988 (
        .y(_T_250),
        .sel(_T_221),
        .a(_T_224),
        .b(_T_249)
    );
    wire _T_251;
    BITWISEAND #(.width(1)) bitwiseand_3989 (
        .y(_T_251),
        .a(_T_220),
        .b(_T_250)
    );
    wire _T_252;
    BITWISEAND #(.width(1)) bitwiseand_3990 (
        .y(_T_252),
        .a(_T_218),
        .b(1'h1)
    );
    wire _T_253;
    BITWISEAND #(.width(1)) bitwiseand_3991 (
        .y(_T_253),
        .a(_T_252),
        .b(io_bp_0_control_w)
    );
    wire _T_254;
    BITS #(.width(2), .high(1), .low(1)) bits_3992 (
        .y(_T_254),
        .in(io_bp_0_control_tmatch)
    );
    wire _T_255;
    GEQ_UNSIGNED #(.width(39)) u_geq_3993 (
        .y(_T_255),
        .a(io_ea),
        .b(io_bp_0_address)
    );
    wire _T_256;
    BITS #(.width(2), .high(0), .low(0)) bits_3994 (
        .y(_T_256),
        .in(io_bp_0_control_tmatch)
    );
    wire _T_257;
    BITWISEXOR #(.width(1)) bitwisexor_3995 (
        .y(_T_257),
        .a(_T_255),
        .b(_T_256)
    );
    wire [38:0] _T_258;
    BITWISENOT #(.width(39)) bitwisenot_3996 (
        .y(_T_258),
        .in(io_ea)
    );
    wire _T_259;
    BITS #(.width(2), .high(0), .low(0)) bits_3997 (
        .y(_T_259),
        .in(io_bp_0_control_tmatch)
    );
    wire _T_260;
    BITS #(.width(39), .high(0), .low(0)) bits_3998 (
        .y(_T_260),
        .in(io_bp_0_address)
    );
    wire _T_261;
    BITWISEAND #(.width(1)) bitwiseand_3999 (
        .y(_T_261),
        .a(_T_259),
        .b(_T_260)
    );
    wire _T_262;
    BITS #(.width(39), .high(1), .low(1)) bits_4000 (
        .y(_T_262),
        .in(io_bp_0_address)
    );
    wire _T_263;
    BITWISEAND #(.width(1)) bitwiseand_4001 (
        .y(_T_263),
        .a(_T_261),
        .b(_T_262)
    );
    wire _T_264;
    BITS #(.width(39), .high(2), .low(2)) bits_4002 (
        .y(_T_264),
        .in(io_bp_0_address)
    );
    wire _T_265;
    BITWISEAND #(.width(1)) bitwiseand_4003 (
        .y(_T_265),
        .a(_T_263),
        .b(_T_264)
    );
    wire [1:0] _T_266;
    CAT #(.width_a(1), .width_b(1)) cat_4004 (
        .y(_T_266),
        .a(_T_261),
        .b(_T_259)
    );
    wire [1:0] _T_267;
    CAT #(.width_a(1), .width_b(1)) cat_4005 (
        .y(_T_267),
        .a(_T_265),
        .b(_T_263)
    );
    wire [3:0] _T_268;
    CAT #(.width_a(2), .width_b(2)) cat_4006 (
        .y(_T_268),
        .a(_T_267),
        .b(_T_266)
    );
    wire [38:0] _T_269;
    wire [38:0] _WTEMP_566;
    PAD_UNSIGNED #(.width(4), .n(39)) u_pad_4007 (
        .y(_WTEMP_566),
        .in(_T_268)
    );
    BITWISEOR #(.width(39)) bitwiseor_4008 (
        .y(_T_269),
        .a(_T_258),
        .b(_WTEMP_566)
    );
    wire [38:0] _T_270;
    BITWISENOT #(.width(39)) bitwisenot_4009 (
        .y(_T_270),
        .in(io_bp_0_address)
    );
    wire _T_271;
    BITS #(.width(2), .high(0), .low(0)) bits_4010 (
        .y(_T_271),
        .in(io_bp_0_control_tmatch)
    );
    wire _T_272;
    BITS #(.width(39), .high(0), .low(0)) bits_4011 (
        .y(_T_272),
        .in(io_bp_0_address)
    );
    wire _T_273;
    BITWISEAND #(.width(1)) bitwiseand_4012 (
        .y(_T_273),
        .a(_T_271),
        .b(_T_272)
    );
    wire _T_274;
    BITS #(.width(39), .high(1), .low(1)) bits_4013 (
        .y(_T_274),
        .in(io_bp_0_address)
    );
    wire _T_275;
    BITWISEAND #(.width(1)) bitwiseand_4014 (
        .y(_T_275),
        .a(_T_273),
        .b(_T_274)
    );
    wire _T_276;
    BITS #(.width(39), .high(2), .low(2)) bits_4015 (
        .y(_T_276),
        .in(io_bp_0_address)
    );
    wire _T_277;
    BITWISEAND #(.width(1)) bitwiseand_4016 (
        .y(_T_277),
        .a(_T_275),
        .b(_T_276)
    );
    wire [1:0] _T_278;
    CAT #(.width_a(1), .width_b(1)) cat_4017 (
        .y(_T_278),
        .a(_T_273),
        .b(_T_271)
    );
    wire [1:0] _T_279;
    CAT #(.width_a(1), .width_b(1)) cat_4018 (
        .y(_T_279),
        .a(_T_277),
        .b(_T_275)
    );
    wire [3:0] _T_280;
    CAT #(.width_a(2), .width_b(2)) cat_4019 (
        .y(_T_280),
        .a(_T_279),
        .b(_T_278)
    );
    wire [38:0] _T_281;
    wire [38:0] _WTEMP_567;
    PAD_UNSIGNED #(.width(4), .n(39)) u_pad_4020 (
        .y(_WTEMP_567),
        .in(_T_280)
    );
    BITWISEOR #(.width(39)) bitwiseor_4021 (
        .y(_T_281),
        .a(_T_270),
        .b(_WTEMP_567)
    );
    wire _T_282;
    EQ_UNSIGNED #(.width(39)) u_eq_4022 (
        .y(_T_282),
        .a(_T_269),
        .b(_T_281)
    );
    wire _T_283;
    MUX_UNSIGNED #(.width(1)) u_mux_4023 (
        .y(_T_283),
        .sel(_T_254),
        .a(_T_257),
        .b(_T_282)
    );
    wire _T_284;
    BITWISEAND #(.width(1)) bitwiseand_4024 (
        .y(_T_284),
        .a(_T_253),
        .b(_T_283)
    );
    wire _T_285;
    BITWISEAND #(.width(1)) bitwiseand_4025 (
        .y(_T_285),
        .a(_T_218),
        .b(1'h1)
    );
    wire _T_286;
    BITWISEAND #(.width(1)) bitwiseand_4026 (
        .y(_T_286),
        .a(_T_285),
        .b(io_bp_0_control_x)
    );
    wire _T_287;
    BITS #(.width(2), .high(1), .low(1)) bits_4027 (
        .y(_T_287),
        .in(io_bp_0_control_tmatch)
    );
    wire _T_288;
    GEQ_UNSIGNED #(.width(39)) u_geq_4028 (
        .y(_T_288),
        .a(io_pc),
        .b(io_bp_0_address)
    );
    wire _T_289;
    BITS #(.width(2), .high(0), .low(0)) bits_4029 (
        .y(_T_289),
        .in(io_bp_0_control_tmatch)
    );
    wire _T_290;
    BITWISEXOR #(.width(1)) bitwisexor_4030 (
        .y(_T_290),
        .a(_T_288),
        .b(_T_289)
    );
    wire [38:0] _T_291;
    BITWISENOT #(.width(39)) bitwisenot_4031 (
        .y(_T_291),
        .in(io_pc)
    );
    wire _T_292;
    BITS #(.width(2), .high(0), .low(0)) bits_4032 (
        .y(_T_292),
        .in(io_bp_0_control_tmatch)
    );
    wire _T_293;
    BITS #(.width(39), .high(0), .low(0)) bits_4033 (
        .y(_T_293),
        .in(io_bp_0_address)
    );
    wire _T_294;
    BITWISEAND #(.width(1)) bitwiseand_4034 (
        .y(_T_294),
        .a(_T_292),
        .b(_T_293)
    );
    wire _T_295;
    BITS #(.width(39), .high(1), .low(1)) bits_4035 (
        .y(_T_295),
        .in(io_bp_0_address)
    );
    wire _T_296;
    BITWISEAND #(.width(1)) bitwiseand_4036 (
        .y(_T_296),
        .a(_T_294),
        .b(_T_295)
    );
    wire _T_297;
    BITS #(.width(39), .high(2), .low(2)) bits_4037 (
        .y(_T_297),
        .in(io_bp_0_address)
    );
    wire _T_298;
    BITWISEAND #(.width(1)) bitwiseand_4038 (
        .y(_T_298),
        .a(_T_296),
        .b(_T_297)
    );
    wire [1:0] _T_299;
    CAT #(.width_a(1), .width_b(1)) cat_4039 (
        .y(_T_299),
        .a(_T_294),
        .b(_T_292)
    );
    wire [1:0] _T_300;
    CAT #(.width_a(1), .width_b(1)) cat_4040 (
        .y(_T_300),
        .a(_T_298),
        .b(_T_296)
    );
    wire [3:0] _T_301;
    CAT #(.width_a(2), .width_b(2)) cat_4041 (
        .y(_T_301),
        .a(_T_300),
        .b(_T_299)
    );
    wire [38:0] _T_302;
    wire [38:0] _WTEMP_568;
    PAD_UNSIGNED #(.width(4), .n(39)) u_pad_4042 (
        .y(_WTEMP_568),
        .in(_T_301)
    );
    BITWISEOR #(.width(39)) bitwiseor_4043 (
        .y(_T_302),
        .a(_T_291),
        .b(_WTEMP_568)
    );
    wire [38:0] _T_303;
    BITWISENOT #(.width(39)) bitwisenot_4044 (
        .y(_T_303),
        .in(io_bp_0_address)
    );
    wire _T_304;
    BITS #(.width(2), .high(0), .low(0)) bits_4045 (
        .y(_T_304),
        .in(io_bp_0_control_tmatch)
    );
    wire _T_305;
    BITS #(.width(39), .high(0), .low(0)) bits_4046 (
        .y(_T_305),
        .in(io_bp_0_address)
    );
    wire _T_306;
    BITWISEAND #(.width(1)) bitwiseand_4047 (
        .y(_T_306),
        .a(_T_304),
        .b(_T_305)
    );
    wire _T_307;
    BITS #(.width(39), .high(1), .low(1)) bits_4048 (
        .y(_T_307),
        .in(io_bp_0_address)
    );
    wire _T_308;
    BITWISEAND #(.width(1)) bitwiseand_4049 (
        .y(_T_308),
        .a(_T_306),
        .b(_T_307)
    );
    wire _T_309;
    BITS #(.width(39), .high(2), .low(2)) bits_4050 (
        .y(_T_309),
        .in(io_bp_0_address)
    );
    wire _T_310;
    BITWISEAND #(.width(1)) bitwiseand_4051 (
        .y(_T_310),
        .a(_T_308),
        .b(_T_309)
    );
    wire [1:0] _T_311;
    CAT #(.width_a(1), .width_b(1)) cat_4052 (
        .y(_T_311),
        .a(_T_306),
        .b(_T_304)
    );
    wire [1:0] _T_312;
    CAT #(.width_a(1), .width_b(1)) cat_4053 (
        .y(_T_312),
        .a(_T_310),
        .b(_T_308)
    );
    wire [3:0] _T_313;
    CAT #(.width_a(2), .width_b(2)) cat_4054 (
        .y(_T_313),
        .a(_T_312),
        .b(_T_311)
    );
    wire [38:0] _T_314;
    wire [38:0] _WTEMP_569;
    PAD_UNSIGNED #(.width(4), .n(39)) u_pad_4055 (
        .y(_WTEMP_569),
        .in(_T_313)
    );
    BITWISEOR #(.width(39)) bitwiseor_4056 (
        .y(_T_314),
        .a(_T_303),
        .b(_WTEMP_569)
    );
    wire _T_315;
    EQ_UNSIGNED #(.width(39)) u_eq_4057 (
        .y(_T_315),
        .a(_T_302),
        .b(_T_314)
    );
    wire _T_316;
    MUX_UNSIGNED #(.width(1)) u_mux_4058 (
        .y(_T_316),
        .sel(_T_287),
        .a(_T_290),
        .b(_T_315)
    );
    wire _T_317;
    BITWISEAND #(.width(1)) bitwiseand_4059 (
        .y(_T_317),
        .a(_T_286),
        .b(_T_316)
    );
    wire _T_319;
    EQ_UNSIGNED #(.width(1)) u_eq_4060 (
        .y(_T_319),
        .a(io_bp_0_control_chain),
        .b(1'h0)
    );
    wire _T_320;
    BITWISEAND #(.width(1)) bitwiseand_4061 (
        .y(_T_320),
        .a(_T_319),
        .b(_T_251)
    );
    wire _T_322;
    EQ_UNSIGNED #(.width(1)) u_eq_4062 (
        .y(_T_322),
        .a(io_bp_0_control_action),
        .b(1'h0)
    );
    wire _T_323;
    BITWISEAND #(.width(1)) bitwiseand_4063 (
        .y(_T_323),
        .a(_T_319),
        .b(_T_284)
    );
    wire _T_325;
    EQ_UNSIGNED #(.width(1)) u_eq_4064 (
        .y(_T_325),
        .a(io_bp_0_control_action),
        .b(1'h0)
    );
    wire _T_326;
    BITWISEAND #(.width(1)) bitwiseand_4065 (
        .y(_T_326),
        .a(_T_319),
        .b(_T_317)
    );
    wire _T_328;
    EQ_UNSIGNED #(.width(1)) u_eq_4066 (
        .y(_T_328),
        .a(io_bp_0_control_action),
        .b(1'h0)
    );
    wire _T_329;
    BITWISEOR #(.width(1)) bitwiseor_4067 (
        .y(_T_329),
        .a(_T_319),
        .b(_T_251)
    );
    wire _T_330;
    BITWISEOR #(.width(1)) bitwiseor_4068 (
        .y(_T_330),
        .a(_T_319),
        .b(_T_284)
    );
    wire _T_331;
    BITWISEOR #(.width(1)) bitwiseor_4069 (
        .y(_T_331),
        .a(_T_319),
        .b(_T_317)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_4070 (
        .y(io_debug_if),
        .sel(_T_326),
        .a(io_bp_0_control_action),
        .b(1'h0)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_4071 (
        .y(io_debug_ld),
        .sel(_T_320),
        .a(io_bp_0_control_action),
        .b(1'h0)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_4072 (
        .y(io_debug_st),
        .sel(_T_323),
        .a(io_bp_0_control_action),
        .b(1'h0)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_4073 (
        .y(io_xcpt_if),
        .sel(_T_326),
        .a(_T_328),
        .b(1'h0)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_4074 (
        .y(io_xcpt_ld),
        .sel(_T_320),
        .a(_T_322),
        .b(1'h0)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_4075 (
        .y(io_xcpt_st),
        .sel(_T_323),
        .a(_T_325),
        .b(1'h0)
    );
endmodule //BreakpointUnit
module BITWISEXOR(y, a, b);
    parameter width = 4;
    output [width-1:0] y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a ^ b;
endmodule // BITWISEXOR
module MUX_SIGNED(y, sel, a, b);
    parameter width = 4;
    output [width-1:0] y;
    input sel;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = sel ? $signed(a) : $signed(b);
endmodule // MUX_SIGNED
module ALU(
    input clock,
    input reset,
    input io_dw,
    input [3:0] io_fn,
    input [63:0] io_in2,
    input [63:0] io_in1,
    output [63:0] io_out,
    output [63:0] io_adder_out,
    output io_cmp_out
);
    wire _T_16;
    BITS #(.width(4), .high(3), .low(3)) bits_4218 (
        .y(_T_16),
        .in(io_fn)
    );
    wire [63:0] _T_17;
    BITWISENOT #(.width(64)) bitwisenot_4219 (
        .y(_T_17),
        .in(io_in2)
    );
    wire [63:0] in2_inv;
    MUX_UNSIGNED #(.width(64)) u_mux_4220 (
        .y(in2_inv),
        .sel(_T_16),
        .a(_T_17),
        .b(io_in2)
    );
    wire [63:0] in1_xor_in2;
    BITWISEXOR #(.width(64)) bitwisexor_4221 (
        .y(in1_xor_in2),
        .a(io_in1),
        .b(in2_inv)
    );
    wire [64:0] _T_18;
    ADD_UNSIGNED #(.width(64)) u_add_4222 (
        .y(_T_18),
        .a(io_in1),
        .b(in2_inv)
    );
    wire [63:0] _T_19;
    TAIL #(.width(65), .n(1)) tail_4223 (
        .y(_T_19),
        .in(_T_18)
    );
    wire _T_20;
    BITS #(.width(4), .high(3), .low(3)) bits_4224 (
        .y(_T_20),
        .in(io_fn)
    );
    wire [64:0] _T_21;
    wire [63:0] _WTEMP_585;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_4225 (
        .y(_WTEMP_585),
        .in(_T_20)
    );
    ADD_UNSIGNED #(.width(64)) u_add_4226 (
        .y(_T_21),
        .a(_T_19),
        .b(_WTEMP_585)
    );
    wire [63:0] _T_22;
    TAIL #(.width(65), .n(1)) tail_4227 (
        .y(_T_22),
        .in(_T_21)
    );
    wire _T_23;
    BITS #(.width(4), .high(0), .low(0)) bits_4228 (
        .y(_T_23),
        .in(io_fn)
    );
    wire _T_24;
    BITS #(.width(4), .high(3), .low(3)) bits_4229 (
        .y(_T_24),
        .in(io_fn)
    );
    wire _T_26;
    EQ_UNSIGNED #(.width(1)) u_eq_4230 (
        .y(_T_26),
        .a(_T_24),
        .b(1'h0)
    );
    wire _T_28;
    wire [63:0] _WTEMP_586;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_4231 (
        .y(_WTEMP_586),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(64)) u_eq_4232 (
        .y(_T_28),
        .a(in1_xor_in2),
        .b(_WTEMP_586)
    );
    wire _T_29;
    BITS #(.width(64), .high(63), .low(63)) bits_4233 (
        .y(_T_29),
        .in(io_in1)
    );
    wire _T_30;
    BITS #(.width(64), .high(63), .low(63)) bits_4234 (
        .y(_T_30),
        .in(io_in2)
    );
    wire _T_31;
    EQ_UNSIGNED #(.width(1)) u_eq_4235 (
        .y(_T_31),
        .a(_T_29),
        .b(_T_30)
    );
    wire _T_32;
    BITS #(.width(64), .high(63), .low(63)) bits_4236 (
        .y(_T_32),
        .in(io_adder_out)
    );
    wire _T_33;
    BITS #(.width(4), .high(1), .low(1)) bits_4237 (
        .y(_T_33),
        .in(io_fn)
    );
    wire _T_34;
    BITS #(.width(64), .high(63), .low(63)) bits_4238 (
        .y(_T_34),
        .in(io_in2)
    );
    wire _T_35;
    BITS #(.width(64), .high(63), .low(63)) bits_4239 (
        .y(_T_35),
        .in(io_in1)
    );
    wire _T_36;
    MUX_UNSIGNED #(.width(1)) u_mux_4240 (
        .y(_T_36),
        .sel(_T_33),
        .a(_T_34),
        .b(_T_35)
    );
    wire _T_37;
    MUX_UNSIGNED #(.width(1)) u_mux_4241 (
        .y(_T_37),
        .sel(_T_31),
        .a(_T_32),
        .b(_T_36)
    );
    wire _T_38;
    MUX_UNSIGNED #(.width(1)) u_mux_4242 (
        .y(_T_38),
        .sel(_T_26),
        .a(_T_28),
        .b(_T_37)
    );
    wire _T_39;
    BITWISEXOR #(.width(1)) bitwisexor_4243 (
        .y(_T_39),
        .a(_T_23),
        .b(_T_38)
    );
    wire _T_40;
    BITS #(.width(4), .high(3), .low(3)) bits_4244 (
        .y(_T_40),
        .in(io_fn)
    );
    wire _T_41;
    BITS #(.width(64), .high(31), .low(31)) bits_4245 (
        .y(_T_41),
        .in(io_in1)
    );
    wire _T_42;
    BITWISEAND #(.width(1)) bitwiseand_4246 (
        .y(_T_42),
        .a(_T_40),
        .b(_T_41)
    );
    wire _T_43;
    BITS #(.width(1), .high(0), .low(0)) bits_4247 (
        .y(_T_43),
        .in(_T_42)
    );
    wire [31:0] _T_46;
    MUX_UNSIGNED #(.width(32)) u_mux_4248 (
        .y(_T_46),
        .sel(_T_43),
        .a(32'hFFFFFFFF),
        .b(32'h0)
    );
    wire _T_48;
    EQ_UNSIGNED #(.width(1)) u_eq_4249 (
        .y(_T_48),
        .a(io_dw),
        .b(1'h1)
    );
    wire [31:0] _T_49;
    BITS #(.width(64), .high(63), .low(32)) bits_4250 (
        .y(_T_49),
        .in(io_in1)
    );
    wire [31:0] _T_50;
    MUX_UNSIGNED #(.width(32)) u_mux_4251 (
        .y(_T_50),
        .sel(_T_48),
        .a(_T_49),
        .b(_T_46)
    );
    wire _T_51;
    BITS #(.width(64), .high(5), .low(5)) bits_4252 (
        .y(_T_51),
        .in(io_in2)
    );
    wire _T_53;
    EQ_UNSIGNED #(.width(1)) u_eq_4253 (
        .y(_T_53),
        .a(io_dw),
        .b(1'h1)
    );
    wire _T_54;
    BITWISEAND #(.width(1)) bitwiseand_4254 (
        .y(_T_54),
        .a(_T_51),
        .b(_T_53)
    );
    wire [4:0] _T_55;
    BITS #(.width(64), .high(4), .low(0)) bits_4255 (
        .y(_T_55),
        .in(io_in2)
    );
    wire [5:0] shamt;
    CAT #(.width_a(1), .width_b(5)) cat_4256 (
        .y(shamt),
        .a(_T_54),
        .b(_T_55)
    );
    wire [31:0] _T_56;
    BITS #(.width(64), .high(31), .low(0)) bits_4257 (
        .y(_T_56),
        .in(io_in1)
    );
    wire [63:0] shin_r;
    CAT #(.width_a(32), .width_b(32)) cat_4258 (
        .y(shin_r),
        .a(_T_50),
        .b(_T_56)
    );
    wire _T_58;
    wire [3:0] _WTEMP_587;
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_4259 (
        .y(_WTEMP_587),
        .in(3'h5)
    );
    EQ_UNSIGNED #(.width(4)) u_eq_4260 (
        .y(_T_58),
        .a(io_fn),
        .b(_WTEMP_587)
    );
    wire _T_60;
    EQ_UNSIGNED #(.width(4)) u_eq_4261 (
        .y(_T_60),
        .a(io_fn),
        .b(4'hB)
    );
    wire _T_61;
    BITWISEOR #(.width(1)) bitwiseor_4262 (
        .y(_T_61),
        .a(_T_58),
        .b(_T_60)
    );
    wire [63:0] _T_64;
    assign _T_64 = 64'hFFFFFFFF00000000;
    wire [63:0] _T_65;
    assign _T_65 = 64'hFFFFFFFF;
    wire [31:0] _T_66;
    SHR_UNSIGNED #(.width(64), .n(32)) u_shr_4263 (
        .y(_T_66),
        .in(shin_r)
    );
    wire [63:0] _T_67;
    wire [63:0] _WTEMP_588;
    PAD_UNSIGNED #(.width(32), .n(64)) u_pad_4264 (
        .y(_WTEMP_588),
        .in(_T_66)
    );
    BITWISEAND #(.width(64)) bitwiseand_4265 (
        .y(_T_67),
        .a(_WTEMP_588),
        .b(_T_65)
    );
    wire [31:0] _T_68;
    BITS #(.width(64), .high(31), .low(0)) bits_4266 (
        .y(_T_68),
        .in(shin_r)
    );
    wire [63:0] _T_69;
    SHL_UNSIGNED #(.width(32), .n(32)) u_shl_4267 (
        .y(_T_69),
        .in(_T_68)
    );
    wire [63:0] _T_70;
    assign _T_70 = 64'hFFFFFFFF00000000;
    wire [63:0] _T_71;
    BITWISEAND #(.width(64)) bitwiseand_4268 (
        .y(_T_71),
        .a(_T_69),
        .b(_T_70)
    );
    wire [63:0] _T_72;
    BITWISEOR #(.width(64)) bitwiseor_4269 (
        .y(_T_72),
        .a(_T_67),
        .b(_T_71)
    );
    wire [47:0] _T_73;
    assign _T_73 = 48'hFFFFFFFF;
    wire [63:0] _T_74;
    assign _T_74 = 64'hFFFFFFFF0000;
    wire [63:0] _T_75;
    assign _T_75 = 64'hFFFF0000FFFF;
    wire [47:0] _T_76;
    SHR_UNSIGNED #(.width(64), .n(16)) u_shr_4270 (
        .y(_T_76),
        .in(_T_72)
    );
    wire [63:0] _T_77;
    wire [63:0] _WTEMP_589;
    PAD_UNSIGNED #(.width(48), .n(64)) u_pad_4271 (
        .y(_WTEMP_589),
        .in(_T_76)
    );
    BITWISEAND #(.width(64)) bitwiseand_4272 (
        .y(_T_77),
        .a(_WTEMP_589),
        .b(_T_75)
    );
    wire [47:0] _T_78;
    BITS #(.width(64), .high(47), .low(0)) bits_4273 (
        .y(_T_78),
        .in(_T_72)
    );
    wire [63:0] _T_79;
    SHL_UNSIGNED #(.width(48), .n(16)) u_shl_4274 (
        .y(_T_79),
        .in(_T_78)
    );
    wire [63:0] _T_80;
    assign _T_80 = 64'hFFFF0000FFFF0000;
    wire [63:0] _T_81;
    BITWISEAND #(.width(64)) bitwiseand_4275 (
        .y(_T_81),
        .a(_T_79),
        .b(_T_80)
    );
    wire [63:0] _T_82;
    BITWISEOR #(.width(64)) bitwiseor_4276 (
        .y(_T_82),
        .a(_T_77),
        .b(_T_81)
    );
    wire [55:0] _T_83;
    assign _T_83 = 56'hFFFF0000FFFF;
    wire [63:0] _T_84;
    assign _T_84 = 64'hFFFF0000FFFF00;
    wire [63:0] _T_85;
    assign _T_85 = 64'hFF00FF00FF00FF;
    wire [55:0] _T_86;
    SHR_UNSIGNED #(.width(64), .n(8)) u_shr_4277 (
        .y(_T_86),
        .in(_T_82)
    );
    wire [63:0] _T_87;
    wire [63:0] _WTEMP_590;
    PAD_UNSIGNED #(.width(56), .n(64)) u_pad_4278 (
        .y(_WTEMP_590),
        .in(_T_86)
    );
    BITWISEAND #(.width(64)) bitwiseand_4279 (
        .y(_T_87),
        .a(_WTEMP_590),
        .b(_T_85)
    );
    wire [55:0] _T_88;
    BITS #(.width(64), .high(55), .low(0)) bits_4280 (
        .y(_T_88),
        .in(_T_82)
    );
    wire [63:0] _T_89;
    SHL_UNSIGNED #(.width(56), .n(8)) u_shl_4281 (
        .y(_T_89),
        .in(_T_88)
    );
    wire [63:0] _T_90;
    assign _T_90 = 64'hFF00FF00FF00FF00;
    wire [63:0] _T_91;
    BITWISEAND #(.width(64)) bitwiseand_4282 (
        .y(_T_91),
        .a(_T_89),
        .b(_T_90)
    );
    wire [63:0] _T_92;
    BITWISEOR #(.width(64)) bitwiseor_4283 (
        .y(_T_92),
        .a(_T_87),
        .b(_T_91)
    );
    wire [59:0] _T_93;
    assign _T_93 = 60'hFF00FF00FF00FF;
    wire [63:0] _T_94;
    assign _T_94 = 64'hFF00FF00FF00FF0;
    wire [63:0] _T_95;
    assign _T_95 = 64'hF0F0F0F0F0F0F0F;
    wire [59:0] _T_96;
    SHR_UNSIGNED #(.width(64), .n(4)) u_shr_4284 (
        .y(_T_96),
        .in(_T_92)
    );
    wire [63:0] _T_97;
    wire [63:0] _WTEMP_591;
    PAD_UNSIGNED #(.width(60), .n(64)) u_pad_4285 (
        .y(_WTEMP_591),
        .in(_T_96)
    );
    BITWISEAND #(.width(64)) bitwiseand_4286 (
        .y(_T_97),
        .a(_WTEMP_591),
        .b(_T_95)
    );
    wire [59:0] _T_98;
    BITS #(.width(64), .high(59), .low(0)) bits_4287 (
        .y(_T_98),
        .in(_T_92)
    );
    wire [63:0] _T_99;
    SHL_UNSIGNED #(.width(60), .n(4)) u_shl_4288 (
        .y(_T_99),
        .in(_T_98)
    );
    wire [63:0] _T_100;
    assign _T_100 = 64'hF0F0F0F0F0F0F0F0;
    wire [63:0] _T_101;
    BITWISEAND #(.width(64)) bitwiseand_4289 (
        .y(_T_101),
        .a(_T_99),
        .b(_T_100)
    );
    wire [63:0] _T_102;
    BITWISEOR #(.width(64)) bitwiseor_4290 (
        .y(_T_102),
        .a(_T_97),
        .b(_T_101)
    );
    wire [61:0] _T_103;
    assign _T_103 = 62'hF0F0F0F0F0F0F0F;
    wire [63:0] _T_104;
    assign _T_104 = 64'h3C3C3C3C3C3C3C3C;
    wire [63:0] _T_105;
    assign _T_105 = 64'h3333333333333333;
    wire [61:0] _T_106;
    SHR_UNSIGNED #(.width(64), .n(2)) u_shr_4291 (
        .y(_T_106),
        .in(_T_102)
    );
    wire [63:0] _T_107;
    wire [63:0] _WTEMP_592;
    PAD_UNSIGNED #(.width(62), .n(64)) u_pad_4292 (
        .y(_WTEMP_592),
        .in(_T_106)
    );
    BITWISEAND #(.width(64)) bitwiseand_4293 (
        .y(_T_107),
        .a(_WTEMP_592),
        .b(_T_105)
    );
    wire [61:0] _T_108;
    BITS #(.width(64), .high(61), .low(0)) bits_4294 (
        .y(_T_108),
        .in(_T_102)
    );
    wire [63:0] _T_109;
    SHL_UNSIGNED #(.width(62), .n(2)) u_shl_4295 (
        .y(_T_109),
        .in(_T_108)
    );
    wire [63:0] _T_110;
    assign _T_110 = 64'hCCCCCCCCCCCCCCCC;
    wire [63:0] _T_111;
    BITWISEAND #(.width(64)) bitwiseand_4296 (
        .y(_T_111),
        .a(_T_109),
        .b(_T_110)
    );
    wire [63:0] _T_112;
    BITWISEOR #(.width(64)) bitwiseor_4297 (
        .y(_T_112),
        .a(_T_107),
        .b(_T_111)
    );
    wire [62:0] _T_113;
    assign _T_113 = 63'h3333333333333333;
    wire [63:0] _T_114;
    assign _T_114 = 64'h6666666666666666;
    wire [63:0] _T_115;
    assign _T_115 = 64'h5555555555555555;
    wire [62:0] _T_116;
    SHR_UNSIGNED #(.width(64), .n(1)) u_shr_4298 (
        .y(_T_116),
        .in(_T_112)
    );
    wire [63:0] _T_117;
    wire [63:0] _WTEMP_593;
    PAD_UNSIGNED #(.width(63), .n(64)) u_pad_4299 (
        .y(_WTEMP_593),
        .in(_T_116)
    );
    BITWISEAND #(.width(64)) bitwiseand_4300 (
        .y(_T_117),
        .a(_WTEMP_593),
        .b(_T_115)
    );
    wire [62:0] _T_118;
    BITS #(.width(64), .high(62), .low(0)) bits_4301 (
        .y(_T_118),
        .in(_T_112)
    );
    wire [63:0] _T_119;
    SHL_UNSIGNED #(.width(63), .n(1)) u_shl_4302 (
        .y(_T_119),
        .in(_T_118)
    );
    wire [63:0] _T_120;
    assign _T_120 = 64'hAAAAAAAAAAAAAAAA;
    wire [63:0] _T_121;
    BITWISEAND #(.width(64)) bitwiseand_4303 (
        .y(_T_121),
        .a(_T_119),
        .b(_T_120)
    );
    wire [63:0] _T_122;
    BITWISEOR #(.width(64)) bitwiseor_4304 (
        .y(_T_122),
        .a(_T_117),
        .b(_T_121)
    );
    wire [63:0] shin;
    MUX_UNSIGNED #(.width(64)) u_mux_4305 (
        .y(shin),
        .sel(_T_61),
        .a(shin_r),
        .b(_T_122)
    );
    wire _T_123;
    BITS #(.width(4), .high(3), .low(3)) bits_4306 (
        .y(_T_123),
        .in(io_fn)
    );
    wire _T_124;
    BITS #(.width(64), .high(63), .low(63)) bits_4307 (
        .y(_T_124),
        .in(shin)
    );
    wire _T_125;
    BITWISEAND #(.width(1)) bitwiseand_4308 (
        .y(_T_125),
        .a(_T_123),
        .b(_T_124)
    );
    wire [64:0] _T_126;
    CAT #(.width_a(1), .width_b(64)) cat_4309 (
        .y(_T_126),
        .a(_T_125),
        .b(shin)
    );
    wire [64:0] _T_127;
    ASSINT #(.width(65)) assint_4310 (
        .y(_T_127),
        .in(_T_126)
    );
    wire [64:0] _T_128;
    DSHR_SIGNED #(.width_in(65), .width_n(6)) s_dshr_4311 (
        .y(_T_128),
        .in(_T_127),
        .n(shamt)
    );
    wire [63:0] shout_r;
    BITS #(.width(65), .high(63), .low(0)) bits_4312 (
        .y(shout_r),
        .in(_T_128)
    );
    wire [63:0] _T_131;
    assign _T_131 = 64'hFFFFFFFF00000000;
    wire [63:0] _T_132;
    assign _T_132 = 64'hFFFFFFFF;
    wire [31:0] _T_133;
    SHR_UNSIGNED #(.width(64), .n(32)) u_shr_4313 (
        .y(_T_133),
        .in(shout_r)
    );
    wire [63:0] _T_134;
    wire [63:0] _WTEMP_594;
    PAD_UNSIGNED #(.width(32), .n(64)) u_pad_4314 (
        .y(_WTEMP_594),
        .in(_T_133)
    );
    BITWISEAND #(.width(64)) bitwiseand_4315 (
        .y(_T_134),
        .a(_WTEMP_594),
        .b(_T_132)
    );
    wire [31:0] _T_135;
    BITS #(.width(64), .high(31), .low(0)) bits_4316 (
        .y(_T_135),
        .in(shout_r)
    );
    wire [63:0] _T_136;
    SHL_UNSIGNED #(.width(32), .n(32)) u_shl_4317 (
        .y(_T_136),
        .in(_T_135)
    );
    wire [63:0] _T_137;
    assign _T_137 = 64'hFFFFFFFF00000000;
    wire [63:0] _T_138;
    BITWISEAND #(.width(64)) bitwiseand_4318 (
        .y(_T_138),
        .a(_T_136),
        .b(_T_137)
    );
    wire [63:0] _T_139;
    BITWISEOR #(.width(64)) bitwiseor_4319 (
        .y(_T_139),
        .a(_T_134),
        .b(_T_138)
    );
    wire [47:0] _T_140;
    assign _T_140 = 48'hFFFFFFFF;
    wire [63:0] _T_141;
    assign _T_141 = 64'hFFFFFFFF0000;
    wire [63:0] _T_142;
    assign _T_142 = 64'hFFFF0000FFFF;
    wire [47:0] _T_143;
    SHR_UNSIGNED #(.width(64), .n(16)) u_shr_4320 (
        .y(_T_143),
        .in(_T_139)
    );
    wire [63:0] _T_144;
    wire [63:0] _WTEMP_595;
    PAD_UNSIGNED #(.width(48), .n(64)) u_pad_4321 (
        .y(_WTEMP_595),
        .in(_T_143)
    );
    BITWISEAND #(.width(64)) bitwiseand_4322 (
        .y(_T_144),
        .a(_WTEMP_595),
        .b(_T_142)
    );
    wire [47:0] _T_145;
    BITS #(.width(64), .high(47), .low(0)) bits_4323 (
        .y(_T_145),
        .in(_T_139)
    );
    wire [63:0] _T_146;
    SHL_UNSIGNED #(.width(48), .n(16)) u_shl_4324 (
        .y(_T_146),
        .in(_T_145)
    );
    wire [63:0] _T_147;
    assign _T_147 = 64'hFFFF0000FFFF0000;
    wire [63:0] _T_148;
    BITWISEAND #(.width(64)) bitwiseand_4325 (
        .y(_T_148),
        .a(_T_146),
        .b(_T_147)
    );
    wire [63:0] _T_149;
    BITWISEOR #(.width(64)) bitwiseor_4326 (
        .y(_T_149),
        .a(_T_144),
        .b(_T_148)
    );
    wire [55:0] _T_150;
    assign _T_150 = 56'hFFFF0000FFFF;
    wire [63:0] _T_151;
    assign _T_151 = 64'hFFFF0000FFFF00;
    wire [63:0] _T_152;
    assign _T_152 = 64'hFF00FF00FF00FF;
    wire [55:0] _T_153;
    SHR_UNSIGNED #(.width(64), .n(8)) u_shr_4327 (
        .y(_T_153),
        .in(_T_149)
    );
    wire [63:0] _T_154;
    wire [63:0] _WTEMP_596;
    PAD_UNSIGNED #(.width(56), .n(64)) u_pad_4328 (
        .y(_WTEMP_596),
        .in(_T_153)
    );
    BITWISEAND #(.width(64)) bitwiseand_4329 (
        .y(_T_154),
        .a(_WTEMP_596),
        .b(_T_152)
    );
    wire [55:0] _T_155;
    BITS #(.width(64), .high(55), .low(0)) bits_4330 (
        .y(_T_155),
        .in(_T_149)
    );
    wire [63:0] _T_156;
    SHL_UNSIGNED #(.width(56), .n(8)) u_shl_4331 (
        .y(_T_156),
        .in(_T_155)
    );
    wire [63:0] _T_157;
    assign _T_157 = 64'hFF00FF00FF00FF00;
    wire [63:0] _T_158;
    BITWISEAND #(.width(64)) bitwiseand_4332 (
        .y(_T_158),
        .a(_T_156),
        .b(_T_157)
    );
    wire [63:0] _T_159;
    BITWISEOR #(.width(64)) bitwiseor_4333 (
        .y(_T_159),
        .a(_T_154),
        .b(_T_158)
    );
    wire [59:0] _T_160;
    assign _T_160 = 60'hFF00FF00FF00FF;
    wire [63:0] _T_161;
    assign _T_161 = 64'hFF00FF00FF00FF0;
    wire [63:0] _T_162;
    assign _T_162 = 64'hF0F0F0F0F0F0F0F;
    wire [59:0] _T_163;
    SHR_UNSIGNED #(.width(64), .n(4)) u_shr_4334 (
        .y(_T_163),
        .in(_T_159)
    );
    wire [63:0] _T_164;
    wire [63:0] _WTEMP_597;
    PAD_UNSIGNED #(.width(60), .n(64)) u_pad_4335 (
        .y(_WTEMP_597),
        .in(_T_163)
    );
    BITWISEAND #(.width(64)) bitwiseand_4336 (
        .y(_T_164),
        .a(_WTEMP_597),
        .b(_T_162)
    );
    wire [59:0] _T_165;
    BITS #(.width(64), .high(59), .low(0)) bits_4337 (
        .y(_T_165),
        .in(_T_159)
    );
    wire [63:0] _T_166;
    SHL_UNSIGNED #(.width(60), .n(4)) u_shl_4338 (
        .y(_T_166),
        .in(_T_165)
    );
    wire [63:0] _T_167;
    assign _T_167 = 64'hF0F0F0F0F0F0F0F0;
    wire [63:0] _T_168;
    BITWISEAND #(.width(64)) bitwiseand_4339 (
        .y(_T_168),
        .a(_T_166),
        .b(_T_167)
    );
    wire [63:0] _T_169;
    BITWISEOR #(.width(64)) bitwiseor_4340 (
        .y(_T_169),
        .a(_T_164),
        .b(_T_168)
    );
    wire [61:0] _T_170;
    assign _T_170 = 62'hF0F0F0F0F0F0F0F;
    wire [63:0] _T_171;
    assign _T_171 = 64'h3C3C3C3C3C3C3C3C;
    wire [63:0] _T_172;
    assign _T_172 = 64'h3333333333333333;
    wire [61:0] _T_173;
    SHR_UNSIGNED #(.width(64), .n(2)) u_shr_4341 (
        .y(_T_173),
        .in(_T_169)
    );
    wire [63:0] _T_174;
    wire [63:0] _WTEMP_598;
    PAD_UNSIGNED #(.width(62), .n(64)) u_pad_4342 (
        .y(_WTEMP_598),
        .in(_T_173)
    );
    BITWISEAND #(.width(64)) bitwiseand_4343 (
        .y(_T_174),
        .a(_WTEMP_598),
        .b(_T_172)
    );
    wire [61:0] _T_175;
    BITS #(.width(64), .high(61), .low(0)) bits_4344 (
        .y(_T_175),
        .in(_T_169)
    );
    wire [63:0] _T_176;
    SHL_UNSIGNED #(.width(62), .n(2)) u_shl_4345 (
        .y(_T_176),
        .in(_T_175)
    );
    wire [63:0] _T_177;
    assign _T_177 = 64'hCCCCCCCCCCCCCCCC;
    wire [63:0] _T_178;
    BITWISEAND #(.width(64)) bitwiseand_4346 (
        .y(_T_178),
        .a(_T_176),
        .b(_T_177)
    );
    wire [63:0] _T_179;
    BITWISEOR #(.width(64)) bitwiseor_4347 (
        .y(_T_179),
        .a(_T_174),
        .b(_T_178)
    );
    wire [62:0] _T_180;
    assign _T_180 = 63'h3333333333333333;
    wire [63:0] _T_181;
    assign _T_181 = 64'h6666666666666666;
    wire [63:0] _T_182;
    assign _T_182 = 64'h5555555555555555;
    wire [62:0] _T_183;
    SHR_UNSIGNED #(.width(64), .n(1)) u_shr_4348 (
        .y(_T_183),
        .in(_T_179)
    );
    wire [63:0] _T_184;
    wire [63:0] _WTEMP_599;
    PAD_UNSIGNED #(.width(63), .n(64)) u_pad_4349 (
        .y(_WTEMP_599),
        .in(_T_183)
    );
    BITWISEAND #(.width(64)) bitwiseand_4350 (
        .y(_T_184),
        .a(_WTEMP_599),
        .b(_T_182)
    );
    wire [62:0] _T_185;
    BITS #(.width(64), .high(62), .low(0)) bits_4351 (
        .y(_T_185),
        .in(_T_179)
    );
    wire [63:0] _T_186;
    SHL_UNSIGNED #(.width(63), .n(1)) u_shl_4352 (
        .y(_T_186),
        .in(_T_185)
    );
    wire [63:0] _T_187;
    assign _T_187 = 64'hAAAAAAAAAAAAAAAA;
    wire [63:0] _T_188;
    BITWISEAND #(.width(64)) bitwiseand_4353 (
        .y(_T_188),
        .a(_T_186),
        .b(_T_187)
    );
    wire [63:0] shout_l;
    BITWISEOR #(.width(64)) bitwiseor_4354 (
        .y(shout_l),
        .a(_T_184),
        .b(_T_188)
    );
    wire _T_190;
    wire [3:0] _WTEMP_600;
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_4355 (
        .y(_WTEMP_600),
        .in(3'h5)
    );
    EQ_UNSIGNED #(.width(4)) u_eq_4356 (
        .y(_T_190),
        .a(io_fn),
        .b(_WTEMP_600)
    );
    wire _T_192;
    EQ_UNSIGNED #(.width(4)) u_eq_4357 (
        .y(_T_192),
        .a(io_fn),
        .b(4'hB)
    );
    wire _T_193;
    BITWISEOR #(.width(1)) bitwiseor_4358 (
        .y(_T_193),
        .a(_T_190),
        .b(_T_192)
    );
    wire [63:0] _T_195;
    wire [63:0] _WTEMP_601;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_4359 (
        .y(_WTEMP_601),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_4360 (
        .y(_T_195),
        .sel(_T_193),
        .a(shout_r),
        .b(_WTEMP_601)
    );
    wire _T_197;
    wire [3:0] _WTEMP_602;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_4361 (
        .y(_WTEMP_602),
        .in(1'h1)
    );
    EQ_UNSIGNED #(.width(4)) u_eq_4362 (
        .y(_T_197),
        .a(io_fn),
        .b(_WTEMP_602)
    );
    wire [63:0] _T_199;
    wire [63:0] _WTEMP_603;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_4363 (
        .y(_WTEMP_603),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_4364 (
        .y(_T_199),
        .sel(_T_197),
        .a(shout_l),
        .b(_WTEMP_603)
    );
    wire [63:0] shout;
    BITWISEOR #(.width(64)) bitwiseor_4365 (
        .y(shout),
        .a(_T_195),
        .b(_T_199)
    );
    wire _T_201;
    wire [3:0] _WTEMP_604;
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_4366 (
        .y(_WTEMP_604),
        .in(3'h4)
    );
    EQ_UNSIGNED #(.width(4)) u_eq_4367 (
        .y(_T_201),
        .a(io_fn),
        .b(_WTEMP_604)
    );
    wire _T_203;
    wire [3:0] _WTEMP_605;
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_4368 (
        .y(_WTEMP_605),
        .in(3'h6)
    );
    EQ_UNSIGNED #(.width(4)) u_eq_4369 (
        .y(_T_203),
        .a(io_fn),
        .b(_WTEMP_605)
    );
    wire _T_204;
    BITWISEOR #(.width(1)) bitwiseor_4370 (
        .y(_T_204),
        .a(_T_201),
        .b(_T_203)
    );
    wire [63:0] _T_206;
    wire [63:0] _WTEMP_606;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_4371 (
        .y(_WTEMP_606),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_4372 (
        .y(_T_206),
        .sel(_T_204),
        .a(in1_xor_in2),
        .b(_WTEMP_606)
    );
    wire _T_208;
    wire [3:0] _WTEMP_607;
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_4373 (
        .y(_WTEMP_607),
        .in(3'h6)
    );
    EQ_UNSIGNED #(.width(4)) u_eq_4374 (
        .y(_T_208),
        .a(io_fn),
        .b(_WTEMP_607)
    );
    wire _T_210;
    wire [3:0] _WTEMP_608;
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_4375 (
        .y(_WTEMP_608),
        .in(3'h7)
    );
    EQ_UNSIGNED #(.width(4)) u_eq_4376 (
        .y(_T_210),
        .a(io_fn),
        .b(_WTEMP_608)
    );
    wire _T_211;
    BITWISEOR #(.width(1)) bitwiseor_4377 (
        .y(_T_211),
        .a(_T_208),
        .b(_T_210)
    );
    wire [63:0] _T_212;
    BITWISEAND #(.width(64)) bitwiseand_4378 (
        .y(_T_212),
        .a(io_in1),
        .b(io_in2)
    );
    wire [63:0] _T_214;
    wire [63:0] _WTEMP_609;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_4379 (
        .y(_WTEMP_609),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_4380 (
        .y(_T_214),
        .sel(_T_211),
        .a(_T_212),
        .b(_WTEMP_609)
    );
    wire [63:0] logic_;
    BITWISEOR #(.width(64)) bitwiseor_4381 (
        .y(logic_),
        .a(_T_206),
        .b(_T_214)
    );
    wire _T_216;
    wire [3:0] _WTEMP_610;
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_4382 (
        .y(_WTEMP_610),
        .in(2'h2)
    );
    EQ_UNSIGNED #(.width(4)) u_eq_4383 (
        .y(_T_216),
        .a(io_fn),
        .b(_WTEMP_610)
    );
    wire _T_218;
    wire [3:0] _WTEMP_611;
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_4384 (
        .y(_WTEMP_611),
        .in(2'h3)
    );
    EQ_UNSIGNED #(.width(4)) u_eq_4385 (
        .y(_T_218),
        .a(io_fn),
        .b(_WTEMP_611)
    );
    wire _T_219;
    BITWISEOR #(.width(1)) bitwiseor_4386 (
        .y(_T_219),
        .a(_T_216),
        .b(_T_218)
    );
    wire _T_221;
    GEQ_UNSIGNED #(.width(4)) u_geq_4387 (
        .y(_T_221),
        .a(io_fn),
        .b(4'hC)
    );
    wire _T_222;
    BITWISEOR #(.width(1)) bitwiseor_4388 (
        .y(_T_222),
        .a(_T_219),
        .b(_T_221)
    );
    wire _T_223;
    BITWISEAND #(.width(1)) bitwiseand_4389 (
        .y(_T_223),
        .a(_T_222),
        .b(io_cmp_out)
    );
    wire [63:0] _T_224;
    wire [63:0] _WTEMP_612;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_4390 (
        .y(_WTEMP_612),
        .in(_T_223)
    );
    BITWISEOR #(.width(64)) bitwiseor_4391 (
        .y(_T_224),
        .a(_WTEMP_612),
        .b(logic_)
    );
    wire [63:0] shift_logic;
    BITWISEOR #(.width(64)) bitwiseor_4392 (
        .y(shift_logic),
        .a(_T_224),
        .b(shout)
    );
    wire _T_226;
    wire [3:0] _WTEMP_613;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_4393 (
        .y(_WTEMP_613),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(4)) u_eq_4394 (
        .y(_T_226),
        .a(io_fn),
        .b(_WTEMP_613)
    );
    wire _T_228;
    EQ_UNSIGNED #(.width(4)) u_eq_4395 (
        .y(_T_228),
        .a(io_fn),
        .b(4'hA)
    );
    wire _T_229;
    BITWISEOR #(.width(1)) bitwiseor_4396 (
        .y(_T_229),
        .a(_T_226),
        .b(_T_228)
    );
    wire [63:0] out;
    MUX_UNSIGNED #(.width(64)) u_mux_4397 (
        .y(out),
        .sel(_T_229),
        .a(io_adder_out),
        .b(shift_logic)
    );
    wire _T_231;
    EQ_UNSIGNED #(.width(1)) u_eq_4398 (
        .y(_T_231),
        .a(io_dw),
        .b(1'h0)
    );
    wire _T_232;
    BITS #(.width(64), .high(31), .low(31)) bits_4399 (
        .y(_T_232),
        .in(out)
    );
    wire _T_233;
    BITS #(.width(1), .high(0), .low(0)) bits_4400 (
        .y(_T_233),
        .in(_T_232)
    );
    wire [31:0] _T_236;
    MUX_UNSIGNED #(.width(32)) u_mux_4401 (
        .y(_T_236),
        .sel(_T_233),
        .a(32'hFFFFFFFF),
        .b(32'h0)
    );
    wire [31:0] _T_237;
    BITS #(.width(64), .high(31), .low(0)) bits_4402 (
        .y(_T_237),
        .in(out)
    );
    wire [63:0] _T_238;
    CAT #(.width_a(32), .width_b(32)) cat_4403 (
        .y(_T_238),
        .a(_T_236),
        .b(_T_237)
    );
    assign io_adder_out = _T_22;
    assign io_cmp_out = _T_39;
    MUX_UNSIGNED #(.width(64)) u_mux_4404 (
        .y(io_out),
        .sel(_T_231),
        .a(_T_238),
        .b(out)
    );
endmodule //ALU
module DSHR_SIGNED(y, in, n);
    parameter width_in = 4;
    parameter width_n = 2;
    output [width_in-1:0] y;
    input [width_in-1:0] in;
    input [width_n-1:0] n;
    assign y = $signed(in) >>> n;
endmodule // DSHR_SIGNED
module MulDiv(
    input clock,
    input reset,
    output io_req_ready,
    input io_req_valid,
    input [3:0] io_req_bits_fn,
    input io_req_bits_dw,
    input [63:0] io_req_bits_in1,
    input [63:0] io_req_bits_in2,
    input [4:0] io_req_bits_tag,
    input io_kill,
    input io_resp_ready,
    output io_resp_valid,
    output [63:0] io_resp_bits_data,
    output [4:0] io_resp_bits_tag
);
    wire [2:0] _state__q;
    wire [2:0] _state__d;
    DFF_POSCLK #(.width(3)) state (
        .q(_state__q),
        .d(_state__d),
        .clk(clock)
    );
    wire [2:0] _WTEMP_614;
    MUX_UNSIGNED #(.width(3)) u_mux_4407 (
        .y(_state__d),
        .sel(reset),
        .a(3'h0),
        .b(_WTEMP_614)
    );
    wire [3:0] _req_fn__q;
    wire [3:0] _req_fn__d;
    DFF_POSCLK #(.width(4)) req_fn (
        .q(_req_fn__q),
        .d(_req_fn__d),
        .clk(clock)
    );
    wire _req_dw__q;
    wire _req_dw__d;
    DFF_POSCLK #(.width(1)) req_dw (
        .q(_req_dw__q),
        .d(_req_dw__d),
        .clk(clock)
    );
    wire [63:0] _req_in1__q;
    wire [63:0] _req_in1__d;
    DFF_POSCLK #(.width(64)) req_in1 (
        .q(_req_in1__q),
        .d(_req_in1__d),
        .clk(clock)
    );
    wire [63:0] _req_in2__q;
    wire [63:0] _req_in2__d;
    DFF_POSCLK #(.width(64)) req_in2 (
        .q(_req_in2__q),
        .d(_req_in2__d),
        .clk(clock)
    );
    wire [4:0] _req_tag__q;
    wire [4:0] _req_tag__d;
    DFF_POSCLK #(.width(5)) req_tag (
        .q(_req_tag__q),
        .d(_req_tag__d),
        .clk(clock)
    );
    wire [6:0] _count__q;
    wire [6:0] _count__d;
    DFF_POSCLK #(.width(7)) count (
        .q(_count__q),
        .d(_count__d),
        .clk(clock)
    );
    wire _neg_out__q;
    wire _neg_out__d;
    DFF_POSCLK #(.width(1)) neg_out (
        .q(_neg_out__q),
        .d(_neg_out__d),
        .clk(clock)
    );
    wire _isMul__q;
    wire _isMul__d;
    DFF_POSCLK #(.width(1)) isMul (
        .q(_isMul__q),
        .d(_isMul__d),
        .clk(clock)
    );
    wire _isHi__q;
    wire _isHi__d;
    DFF_POSCLK #(.width(1)) isHi (
        .q(_isHi__q),
        .d(_isHi__d),
        .clk(clock)
    );
    wire [64:0] _divisor__q;
    wire [64:0] _divisor__d;
    DFF_POSCLK #(.width(65)) divisor (
        .q(_divisor__q),
        .d(_divisor__d),
        .clk(clock)
    );
    wire [129:0] _remainder__q;
    wire [129:0] _remainder__d;
    DFF_POSCLK #(.width(130)) remainder (
        .q(_remainder__q),
        .d(_remainder__d),
        .clk(clock)
    );
    wire [3:0] _T_79;
    BITWISEAND #(.width(4)) bitwiseand_4408 (
        .y(_T_79),
        .a(io_req_bits_fn),
        .b(4'h4)
    );
    wire _T_81;
    EQ_UNSIGNED #(.width(4)) u_eq_4409 (
        .y(_T_81),
        .a(_T_79),
        .b(4'h0)
    );
    wire [3:0] _T_83;
    BITWISEAND #(.width(4)) bitwiseand_4410 (
        .y(_T_83),
        .a(io_req_bits_fn),
        .b(4'h8)
    );
    wire _T_85;
    EQ_UNSIGNED #(.width(4)) u_eq_4411 (
        .y(_T_85),
        .a(_T_83),
        .b(4'h8)
    );
    wire _T_87;
    BITWISEOR #(.width(1)) bitwiseor_4412 (
        .y(_T_87),
        .a(1'h0),
        .b(_T_81)
    );
    wire _T_88;
    BITWISEOR #(.width(1)) bitwiseor_4413 (
        .y(_T_88),
        .a(_T_87),
        .b(_T_85)
    );
    wire [3:0] _T_90;
    BITWISEAND #(.width(4)) bitwiseand_4414 (
        .y(_T_90),
        .a(io_req_bits_fn),
        .b(4'h5)
    );
    wire _T_92;
    EQ_UNSIGNED #(.width(4)) u_eq_4415 (
        .y(_T_92),
        .a(_T_90),
        .b(4'h1)
    );
    wire [3:0] _T_94;
    BITWISEAND #(.width(4)) bitwiseand_4416 (
        .y(_T_94),
        .a(io_req_bits_fn),
        .b(4'h2)
    );
    wire _T_96;
    EQ_UNSIGNED #(.width(4)) u_eq_4417 (
        .y(_T_96),
        .a(_T_94),
        .b(4'h2)
    );
    wire _T_98;
    BITWISEOR #(.width(1)) bitwiseor_4418 (
        .y(_T_98),
        .a(1'h0),
        .b(_T_92)
    );
    wire _T_99;
    BITWISEOR #(.width(1)) bitwiseor_4419 (
        .y(_T_99),
        .a(_T_98),
        .b(_T_96)
    );
    wire _T_100;
    BITWISEOR #(.width(1)) bitwiseor_4420 (
        .y(_T_100),
        .a(_T_99),
        .b(_T_85)
    );
    wire [3:0] _T_102;
    BITWISEAND #(.width(4)) bitwiseand_4421 (
        .y(_T_102),
        .a(io_req_bits_fn),
        .b(4'h9)
    );
    wire _T_104;
    EQ_UNSIGNED #(.width(4)) u_eq_4422 (
        .y(_T_104),
        .a(_T_102),
        .b(4'h0)
    );
    wire [3:0] _T_106;
    BITWISEAND #(.width(4)) bitwiseand_4423 (
        .y(_T_106),
        .a(io_req_bits_fn),
        .b(4'h3)
    );
    wire _T_108;
    EQ_UNSIGNED #(.width(4)) u_eq_4424 (
        .y(_T_108),
        .a(_T_106),
        .b(4'h0)
    );
    wire _T_110;
    BITWISEOR #(.width(1)) bitwiseor_4425 (
        .y(_T_110),
        .a(1'h0),
        .b(_T_104)
    );
    wire _T_111;
    BITWISEOR #(.width(1)) bitwiseor_4426 (
        .y(_T_111),
        .a(_T_110),
        .b(_T_81)
    );
    wire _T_112;
    BITWISEOR #(.width(1)) bitwiseor_4427 (
        .y(_T_112),
        .a(_T_111),
        .b(_T_108)
    );
    wire _T_114;
    BITWISEOR #(.width(1)) bitwiseor_4428 (
        .y(_T_114),
        .a(1'h0),
        .b(_T_104)
    );
    wire _T_115;
    BITWISEOR #(.width(1)) bitwiseor_4429 (
        .y(_T_115),
        .a(_T_114),
        .b(_T_81)
    );
    wire cmdMul;
    BITS #(.width(1), .high(0), .low(0)) bits_4430 (
        .y(cmdMul),
        .in(_T_88)
    );
    wire cmdHi;
    BITS #(.width(1), .high(0), .low(0)) bits_4431 (
        .y(cmdHi),
        .in(_T_100)
    );
    wire lhsSigned;
    BITS #(.width(1), .high(0), .low(0)) bits_4432 (
        .y(lhsSigned),
        .in(_T_112)
    );
    wire rhsSigned;
    BITS #(.width(1), .high(0), .low(0)) bits_4433 (
        .y(rhsSigned),
        .in(_T_115)
    );
    wire _T_118;
    EQ_UNSIGNED #(.width(1)) u_eq_4434 (
        .y(_T_118),
        .a(io_req_bits_dw),
        .b(1'h0)
    );
    wire _T_119;
    BITWISEAND #(.width(1)) bitwiseand_4435 (
        .y(_T_119),
        .a(1'h1),
        .b(_T_118)
    );
    wire _T_120;
    BITS #(.width(64), .high(31), .low(31)) bits_4436 (
        .y(_T_120),
        .in(io_req_bits_in1)
    );
    wire _T_121;
    BITS #(.width(64), .high(63), .low(63)) bits_4437 (
        .y(_T_121),
        .in(io_req_bits_in1)
    );
    wire _T_122;
    MUX_UNSIGNED #(.width(1)) u_mux_4438 (
        .y(_T_122),
        .sel(_T_119),
        .a(_T_120),
        .b(_T_121)
    );
    wire lhs_sign;
    BITWISEAND #(.width(1)) bitwiseand_4439 (
        .y(lhs_sign),
        .a(lhsSigned),
        .b(_T_122)
    );
    wire _T_123;
    BITS #(.width(1), .high(0), .low(0)) bits_4440 (
        .y(_T_123),
        .in(lhs_sign)
    );
    wire [31:0] _T_126;
    MUX_UNSIGNED #(.width(32)) u_mux_4441 (
        .y(_T_126),
        .sel(_T_123),
        .a(32'hFFFFFFFF),
        .b(32'h0)
    );
    wire [31:0] _T_127;
    BITS #(.width(64), .high(63), .low(32)) bits_4442 (
        .y(_T_127),
        .in(io_req_bits_in1)
    );
    wire [31:0] _T_128;
    MUX_UNSIGNED #(.width(32)) u_mux_4443 (
        .y(_T_128),
        .sel(_T_119),
        .a(_T_126),
        .b(_T_127)
    );
    wire [31:0] _T_129;
    BITS #(.width(64), .high(31), .low(0)) bits_4444 (
        .y(_T_129),
        .in(io_req_bits_in1)
    );
    wire [63:0] lhs_in;
    CAT #(.width_a(32), .width_b(32)) cat_4445 (
        .y(lhs_in),
        .a(_T_128),
        .b(_T_129)
    );
    wire _T_132;
    EQ_UNSIGNED #(.width(1)) u_eq_4446 (
        .y(_T_132),
        .a(io_req_bits_dw),
        .b(1'h0)
    );
    wire _T_133;
    BITWISEAND #(.width(1)) bitwiseand_4447 (
        .y(_T_133),
        .a(1'h1),
        .b(_T_132)
    );
    wire _T_134;
    BITS #(.width(64), .high(31), .low(31)) bits_4448 (
        .y(_T_134),
        .in(io_req_bits_in2)
    );
    wire _T_135;
    BITS #(.width(64), .high(63), .low(63)) bits_4449 (
        .y(_T_135),
        .in(io_req_bits_in2)
    );
    wire _T_136;
    MUX_UNSIGNED #(.width(1)) u_mux_4450 (
        .y(_T_136),
        .sel(_T_133),
        .a(_T_134),
        .b(_T_135)
    );
    wire rhs_sign;
    BITWISEAND #(.width(1)) bitwiseand_4451 (
        .y(rhs_sign),
        .a(rhsSigned),
        .b(_T_136)
    );
    wire _T_137;
    BITS #(.width(1), .high(0), .low(0)) bits_4452 (
        .y(_T_137),
        .in(rhs_sign)
    );
    wire [31:0] _T_140;
    MUX_UNSIGNED #(.width(32)) u_mux_4453 (
        .y(_T_140),
        .sel(_T_137),
        .a(32'hFFFFFFFF),
        .b(32'h0)
    );
    wire [31:0] _T_141;
    BITS #(.width(64), .high(63), .low(32)) bits_4454 (
        .y(_T_141),
        .in(io_req_bits_in2)
    );
    wire [31:0] _T_142;
    MUX_UNSIGNED #(.width(32)) u_mux_4455 (
        .y(_T_142),
        .sel(_T_133),
        .a(_T_140),
        .b(_T_141)
    );
    wire [31:0] _T_143;
    BITS #(.width(64), .high(31), .low(0)) bits_4456 (
        .y(_T_143),
        .in(io_req_bits_in2)
    );
    wire [63:0] rhs_in;
    CAT #(.width_a(32), .width_b(32)) cat_4457 (
        .y(rhs_in),
        .a(_T_142),
        .b(_T_143)
    );
    wire [64:0] _T_144;
    BITS #(.width(130), .high(128), .low(64)) bits_4458 (
        .y(_T_144),
        .in(_remainder__q)
    );
    wire [65:0] _T_145;
    SUB_UNSIGNED #(.width(65)) u_sub_4459 (
        .y(_T_145),
        .a(_T_144),
        .b(_divisor__q)
    );
    wire [65:0] _T_146;
    ASUINT #(.width(66)) asuint_4460 (
        .y(_T_146),
        .in(_T_145)
    );
    wire [64:0] subtractor;
    TAIL #(.width(66), .n(1)) tail_4461 (
        .y(subtractor),
        .in(_T_146)
    );
    wire [63:0] _T_147;
    BITS #(.width(130), .high(63), .low(0)) bits_4462 (
        .y(_T_147),
        .in(_remainder__q)
    );
    wire [64:0] _T_149;
    wire [63:0] _WTEMP_615;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_4463 (
        .y(_WTEMP_615),
        .in(1'h0)
    );
    SUB_UNSIGNED #(.width(64)) u_sub_4464 (
        .y(_T_149),
        .a(_WTEMP_615),
        .b(_T_147)
    );
    wire [64:0] _T_150;
    ASUINT #(.width(65)) asuint_4465 (
        .y(_T_150),
        .in(_T_149)
    );
    wire [63:0] negated_remainder;
    TAIL #(.width(65), .n(1)) tail_4466 (
        .y(negated_remainder),
        .in(_T_150)
    );
    wire _T_151;
    EQ_UNSIGNED #(.width(3)) u_eq_4467 (
        .y(_T_151),
        .a(_state__q),
        .b(3'h1)
    );
    wire _T_152;
    BITS #(.width(130), .high(63), .low(63)) bits_4468 (
        .y(_T_152),
        .in(_remainder__q)
    );
    wire _T_153;
    BITWISEOR #(.width(1)) bitwiseor_4469 (
        .y(_T_153),
        .a(_T_152),
        .b(_isMul__q)
    );
    wire _T_154;
    BITS #(.width(65), .high(63), .low(63)) bits_4470 (
        .y(_T_154),
        .in(_divisor__q)
    );
    wire _T_155;
    BITWISEOR #(.width(1)) bitwiseor_4471 (
        .y(_T_155),
        .a(_T_154),
        .b(_isMul__q)
    );
    wire [64:0] _node_340;
    MUX_UNSIGNED #(.width(65)) u_mux_4472 (
        .y(_node_340),
        .sel(_T_155),
        .a(subtractor),
        .b(_divisor__q)
    );
    wire [129:0] _node_341;
    wire [129:0] _WTEMP_616;
    PAD_UNSIGNED #(.width(64), .n(130)) u_pad_4473 (
        .y(_WTEMP_616),
        .in(negated_remainder)
    );
    MUX_UNSIGNED #(.width(130)) u_mux_4474 (
        .y(_node_341),
        .sel(_T_153),
        .a(_WTEMP_616),
        .b(_remainder__q)
    );
    wire _T_156;
    EQ_UNSIGNED #(.width(3)) u_eq_4475 (
        .y(_T_156),
        .a(_state__q),
        .b(3'h4)
    );
    wire [129:0] _node_342;
    MUX_UNSIGNED #(.width(130)) u_mux_4476 (
        .y(_node_342),
        .sel(_T_151),
        .a(_node_341),
        .b(_remainder__q)
    );
    wire [2:0] _node_343;
    MUX_UNSIGNED #(.width(3)) u_mux_4477 (
        .y(_node_343),
        .sel(_T_151),
        .a(3'h2),
        .b(_state__q)
    );
    wire _T_157;
    EQ_UNSIGNED #(.width(3)) u_eq_4478 (
        .y(_T_157),
        .a(_state__q),
        .b(3'h3)
    );
    wire [63:0] _T_158;
    BITS #(.width(130), .high(128), .low(65)) bits_4479 (
        .y(_T_158),
        .in(_remainder__q)
    );
    wire [2:0] _T_159;
    MUX_UNSIGNED #(.width(3)) u_mux_4480 (
        .y(_T_159),
        .sel(_neg_out__q),
        .a(3'h4),
        .b(3'h5)
    );
    wire [129:0] _node_344;
    wire [129:0] _WTEMP_617;
    PAD_UNSIGNED #(.width(64), .n(130)) u_pad_4481 (
        .y(_WTEMP_617),
        .in(negated_remainder)
    );
    MUX_UNSIGNED #(.width(130)) u_mux_4482 (
        .y(_node_344),
        .sel(_T_156),
        .a(_WTEMP_617),
        .b(_node_342)
    );
    wire [2:0] _node_345;
    MUX_UNSIGNED #(.width(3)) u_mux_4483 (
        .y(_node_345),
        .sel(_T_156),
        .a(3'h5),
        .b(_node_343)
    );
    wire _T_160;
    EQ_UNSIGNED #(.width(3)) u_eq_4484 (
        .y(_T_160),
        .a(_state__q),
        .b(3'h2)
    );
    wire _T_161;
    BITWISEAND #(.width(1)) bitwiseand_4485 (
        .y(_T_161),
        .a(_T_160),
        .b(_isMul__q)
    );
    wire [64:0] _T_162;
    BITS #(.width(130), .high(129), .low(65)) bits_4486 (
        .y(_T_162),
        .in(_remainder__q)
    );
    wire [63:0] _T_163;
    BITS #(.width(130), .high(63), .low(0)) bits_4487 (
        .y(_T_163),
        .in(_remainder__q)
    );
    wire [128:0] _T_164;
    CAT #(.width_a(65), .width_b(64)) cat_4488 (
        .y(_T_164),
        .a(_T_162),
        .b(_T_163)
    );
    wire [63:0] _T_165;
    BITS #(.width(129), .high(63), .low(0)) bits_4489 (
        .y(_T_165),
        .in(_T_164)
    );
    wire [64:0] _T_166;
    BITS #(.width(129), .high(128), .low(64)) bits_4490 (
        .y(_T_166),
        .in(_T_164)
    );
    wire [64:0] _T_167;
    ASSINT #(.width(65)) assint_4491 (
        .y(_T_167),
        .in(_T_166)
    );
    wire [64:0] _T_168;
    ASSINT #(.width(65)) assint_4492 (
        .y(_T_168),
        .in(_divisor__q)
    );
    wire [7:0] _T_169;
    BITS #(.width(64), .high(7), .low(0)) bits_4493 (
        .y(_T_169),
        .in(_T_165)
    );
    wire [7:0] _M_170;
    ASSINT #(.width(8)) assint_4494 (
        .y(_M_170),
        .in(_T_169)
    );
    wire [72:0] _T_170;
    MUL2_SIGNED #(.width_a(65), .width_b(8)) s_mul2_4495 (
        .y(_T_170),
        .a(_T_168),
        .b(_M_170)
    );
    wire [73:0] _T_171;
    wire [72:0] _WTEMP_618;
    PAD_SIGNED #(.width(65), .n(73)) s_pad_4496 (
        .y(_WTEMP_618),
        .in(_T_167)
    );
    ADD_SIGNED #(.width(73)) s_add_4497 (
        .y(_T_171),
        .a(_T_170),
        .b(_WTEMP_618)
    );
    wire [72:0] _T_172;
    TAIL #(.width(74), .n(1)) tail_4498 (
        .y(_T_172),
        .in(_T_171)
    );
    wire [72:0] _T_173;
    ASSINT #(.width(73)) assint_4499 (
        .y(_T_173),
        .in(_T_172)
    );
    wire [55:0] _T_174;
    BITS #(.width(64), .high(63), .low(8)) bits_4500 (
        .y(_T_174),
        .in(_T_165)
    );
    wire [72:0] _T_175;
    ASUINT #(.width(73)) asuint_4501 (
        .y(_T_175),
        .in(_T_173)
    );
    wire [128:0] _T_176;
    CAT #(.width_a(73), .width_b(56)) cat_4502 (
        .y(_T_176),
        .a(_T_175),
        .b(_T_174)
    );
    wire [10:0] _T_179;
    MUL2_UNSIGNED #(.width_a(7), .width_b(4)) u_mul2_4503 (
        .y(_T_179),
        .a(_count__q),
        .b(4'h8)
    );
    wire [5:0] _T_180;
    BITS #(.width(11), .high(5), .low(0)) bits_4504 (
        .y(_T_180),
        .in(_T_179)
    );
    wire [64:0] _T_181;
    DSHR_SIGNED #(.width_in(65), .width_n(6)) s_dshr_4505 (
        .y(_T_181),
        .in(-65'sh10000000000000000),
        .n(_T_180)
    );
    wire [63:0] _T_182;
    BITS #(.width(65), .high(63), .low(0)) bits_4506 (
        .y(_T_182),
        .in(_T_181)
    );
    wire _T_185;
    wire [6:0] _WTEMP_619;
    PAD_UNSIGNED #(.width(3), .n(7)) u_pad_4507 (
        .y(_WTEMP_619),
        .in(3'h7)
    );
    NEQ_UNSIGNED #(.width(7)) u_neq_4508 (
        .y(_T_185),
        .a(_count__q),
        .b(_WTEMP_619)
    );
    wire _T_186;
    BITWISEAND #(.width(1)) bitwiseand_4509 (
        .y(_T_186),
        .a(1'h1),
        .b(_T_185)
    );
    wire _T_188;
    wire [6:0] _WTEMP_620;
    PAD_UNSIGNED #(.width(1), .n(7)) u_pad_4510 (
        .y(_WTEMP_620),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(7)) u_neq_4511 (
        .y(_T_188),
        .a(_count__q),
        .b(_WTEMP_620)
    );
    wire _T_189;
    BITWISEAND #(.width(1)) bitwiseand_4512 (
        .y(_T_189),
        .a(_T_186),
        .b(_T_188)
    );
    wire _T_191;
    EQ_UNSIGNED #(.width(1)) u_eq_4513 (
        .y(_T_191),
        .a(_isHi__q),
        .b(1'h0)
    );
    wire _T_192;
    BITWISEAND #(.width(1)) bitwiseand_4514 (
        .y(_T_192),
        .a(_T_189),
        .b(_T_191)
    );
    wire [63:0] _T_193;
    BITWISENOT #(.width(64)) bitwisenot_4515 (
        .y(_T_193),
        .in(_T_182)
    );
    wire [63:0] _T_194;
    BITWISEAND #(.width(64)) bitwiseand_4516 (
        .y(_T_194),
        .a(_T_165),
        .b(_T_193)
    );
    wire _T_196;
    wire [63:0] _WTEMP_621;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_4517 (
        .y(_WTEMP_621),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(64)) u_eq_4518 (
        .y(_T_196),
        .a(_T_194),
        .b(_WTEMP_621)
    );
    wire _T_197;
    BITWISEAND #(.width(1)) bitwiseand_4519 (
        .y(_T_197),
        .a(_T_192),
        .b(_T_196)
    );
    wire [10:0] _T_200;
    MUL2_UNSIGNED #(.width_a(7), .width_b(4)) u_mul2_4520 (
        .y(_T_200),
        .a(_count__q),
        .b(4'h8)
    );
    wire [11:0] _T_201;
    wire [10:0] _WTEMP_622;
    PAD_UNSIGNED #(.width(7), .n(11)) u_pad_4521 (
        .y(_WTEMP_622),
        .in(7'h40)
    );
    SUB_UNSIGNED #(.width(11)) u_sub_4522 (
        .y(_T_201),
        .a(_WTEMP_622),
        .b(_T_200)
    );
    wire [11:0] _T_202;
    ASUINT #(.width(12)) asuint_4523 (
        .y(_T_202),
        .in(_T_201)
    );
    wire [10:0] _T_203;
    TAIL #(.width(12), .n(1)) tail_4524 (
        .y(_T_203),
        .in(_T_202)
    );
    wire [5:0] _T_204;
    BITS #(.width(11), .high(5), .low(0)) bits_4525 (
        .y(_T_204),
        .in(_T_203)
    );
    wire [128:0] _T_205;
    DSHR_UNSIGNED #(.width_in(129), .width_n(6)) u_dshr_4526 (
        .y(_T_205),
        .in(_T_164),
        .n(_T_204)
    );
    wire [64:0] _T_206;
    BITS #(.width(129), .high(128), .low(64)) bits_4527 (
        .y(_T_206),
        .in(_T_176)
    );
    wire [128:0] _T_207;
    MUX_UNSIGNED #(.width(129)) u_mux_4528 (
        .y(_T_207),
        .sel(_T_197),
        .a(_T_205),
        .b(_T_176)
    );
    wire [63:0] _T_208;
    BITS #(.width(129), .high(63), .low(0)) bits_4529 (
        .y(_T_208),
        .in(_T_207)
    );
    wire [128:0] _T_209;
    CAT #(.width_a(65), .width_b(64)) cat_4530 (
        .y(_T_209),
        .a(_T_206),
        .b(_T_208)
    );
    wire [64:0] _T_210;
    SHR_UNSIGNED #(.width(129), .n(64)) u_shr_4531 (
        .y(_T_210),
        .in(_T_209)
    );
    wire [63:0] _T_212;
    BITS #(.width(129), .high(63), .low(0)) bits_4532 (
        .y(_T_212),
        .in(_T_209)
    );
    wire [65:0] _T_213;
    CAT #(.width_a(65), .width_b(1)) cat_4533 (
        .y(_T_213),
        .a(_T_210),
        .b(1'h0)
    );
    wire [129:0] _T_214;
    CAT #(.width_a(66), .width_b(64)) cat_4534 (
        .y(_T_214),
        .a(_T_213),
        .b(_T_212)
    );
    wire [7:0] _T_216;
    wire [6:0] _WTEMP_623;
    PAD_UNSIGNED #(.width(1), .n(7)) u_pad_4535 (
        .y(_WTEMP_623),
        .in(1'h1)
    );
    ADD_UNSIGNED #(.width(7)) u_add_4536 (
        .y(_T_216),
        .a(_count__q),
        .b(_WTEMP_623)
    );
    wire [6:0] _T_217;
    TAIL #(.width(8), .n(1)) tail_4537 (
        .y(_T_217),
        .in(_T_216)
    );
    wire _T_219;
    wire [6:0] _WTEMP_624;
    PAD_UNSIGNED #(.width(3), .n(7)) u_pad_4538 (
        .y(_WTEMP_624),
        .in(3'h7)
    );
    EQ_UNSIGNED #(.width(7)) u_eq_4539 (
        .y(_T_219),
        .a(_count__q),
        .b(_WTEMP_624)
    );
    wire _T_220;
    BITWISEOR #(.width(1)) bitwiseor_4540 (
        .y(_T_220),
        .a(_T_197),
        .b(_T_219)
    );
    wire [2:0] _T_221;
    MUX_UNSIGNED #(.width(3)) u_mux_4541 (
        .y(_T_221),
        .sel(_isHi__q),
        .a(3'h3),
        .b(3'h5)
    );
    wire [2:0] _node_346;
    MUX_UNSIGNED #(.width(3)) u_mux_4542 (
        .y(_node_346),
        .sel(_T_157),
        .a(_T_159),
        .b(_node_345)
    );
    wire [129:0] _node_347;
    wire [129:0] _WTEMP_625;
    PAD_UNSIGNED #(.width(64), .n(130)) u_pad_4543 (
        .y(_WTEMP_625),
        .in(_T_158)
    );
    MUX_UNSIGNED #(.width(130)) u_mux_4544 (
        .y(_node_347),
        .sel(_T_157),
        .a(_WTEMP_625),
        .b(_node_344)
    );
    wire [2:0] _node_348;
    MUX_UNSIGNED #(.width(3)) u_mux_4545 (
        .y(_node_348),
        .sel(_T_220),
        .a(_T_221),
        .b(_node_346)
    );
    wire [2:0] _node_349;
    MUX_UNSIGNED #(.width(3)) u_mux_4546 (
        .y(_node_349),
        .sel(_T_157),
        .a(_T_159),
        .b(_node_345)
    );
    wire _T_222;
    EQ_UNSIGNED #(.width(3)) u_eq_4547 (
        .y(_T_222),
        .a(_state__q),
        .b(3'h2)
    );
    wire _T_224;
    EQ_UNSIGNED #(.width(1)) u_eq_4548 (
        .y(_T_224),
        .a(_isMul__q),
        .b(1'h0)
    );
    wire _T_225;
    BITWISEAND #(.width(1)) bitwiseand_4549 (
        .y(_T_225),
        .a(_T_222),
        .b(_T_224)
    );
    wire _T_226;
    BITS #(.width(65), .high(64), .low(64)) bits_4550 (
        .y(_T_226),
        .in(subtractor)
    );
    wire [63:0] _T_227;
    BITS #(.width(130), .high(127), .low(64)) bits_4551 (
        .y(_T_227),
        .in(_remainder__q)
    );
    wire [63:0] _T_228;
    BITS #(.width(65), .high(63), .low(0)) bits_4552 (
        .y(_T_228),
        .in(subtractor)
    );
    wire [63:0] _T_229;
    MUX_UNSIGNED #(.width(64)) u_mux_4553 (
        .y(_T_229),
        .sel(_T_226),
        .a(_T_227),
        .b(_T_228)
    );
    wire [63:0] _T_230;
    BITS #(.width(130), .high(63), .low(0)) bits_4554 (
        .y(_T_230),
        .in(_remainder__q)
    );
    wire _T_232;
    EQ_UNSIGNED #(.width(1)) u_eq_4555 (
        .y(_T_232),
        .a(_T_226),
        .b(1'h0)
    );
    wire [127:0] _T_233;
    CAT #(.width_a(64), .width_b(64)) cat_4556 (
        .y(_T_233),
        .a(_T_229),
        .b(_T_230)
    );
    wire [128:0] _T_234;
    CAT #(.width_a(128), .width_b(1)) cat_4557 (
        .y(_T_234),
        .a(_T_233),
        .b(_T_232)
    );
    wire _T_236;
    EQ_UNSIGNED #(.width(7)) u_eq_4558 (
        .y(_T_236),
        .a(_count__q),
        .b(7'h40)
    );
    wire [2:0] _T_237;
    MUX_UNSIGNED #(.width(3)) u_mux_4559 (
        .y(_T_237),
        .sel(_neg_out__q),
        .a(3'h4),
        .b(3'h5)
    );
    wire [2:0] _T_238;
    MUX_UNSIGNED #(.width(3)) u_mux_4560 (
        .y(_T_238),
        .sel(_isHi__q),
        .a(3'h3),
        .b(_T_237)
    );
    wire [2:0] _node_350;
    MUX_UNSIGNED #(.width(3)) u_mux_4561 (
        .y(_node_350),
        .sel(_T_161),
        .a(_node_348),
        .b(_node_349)
    );
    wire [7:0] _T_240;
    wire [6:0] _WTEMP_626;
    PAD_UNSIGNED #(.width(1), .n(7)) u_pad_4562 (
        .y(_WTEMP_626),
        .in(1'h1)
    );
    ADD_UNSIGNED #(.width(7)) u_add_4563 (
        .y(_T_240),
        .a(_count__q),
        .b(_WTEMP_626)
    );
    wire [6:0] _T_241;
    TAIL #(.width(8), .n(1)) tail_4564 (
        .y(_T_241),
        .in(_T_240)
    );
    wire _T_243;
    wire [6:0] _WTEMP_627;
    PAD_UNSIGNED #(.width(1), .n(7)) u_pad_4565 (
        .y(_WTEMP_627),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(7)) u_eq_4566 (
        .y(_T_243),
        .a(_count__q),
        .b(_WTEMP_627)
    );
    wire _T_244;
    BITS #(.width(65), .high(64), .low(64)) bits_4567 (
        .y(_T_244),
        .in(subtractor)
    );
    wire _T_246;
    EQ_UNSIGNED #(.width(1)) u_eq_4568 (
        .y(_T_246),
        .a(_T_244),
        .b(1'h0)
    );
    wire _T_247;
    BITWISEAND #(.width(1)) bitwiseand_4569 (
        .y(_T_247),
        .a(_T_243),
        .b(_T_246)
    );
    wire [63:0] _T_248;
    BITS #(.width(65), .high(63), .low(0)) bits_4570 (
        .y(_T_248),
        .in(_divisor__q)
    );
    wire [31:0] _T_249;
    BITS #(.width(64), .high(63), .low(32)) bits_4571 (
        .y(_T_249),
        .in(_T_248)
    );
    wire [31:0] _T_250;
    BITS #(.width(64), .high(31), .low(0)) bits_4572 (
        .y(_T_250),
        .in(_T_248)
    );
    wire _T_252;
    wire [31:0] _WTEMP_628;
    PAD_UNSIGNED #(.width(1), .n(32)) u_pad_4573 (
        .y(_WTEMP_628),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(32)) u_neq_4574 (
        .y(_T_252),
        .a(_T_249),
        .b(_WTEMP_628)
    );
    wire [15:0] _T_253;
    BITS #(.width(32), .high(31), .low(16)) bits_4575 (
        .y(_T_253),
        .in(_T_249)
    );
    wire [15:0] _T_254;
    BITS #(.width(32), .high(15), .low(0)) bits_4576 (
        .y(_T_254),
        .in(_T_249)
    );
    wire _T_256;
    wire [15:0] _WTEMP_629;
    PAD_UNSIGNED #(.width(1), .n(16)) u_pad_4577 (
        .y(_WTEMP_629),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(16)) u_neq_4578 (
        .y(_T_256),
        .a(_T_253),
        .b(_WTEMP_629)
    );
    wire [7:0] _T_257;
    BITS #(.width(16), .high(15), .low(8)) bits_4579 (
        .y(_T_257),
        .in(_T_253)
    );
    wire [7:0] _T_258;
    BITS #(.width(16), .high(7), .low(0)) bits_4580 (
        .y(_T_258),
        .in(_T_253)
    );
    wire _T_260;
    wire [7:0] _WTEMP_630;
    PAD_UNSIGNED #(.width(1), .n(8)) u_pad_4581 (
        .y(_WTEMP_630),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(8)) u_neq_4582 (
        .y(_T_260),
        .a(_T_257),
        .b(_WTEMP_630)
    );
    wire [3:0] _T_261;
    BITS #(.width(8), .high(7), .low(4)) bits_4583 (
        .y(_T_261),
        .in(_T_257)
    );
    wire [3:0] _T_262;
    BITS #(.width(8), .high(3), .low(0)) bits_4584 (
        .y(_T_262),
        .in(_T_257)
    );
    wire _T_264;
    wire [3:0] _WTEMP_631;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_4585 (
        .y(_WTEMP_631),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_4586 (
        .y(_T_264),
        .a(_T_261),
        .b(_WTEMP_631)
    );
    wire _T_265;
    BITS #(.width(4), .high(3), .low(3)) bits_4587 (
        .y(_T_265),
        .in(_T_261)
    );
    wire _T_267;
    BITS #(.width(4), .high(2), .low(2)) bits_4588 (
        .y(_T_267),
        .in(_T_261)
    );
    wire _T_269;
    BITS #(.width(4), .high(1), .low(1)) bits_4589 (
        .y(_T_269),
        .in(_T_261)
    );
    wire [1:0] _T_270;
    wire [1:0] _WTEMP_632;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_4590 (
        .y(_WTEMP_632),
        .in(_T_269)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_4591 (
        .y(_T_270),
        .sel(_T_267),
        .a(2'h2),
        .b(_WTEMP_632)
    );
    wire [1:0] _T_271;
    MUX_UNSIGNED #(.width(2)) u_mux_4592 (
        .y(_T_271),
        .sel(_T_265),
        .a(2'h3),
        .b(_T_270)
    );
    wire _T_272;
    BITS #(.width(4), .high(3), .low(3)) bits_4593 (
        .y(_T_272),
        .in(_T_262)
    );
    wire _T_274;
    BITS #(.width(4), .high(2), .low(2)) bits_4594 (
        .y(_T_274),
        .in(_T_262)
    );
    wire _T_276;
    BITS #(.width(4), .high(1), .low(1)) bits_4595 (
        .y(_T_276),
        .in(_T_262)
    );
    wire [1:0] _T_277;
    wire [1:0] _WTEMP_633;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_4596 (
        .y(_WTEMP_633),
        .in(_T_276)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_4597 (
        .y(_T_277),
        .sel(_T_274),
        .a(2'h2),
        .b(_WTEMP_633)
    );
    wire [1:0] _T_278;
    MUX_UNSIGNED #(.width(2)) u_mux_4598 (
        .y(_T_278),
        .sel(_T_272),
        .a(2'h3),
        .b(_T_277)
    );
    wire [1:0] _T_279;
    MUX_UNSIGNED #(.width(2)) u_mux_4599 (
        .y(_T_279),
        .sel(_T_264),
        .a(_T_271),
        .b(_T_278)
    );
    wire [2:0] _T_280;
    CAT #(.width_a(1), .width_b(2)) cat_4600 (
        .y(_T_280),
        .a(_T_264),
        .b(_T_279)
    );
    wire [3:0] _T_281;
    BITS #(.width(8), .high(7), .low(4)) bits_4601 (
        .y(_T_281),
        .in(_T_258)
    );
    wire [3:0] _T_282;
    BITS #(.width(8), .high(3), .low(0)) bits_4602 (
        .y(_T_282),
        .in(_T_258)
    );
    wire _T_284;
    wire [3:0] _WTEMP_634;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_4603 (
        .y(_WTEMP_634),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_4604 (
        .y(_T_284),
        .a(_T_281),
        .b(_WTEMP_634)
    );
    wire _T_285;
    BITS #(.width(4), .high(3), .low(3)) bits_4605 (
        .y(_T_285),
        .in(_T_281)
    );
    wire _T_287;
    BITS #(.width(4), .high(2), .low(2)) bits_4606 (
        .y(_T_287),
        .in(_T_281)
    );
    wire _T_289;
    BITS #(.width(4), .high(1), .low(1)) bits_4607 (
        .y(_T_289),
        .in(_T_281)
    );
    wire [1:0] _T_290;
    wire [1:0] _WTEMP_635;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_4608 (
        .y(_WTEMP_635),
        .in(_T_289)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_4609 (
        .y(_T_290),
        .sel(_T_287),
        .a(2'h2),
        .b(_WTEMP_635)
    );
    wire [1:0] _T_291;
    MUX_UNSIGNED #(.width(2)) u_mux_4610 (
        .y(_T_291),
        .sel(_T_285),
        .a(2'h3),
        .b(_T_290)
    );
    wire _T_292;
    BITS #(.width(4), .high(3), .low(3)) bits_4611 (
        .y(_T_292),
        .in(_T_282)
    );
    wire _T_294;
    BITS #(.width(4), .high(2), .low(2)) bits_4612 (
        .y(_T_294),
        .in(_T_282)
    );
    wire _T_296;
    BITS #(.width(4), .high(1), .low(1)) bits_4613 (
        .y(_T_296),
        .in(_T_282)
    );
    wire [1:0] _T_297;
    wire [1:0] _WTEMP_636;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_4614 (
        .y(_WTEMP_636),
        .in(_T_296)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_4615 (
        .y(_T_297),
        .sel(_T_294),
        .a(2'h2),
        .b(_WTEMP_636)
    );
    wire [1:0] _T_298;
    MUX_UNSIGNED #(.width(2)) u_mux_4616 (
        .y(_T_298),
        .sel(_T_292),
        .a(2'h3),
        .b(_T_297)
    );
    wire [1:0] _T_299;
    MUX_UNSIGNED #(.width(2)) u_mux_4617 (
        .y(_T_299),
        .sel(_T_284),
        .a(_T_291),
        .b(_T_298)
    );
    wire [2:0] _T_300;
    CAT #(.width_a(1), .width_b(2)) cat_4618 (
        .y(_T_300),
        .a(_T_284),
        .b(_T_299)
    );
    wire [2:0] _T_301;
    MUX_UNSIGNED #(.width(3)) u_mux_4619 (
        .y(_T_301),
        .sel(_T_260),
        .a(_T_280),
        .b(_T_300)
    );
    wire [3:0] _T_302;
    CAT #(.width_a(1), .width_b(3)) cat_4620 (
        .y(_T_302),
        .a(_T_260),
        .b(_T_301)
    );
    wire [7:0] _T_303;
    BITS #(.width(16), .high(15), .low(8)) bits_4621 (
        .y(_T_303),
        .in(_T_254)
    );
    wire [7:0] _T_304;
    BITS #(.width(16), .high(7), .low(0)) bits_4622 (
        .y(_T_304),
        .in(_T_254)
    );
    wire _T_306;
    wire [7:0] _WTEMP_637;
    PAD_UNSIGNED #(.width(1), .n(8)) u_pad_4623 (
        .y(_WTEMP_637),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(8)) u_neq_4624 (
        .y(_T_306),
        .a(_T_303),
        .b(_WTEMP_637)
    );
    wire [3:0] _T_307;
    BITS #(.width(8), .high(7), .low(4)) bits_4625 (
        .y(_T_307),
        .in(_T_303)
    );
    wire [3:0] _T_308;
    BITS #(.width(8), .high(3), .low(0)) bits_4626 (
        .y(_T_308),
        .in(_T_303)
    );
    wire _T_310;
    wire [3:0] _WTEMP_638;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_4627 (
        .y(_WTEMP_638),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_4628 (
        .y(_T_310),
        .a(_T_307),
        .b(_WTEMP_638)
    );
    wire _T_311;
    BITS #(.width(4), .high(3), .low(3)) bits_4629 (
        .y(_T_311),
        .in(_T_307)
    );
    wire _T_313;
    BITS #(.width(4), .high(2), .low(2)) bits_4630 (
        .y(_T_313),
        .in(_T_307)
    );
    wire _T_315;
    BITS #(.width(4), .high(1), .low(1)) bits_4631 (
        .y(_T_315),
        .in(_T_307)
    );
    wire [1:0] _T_316;
    wire [1:0] _WTEMP_639;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_4632 (
        .y(_WTEMP_639),
        .in(_T_315)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_4633 (
        .y(_T_316),
        .sel(_T_313),
        .a(2'h2),
        .b(_WTEMP_639)
    );
    wire [1:0] _T_317;
    MUX_UNSIGNED #(.width(2)) u_mux_4634 (
        .y(_T_317),
        .sel(_T_311),
        .a(2'h3),
        .b(_T_316)
    );
    wire _T_318;
    BITS #(.width(4), .high(3), .low(3)) bits_4635 (
        .y(_T_318),
        .in(_T_308)
    );
    wire _T_320;
    BITS #(.width(4), .high(2), .low(2)) bits_4636 (
        .y(_T_320),
        .in(_T_308)
    );
    wire _T_322;
    BITS #(.width(4), .high(1), .low(1)) bits_4637 (
        .y(_T_322),
        .in(_T_308)
    );
    wire [1:0] _T_323;
    wire [1:0] _WTEMP_640;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_4638 (
        .y(_WTEMP_640),
        .in(_T_322)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_4639 (
        .y(_T_323),
        .sel(_T_320),
        .a(2'h2),
        .b(_WTEMP_640)
    );
    wire [1:0] _T_324;
    MUX_UNSIGNED #(.width(2)) u_mux_4640 (
        .y(_T_324),
        .sel(_T_318),
        .a(2'h3),
        .b(_T_323)
    );
    wire [1:0] _T_325;
    MUX_UNSIGNED #(.width(2)) u_mux_4641 (
        .y(_T_325),
        .sel(_T_310),
        .a(_T_317),
        .b(_T_324)
    );
    wire [2:0] _T_326;
    CAT #(.width_a(1), .width_b(2)) cat_4642 (
        .y(_T_326),
        .a(_T_310),
        .b(_T_325)
    );
    wire [3:0] _T_327;
    BITS #(.width(8), .high(7), .low(4)) bits_4643 (
        .y(_T_327),
        .in(_T_304)
    );
    wire [3:0] _T_328;
    BITS #(.width(8), .high(3), .low(0)) bits_4644 (
        .y(_T_328),
        .in(_T_304)
    );
    wire _T_330;
    wire [3:0] _WTEMP_641;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_4645 (
        .y(_WTEMP_641),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_4646 (
        .y(_T_330),
        .a(_T_327),
        .b(_WTEMP_641)
    );
    wire _T_331;
    BITS #(.width(4), .high(3), .low(3)) bits_4647 (
        .y(_T_331),
        .in(_T_327)
    );
    wire _T_333;
    BITS #(.width(4), .high(2), .low(2)) bits_4648 (
        .y(_T_333),
        .in(_T_327)
    );
    wire _T_335;
    BITS #(.width(4), .high(1), .low(1)) bits_4649 (
        .y(_T_335),
        .in(_T_327)
    );
    wire [1:0] _T_336;
    wire [1:0] _WTEMP_642;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_4650 (
        .y(_WTEMP_642),
        .in(_T_335)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_4651 (
        .y(_T_336),
        .sel(_T_333),
        .a(2'h2),
        .b(_WTEMP_642)
    );
    wire [1:0] _T_337;
    MUX_UNSIGNED #(.width(2)) u_mux_4652 (
        .y(_T_337),
        .sel(_T_331),
        .a(2'h3),
        .b(_T_336)
    );
    wire _T_338;
    BITS #(.width(4), .high(3), .low(3)) bits_4653 (
        .y(_T_338),
        .in(_T_328)
    );
    wire _T_340;
    BITS #(.width(4), .high(2), .low(2)) bits_4654 (
        .y(_T_340),
        .in(_T_328)
    );
    wire _T_342;
    BITS #(.width(4), .high(1), .low(1)) bits_4655 (
        .y(_T_342),
        .in(_T_328)
    );
    wire [1:0] _T_343;
    wire [1:0] _WTEMP_643;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_4656 (
        .y(_WTEMP_643),
        .in(_T_342)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_4657 (
        .y(_T_343),
        .sel(_T_340),
        .a(2'h2),
        .b(_WTEMP_643)
    );
    wire [1:0] _T_344;
    MUX_UNSIGNED #(.width(2)) u_mux_4658 (
        .y(_T_344),
        .sel(_T_338),
        .a(2'h3),
        .b(_T_343)
    );
    wire [1:0] _T_345;
    MUX_UNSIGNED #(.width(2)) u_mux_4659 (
        .y(_T_345),
        .sel(_T_330),
        .a(_T_337),
        .b(_T_344)
    );
    wire [2:0] _T_346;
    CAT #(.width_a(1), .width_b(2)) cat_4660 (
        .y(_T_346),
        .a(_T_330),
        .b(_T_345)
    );
    wire [2:0] _T_347;
    MUX_UNSIGNED #(.width(3)) u_mux_4661 (
        .y(_T_347),
        .sel(_T_306),
        .a(_T_326),
        .b(_T_346)
    );
    wire [3:0] _T_348;
    CAT #(.width_a(1), .width_b(3)) cat_4662 (
        .y(_T_348),
        .a(_T_306),
        .b(_T_347)
    );
    wire [3:0] _T_349;
    MUX_UNSIGNED #(.width(4)) u_mux_4663 (
        .y(_T_349),
        .sel(_T_256),
        .a(_T_302),
        .b(_T_348)
    );
    wire [4:0] _T_350;
    CAT #(.width_a(1), .width_b(4)) cat_4664 (
        .y(_T_350),
        .a(_T_256),
        .b(_T_349)
    );
    wire [15:0] _T_351;
    BITS #(.width(32), .high(31), .low(16)) bits_4665 (
        .y(_T_351),
        .in(_T_250)
    );
    wire [15:0] _T_352;
    BITS #(.width(32), .high(15), .low(0)) bits_4666 (
        .y(_T_352),
        .in(_T_250)
    );
    wire _T_354;
    wire [15:0] _WTEMP_644;
    PAD_UNSIGNED #(.width(1), .n(16)) u_pad_4667 (
        .y(_WTEMP_644),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(16)) u_neq_4668 (
        .y(_T_354),
        .a(_T_351),
        .b(_WTEMP_644)
    );
    wire [7:0] _T_355;
    BITS #(.width(16), .high(15), .low(8)) bits_4669 (
        .y(_T_355),
        .in(_T_351)
    );
    wire [7:0] _T_356;
    BITS #(.width(16), .high(7), .low(0)) bits_4670 (
        .y(_T_356),
        .in(_T_351)
    );
    wire _T_358;
    wire [7:0] _WTEMP_645;
    PAD_UNSIGNED #(.width(1), .n(8)) u_pad_4671 (
        .y(_WTEMP_645),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(8)) u_neq_4672 (
        .y(_T_358),
        .a(_T_355),
        .b(_WTEMP_645)
    );
    wire [3:0] _T_359;
    BITS #(.width(8), .high(7), .low(4)) bits_4673 (
        .y(_T_359),
        .in(_T_355)
    );
    wire [3:0] _T_360;
    BITS #(.width(8), .high(3), .low(0)) bits_4674 (
        .y(_T_360),
        .in(_T_355)
    );
    wire _T_362;
    wire [3:0] _WTEMP_646;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_4675 (
        .y(_WTEMP_646),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_4676 (
        .y(_T_362),
        .a(_T_359),
        .b(_WTEMP_646)
    );
    wire _T_363;
    BITS #(.width(4), .high(3), .low(3)) bits_4677 (
        .y(_T_363),
        .in(_T_359)
    );
    wire _T_365;
    BITS #(.width(4), .high(2), .low(2)) bits_4678 (
        .y(_T_365),
        .in(_T_359)
    );
    wire _T_367;
    BITS #(.width(4), .high(1), .low(1)) bits_4679 (
        .y(_T_367),
        .in(_T_359)
    );
    wire [1:0] _T_368;
    wire [1:0] _WTEMP_647;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_4680 (
        .y(_WTEMP_647),
        .in(_T_367)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_4681 (
        .y(_T_368),
        .sel(_T_365),
        .a(2'h2),
        .b(_WTEMP_647)
    );
    wire [1:0] _T_369;
    MUX_UNSIGNED #(.width(2)) u_mux_4682 (
        .y(_T_369),
        .sel(_T_363),
        .a(2'h3),
        .b(_T_368)
    );
    wire _T_370;
    BITS #(.width(4), .high(3), .low(3)) bits_4683 (
        .y(_T_370),
        .in(_T_360)
    );
    wire _T_372;
    BITS #(.width(4), .high(2), .low(2)) bits_4684 (
        .y(_T_372),
        .in(_T_360)
    );
    wire _T_374;
    BITS #(.width(4), .high(1), .low(1)) bits_4685 (
        .y(_T_374),
        .in(_T_360)
    );
    wire [1:0] _T_375;
    wire [1:0] _WTEMP_648;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_4686 (
        .y(_WTEMP_648),
        .in(_T_374)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_4687 (
        .y(_T_375),
        .sel(_T_372),
        .a(2'h2),
        .b(_WTEMP_648)
    );
    wire [1:0] _T_376;
    MUX_UNSIGNED #(.width(2)) u_mux_4688 (
        .y(_T_376),
        .sel(_T_370),
        .a(2'h3),
        .b(_T_375)
    );
    wire [1:0] _T_377;
    MUX_UNSIGNED #(.width(2)) u_mux_4689 (
        .y(_T_377),
        .sel(_T_362),
        .a(_T_369),
        .b(_T_376)
    );
    wire [2:0] _T_378;
    CAT #(.width_a(1), .width_b(2)) cat_4690 (
        .y(_T_378),
        .a(_T_362),
        .b(_T_377)
    );
    wire [3:0] _T_379;
    BITS #(.width(8), .high(7), .low(4)) bits_4691 (
        .y(_T_379),
        .in(_T_356)
    );
    wire [3:0] _T_380;
    BITS #(.width(8), .high(3), .low(0)) bits_4692 (
        .y(_T_380),
        .in(_T_356)
    );
    wire _T_382;
    wire [3:0] _WTEMP_649;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_4693 (
        .y(_WTEMP_649),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_4694 (
        .y(_T_382),
        .a(_T_379),
        .b(_WTEMP_649)
    );
    wire _T_383;
    BITS #(.width(4), .high(3), .low(3)) bits_4695 (
        .y(_T_383),
        .in(_T_379)
    );
    wire _T_385;
    BITS #(.width(4), .high(2), .low(2)) bits_4696 (
        .y(_T_385),
        .in(_T_379)
    );
    wire _T_387;
    BITS #(.width(4), .high(1), .low(1)) bits_4697 (
        .y(_T_387),
        .in(_T_379)
    );
    wire [1:0] _T_388;
    wire [1:0] _WTEMP_650;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_4698 (
        .y(_WTEMP_650),
        .in(_T_387)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_4699 (
        .y(_T_388),
        .sel(_T_385),
        .a(2'h2),
        .b(_WTEMP_650)
    );
    wire [1:0] _T_389;
    MUX_UNSIGNED #(.width(2)) u_mux_4700 (
        .y(_T_389),
        .sel(_T_383),
        .a(2'h3),
        .b(_T_388)
    );
    wire _T_390;
    BITS #(.width(4), .high(3), .low(3)) bits_4701 (
        .y(_T_390),
        .in(_T_380)
    );
    wire _T_392;
    BITS #(.width(4), .high(2), .low(2)) bits_4702 (
        .y(_T_392),
        .in(_T_380)
    );
    wire _T_394;
    BITS #(.width(4), .high(1), .low(1)) bits_4703 (
        .y(_T_394),
        .in(_T_380)
    );
    wire [1:0] _T_395;
    wire [1:0] _WTEMP_651;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_4704 (
        .y(_WTEMP_651),
        .in(_T_394)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_4705 (
        .y(_T_395),
        .sel(_T_392),
        .a(2'h2),
        .b(_WTEMP_651)
    );
    wire [1:0] _T_396;
    MUX_UNSIGNED #(.width(2)) u_mux_4706 (
        .y(_T_396),
        .sel(_T_390),
        .a(2'h3),
        .b(_T_395)
    );
    wire [1:0] _T_397;
    MUX_UNSIGNED #(.width(2)) u_mux_4707 (
        .y(_T_397),
        .sel(_T_382),
        .a(_T_389),
        .b(_T_396)
    );
    wire [2:0] _T_398;
    CAT #(.width_a(1), .width_b(2)) cat_4708 (
        .y(_T_398),
        .a(_T_382),
        .b(_T_397)
    );
    wire [2:0] _T_399;
    MUX_UNSIGNED #(.width(3)) u_mux_4709 (
        .y(_T_399),
        .sel(_T_358),
        .a(_T_378),
        .b(_T_398)
    );
    wire [3:0] _T_400;
    CAT #(.width_a(1), .width_b(3)) cat_4710 (
        .y(_T_400),
        .a(_T_358),
        .b(_T_399)
    );
    wire [7:0] _T_401;
    BITS #(.width(16), .high(15), .low(8)) bits_4711 (
        .y(_T_401),
        .in(_T_352)
    );
    wire [7:0] _T_402;
    BITS #(.width(16), .high(7), .low(0)) bits_4712 (
        .y(_T_402),
        .in(_T_352)
    );
    wire _T_404;
    wire [7:0] _WTEMP_652;
    PAD_UNSIGNED #(.width(1), .n(8)) u_pad_4713 (
        .y(_WTEMP_652),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(8)) u_neq_4714 (
        .y(_T_404),
        .a(_T_401),
        .b(_WTEMP_652)
    );
    wire [3:0] _T_405;
    BITS #(.width(8), .high(7), .low(4)) bits_4715 (
        .y(_T_405),
        .in(_T_401)
    );
    wire [3:0] _T_406;
    BITS #(.width(8), .high(3), .low(0)) bits_4716 (
        .y(_T_406),
        .in(_T_401)
    );
    wire _T_408;
    wire [3:0] _WTEMP_653;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_4717 (
        .y(_WTEMP_653),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_4718 (
        .y(_T_408),
        .a(_T_405),
        .b(_WTEMP_653)
    );
    wire _T_409;
    BITS #(.width(4), .high(3), .low(3)) bits_4719 (
        .y(_T_409),
        .in(_T_405)
    );
    wire _T_411;
    BITS #(.width(4), .high(2), .low(2)) bits_4720 (
        .y(_T_411),
        .in(_T_405)
    );
    wire _T_413;
    BITS #(.width(4), .high(1), .low(1)) bits_4721 (
        .y(_T_413),
        .in(_T_405)
    );
    wire [1:0] _T_414;
    wire [1:0] _WTEMP_654;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_4722 (
        .y(_WTEMP_654),
        .in(_T_413)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_4723 (
        .y(_T_414),
        .sel(_T_411),
        .a(2'h2),
        .b(_WTEMP_654)
    );
    wire [1:0] _T_415;
    MUX_UNSIGNED #(.width(2)) u_mux_4724 (
        .y(_T_415),
        .sel(_T_409),
        .a(2'h3),
        .b(_T_414)
    );
    wire _T_416;
    BITS #(.width(4), .high(3), .low(3)) bits_4725 (
        .y(_T_416),
        .in(_T_406)
    );
    wire _T_418;
    BITS #(.width(4), .high(2), .low(2)) bits_4726 (
        .y(_T_418),
        .in(_T_406)
    );
    wire _T_420;
    BITS #(.width(4), .high(1), .low(1)) bits_4727 (
        .y(_T_420),
        .in(_T_406)
    );
    wire [1:0] _T_421;
    wire [1:0] _WTEMP_655;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_4728 (
        .y(_WTEMP_655),
        .in(_T_420)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_4729 (
        .y(_T_421),
        .sel(_T_418),
        .a(2'h2),
        .b(_WTEMP_655)
    );
    wire [1:0] _T_422;
    MUX_UNSIGNED #(.width(2)) u_mux_4730 (
        .y(_T_422),
        .sel(_T_416),
        .a(2'h3),
        .b(_T_421)
    );
    wire [1:0] _T_423;
    MUX_UNSIGNED #(.width(2)) u_mux_4731 (
        .y(_T_423),
        .sel(_T_408),
        .a(_T_415),
        .b(_T_422)
    );
    wire [2:0] _T_424;
    CAT #(.width_a(1), .width_b(2)) cat_4732 (
        .y(_T_424),
        .a(_T_408),
        .b(_T_423)
    );
    wire [3:0] _T_425;
    BITS #(.width(8), .high(7), .low(4)) bits_4733 (
        .y(_T_425),
        .in(_T_402)
    );
    wire [3:0] _T_426;
    BITS #(.width(8), .high(3), .low(0)) bits_4734 (
        .y(_T_426),
        .in(_T_402)
    );
    wire _T_428;
    wire [3:0] _WTEMP_656;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_4735 (
        .y(_WTEMP_656),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_4736 (
        .y(_T_428),
        .a(_T_425),
        .b(_WTEMP_656)
    );
    wire _T_429;
    BITS #(.width(4), .high(3), .low(3)) bits_4737 (
        .y(_T_429),
        .in(_T_425)
    );
    wire _T_431;
    BITS #(.width(4), .high(2), .low(2)) bits_4738 (
        .y(_T_431),
        .in(_T_425)
    );
    wire _T_433;
    BITS #(.width(4), .high(1), .low(1)) bits_4739 (
        .y(_T_433),
        .in(_T_425)
    );
    wire [1:0] _T_434;
    wire [1:0] _WTEMP_657;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_4740 (
        .y(_WTEMP_657),
        .in(_T_433)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_4741 (
        .y(_T_434),
        .sel(_T_431),
        .a(2'h2),
        .b(_WTEMP_657)
    );
    wire [1:0] _T_435;
    MUX_UNSIGNED #(.width(2)) u_mux_4742 (
        .y(_T_435),
        .sel(_T_429),
        .a(2'h3),
        .b(_T_434)
    );
    wire _T_436;
    BITS #(.width(4), .high(3), .low(3)) bits_4743 (
        .y(_T_436),
        .in(_T_426)
    );
    wire _T_438;
    BITS #(.width(4), .high(2), .low(2)) bits_4744 (
        .y(_T_438),
        .in(_T_426)
    );
    wire _T_440;
    BITS #(.width(4), .high(1), .low(1)) bits_4745 (
        .y(_T_440),
        .in(_T_426)
    );
    wire [1:0] _T_441;
    wire [1:0] _WTEMP_658;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_4746 (
        .y(_WTEMP_658),
        .in(_T_440)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_4747 (
        .y(_T_441),
        .sel(_T_438),
        .a(2'h2),
        .b(_WTEMP_658)
    );
    wire [1:0] _T_442;
    MUX_UNSIGNED #(.width(2)) u_mux_4748 (
        .y(_T_442),
        .sel(_T_436),
        .a(2'h3),
        .b(_T_441)
    );
    wire [1:0] _T_443;
    MUX_UNSIGNED #(.width(2)) u_mux_4749 (
        .y(_T_443),
        .sel(_T_428),
        .a(_T_435),
        .b(_T_442)
    );
    wire [2:0] _T_444;
    CAT #(.width_a(1), .width_b(2)) cat_4750 (
        .y(_T_444),
        .a(_T_428),
        .b(_T_443)
    );
    wire [2:0] _T_445;
    MUX_UNSIGNED #(.width(3)) u_mux_4751 (
        .y(_T_445),
        .sel(_T_404),
        .a(_T_424),
        .b(_T_444)
    );
    wire [3:0] _T_446;
    CAT #(.width_a(1), .width_b(3)) cat_4752 (
        .y(_T_446),
        .a(_T_404),
        .b(_T_445)
    );
    wire [3:0] _T_447;
    MUX_UNSIGNED #(.width(4)) u_mux_4753 (
        .y(_T_447),
        .sel(_T_354),
        .a(_T_400),
        .b(_T_446)
    );
    wire [4:0] _T_448;
    CAT #(.width_a(1), .width_b(4)) cat_4754 (
        .y(_T_448),
        .a(_T_354),
        .b(_T_447)
    );
    wire [4:0] _T_449;
    MUX_UNSIGNED #(.width(5)) u_mux_4755 (
        .y(_T_449),
        .sel(_T_252),
        .a(_T_350),
        .b(_T_448)
    );
    wire [5:0] _T_450;
    CAT #(.width_a(1), .width_b(5)) cat_4756 (
        .y(_T_450),
        .a(_T_252),
        .b(_T_449)
    );
    wire [63:0] _T_451;
    BITS #(.width(130), .high(63), .low(0)) bits_4757 (
        .y(_T_451),
        .in(_remainder__q)
    );
    wire [31:0] _T_452;
    BITS #(.width(64), .high(63), .low(32)) bits_4758 (
        .y(_T_452),
        .in(_T_451)
    );
    wire [31:0] _T_453;
    BITS #(.width(64), .high(31), .low(0)) bits_4759 (
        .y(_T_453),
        .in(_T_451)
    );
    wire _T_455;
    wire [31:0] _WTEMP_659;
    PAD_UNSIGNED #(.width(1), .n(32)) u_pad_4760 (
        .y(_WTEMP_659),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(32)) u_neq_4761 (
        .y(_T_455),
        .a(_T_452),
        .b(_WTEMP_659)
    );
    wire [15:0] _T_456;
    BITS #(.width(32), .high(31), .low(16)) bits_4762 (
        .y(_T_456),
        .in(_T_452)
    );
    wire [15:0] _T_457;
    BITS #(.width(32), .high(15), .low(0)) bits_4763 (
        .y(_T_457),
        .in(_T_452)
    );
    wire _T_459;
    wire [15:0] _WTEMP_660;
    PAD_UNSIGNED #(.width(1), .n(16)) u_pad_4764 (
        .y(_WTEMP_660),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(16)) u_neq_4765 (
        .y(_T_459),
        .a(_T_456),
        .b(_WTEMP_660)
    );
    wire [7:0] _T_460;
    BITS #(.width(16), .high(15), .low(8)) bits_4766 (
        .y(_T_460),
        .in(_T_456)
    );
    wire [7:0] _T_461;
    BITS #(.width(16), .high(7), .low(0)) bits_4767 (
        .y(_T_461),
        .in(_T_456)
    );
    wire _T_463;
    wire [7:0] _WTEMP_661;
    PAD_UNSIGNED #(.width(1), .n(8)) u_pad_4768 (
        .y(_WTEMP_661),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(8)) u_neq_4769 (
        .y(_T_463),
        .a(_T_460),
        .b(_WTEMP_661)
    );
    wire [3:0] _T_464;
    BITS #(.width(8), .high(7), .low(4)) bits_4770 (
        .y(_T_464),
        .in(_T_460)
    );
    wire [3:0] _T_465;
    BITS #(.width(8), .high(3), .low(0)) bits_4771 (
        .y(_T_465),
        .in(_T_460)
    );
    wire _T_467;
    wire [3:0] _WTEMP_662;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_4772 (
        .y(_WTEMP_662),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_4773 (
        .y(_T_467),
        .a(_T_464),
        .b(_WTEMP_662)
    );
    wire _T_468;
    BITS #(.width(4), .high(3), .low(3)) bits_4774 (
        .y(_T_468),
        .in(_T_464)
    );
    wire _T_470;
    BITS #(.width(4), .high(2), .low(2)) bits_4775 (
        .y(_T_470),
        .in(_T_464)
    );
    wire _T_472;
    BITS #(.width(4), .high(1), .low(1)) bits_4776 (
        .y(_T_472),
        .in(_T_464)
    );
    wire [1:0] _T_473;
    wire [1:0] _WTEMP_663;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_4777 (
        .y(_WTEMP_663),
        .in(_T_472)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_4778 (
        .y(_T_473),
        .sel(_T_470),
        .a(2'h2),
        .b(_WTEMP_663)
    );
    wire [1:0] _T_474;
    MUX_UNSIGNED #(.width(2)) u_mux_4779 (
        .y(_T_474),
        .sel(_T_468),
        .a(2'h3),
        .b(_T_473)
    );
    wire _T_475;
    BITS #(.width(4), .high(3), .low(3)) bits_4780 (
        .y(_T_475),
        .in(_T_465)
    );
    wire _T_477;
    BITS #(.width(4), .high(2), .low(2)) bits_4781 (
        .y(_T_477),
        .in(_T_465)
    );
    wire _T_479;
    BITS #(.width(4), .high(1), .low(1)) bits_4782 (
        .y(_T_479),
        .in(_T_465)
    );
    wire [1:0] _T_480;
    wire [1:0] _WTEMP_664;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_4783 (
        .y(_WTEMP_664),
        .in(_T_479)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_4784 (
        .y(_T_480),
        .sel(_T_477),
        .a(2'h2),
        .b(_WTEMP_664)
    );
    wire [1:0] _T_481;
    MUX_UNSIGNED #(.width(2)) u_mux_4785 (
        .y(_T_481),
        .sel(_T_475),
        .a(2'h3),
        .b(_T_480)
    );
    wire [1:0] _T_482;
    MUX_UNSIGNED #(.width(2)) u_mux_4786 (
        .y(_T_482),
        .sel(_T_467),
        .a(_T_474),
        .b(_T_481)
    );
    wire [2:0] _T_483;
    CAT #(.width_a(1), .width_b(2)) cat_4787 (
        .y(_T_483),
        .a(_T_467),
        .b(_T_482)
    );
    wire [3:0] _T_484;
    BITS #(.width(8), .high(7), .low(4)) bits_4788 (
        .y(_T_484),
        .in(_T_461)
    );
    wire [3:0] _T_485;
    BITS #(.width(8), .high(3), .low(0)) bits_4789 (
        .y(_T_485),
        .in(_T_461)
    );
    wire _T_487;
    wire [3:0] _WTEMP_665;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_4790 (
        .y(_WTEMP_665),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_4791 (
        .y(_T_487),
        .a(_T_484),
        .b(_WTEMP_665)
    );
    wire _T_488;
    BITS #(.width(4), .high(3), .low(3)) bits_4792 (
        .y(_T_488),
        .in(_T_484)
    );
    wire _T_490;
    BITS #(.width(4), .high(2), .low(2)) bits_4793 (
        .y(_T_490),
        .in(_T_484)
    );
    wire _T_492;
    BITS #(.width(4), .high(1), .low(1)) bits_4794 (
        .y(_T_492),
        .in(_T_484)
    );
    wire [1:0] _T_493;
    wire [1:0] _WTEMP_666;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_4795 (
        .y(_WTEMP_666),
        .in(_T_492)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_4796 (
        .y(_T_493),
        .sel(_T_490),
        .a(2'h2),
        .b(_WTEMP_666)
    );
    wire [1:0] _T_494;
    MUX_UNSIGNED #(.width(2)) u_mux_4797 (
        .y(_T_494),
        .sel(_T_488),
        .a(2'h3),
        .b(_T_493)
    );
    wire _T_495;
    BITS #(.width(4), .high(3), .low(3)) bits_4798 (
        .y(_T_495),
        .in(_T_485)
    );
    wire _T_497;
    BITS #(.width(4), .high(2), .low(2)) bits_4799 (
        .y(_T_497),
        .in(_T_485)
    );
    wire _T_499;
    BITS #(.width(4), .high(1), .low(1)) bits_4800 (
        .y(_T_499),
        .in(_T_485)
    );
    wire [1:0] _T_500;
    wire [1:0] _WTEMP_667;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_4801 (
        .y(_WTEMP_667),
        .in(_T_499)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_4802 (
        .y(_T_500),
        .sel(_T_497),
        .a(2'h2),
        .b(_WTEMP_667)
    );
    wire [1:0] _T_501;
    MUX_UNSIGNED #(.width(2)) u_mux_4803 (
        .y(_T_501),
        .sel(_T_495),
        .a(2'h3),
        .b(_T_500)
    );
    wire [1:0] _T_502;
    MUX_UNSIGNED #(.width(2)) u_mux_4804 (
        .y(_T_502),
        .sel(_T_487),
        .a(_T_494),
        .b(_T_501)
    );
    wire [2:0] _T_503;
    CAT #(.width_a(1), .width_b(2)) cat_4805 (
        .y(_T_503),
        .a(_T_487),
        .b(_T_502)
    );
    wire [2:0] _T_504;
    MUX_UNSIGNED #(.width(3)) u_mux_4806 (
        .y(_T_504),
        .sel(_T_463),
        .a(_T_483),
        .b(_T_503)
    );
    wire [3:0] _T_505;
    CAT #(.width_a(1), .width_b(3)) cat_4807 (
        .y(_T_505),
        .a(_T_463),
        .b(_T_504)
    );
    wire [7:0] _T_506;
    BITS #(.width(16), .high(15), .low(8)) bits_4808 (
        .y(_T_506),
        .in(_T_457)
    );
    wire [7:0] _T_507;
    BITS #(.width(16), .high(7), .low(0)) bits_4809 (
        .y(_T_507),
        .in(_T_457)
    );
    wire _T_509;
    wire [7:0] _WTEMP_668;
    PAD_UNSIGNED #(.width(1), .n(8)) u_pad_4810 (
        .y(_WTEMP_668),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(8)) u_neq_4811 (
        .y(_T_509),
        .a(_T_506),
        .b(_WTEMP_668)
    );
    wire [3:0] _T_510;
    BITS #(.width(8), .high(7), .low(4)) bits_4812 (
        .y(_T_510),
        .in(_T_506)
    );
    wire [3:0] _T_511;
    BITS #(.width(8), .high(3), .low(0)) bits_4813 (
        .y(_T_511),
        .in(_T_506)
    );
    wire _T_513;
    wire [3:0] _WTEMP_669;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_4814 (
        .y(_WTEMP_669),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_4815 (
        .y(_T_513),
        .a(_T_510),
        .b(_WTEMP_669)
    );
    wire _T_514;
    BITS #(.width(4), .high(3), .low(3)) bits_4816 (
        .y(_T_514),
        .in(_T_510)
    );
    wire _T_516;
    BITS #(.width(4), .high(2), .low(2)) bits_4817 (
        .y(_T_516),
        .in(_T_510)
    );
    wire _T_518;
    BITS #(.width(4), .high(1), .low(1)) bits_4818 (
        .y(_T_518),
        .in(_T_510)
    );
    wire [1:0] _T_519;
    wire [1:0] _WTEMP_670;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_4819 (
        .y(_WTEMP_670),
        .in(_T_518)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_4820 (
        .y(_T_519),
        .sel(_T_516),
        .a(2'h2),
        .b(_WTEMP_670)
    );
    wire [1:0] _T_520;
    MUX_UNSIGNED #(.width(2)) u_mux_4821 (
        .y(_T_520),
        .sel(_T_514),
        .a(2'h3),
        .b(_T_519)
    );
    wire _T_521;
    BITS #(.width(4), .high(3), .low(3)) bits_4822 (
        .y(_T_521),
        .in(_T_511)
    );
    wire _T_523;
    BITS #(.width(4), .high(2), .low(2)) bits_4823 (
        .y(_T_523),
        .in(_T_511)
    );
    wire _T_525;
    BITS #(.width(4), .high(1), .low(1)) bits_4824 (
        .y(_T_525),
        .in(_T_511)
    );
    wire [1:0] _T_526;
    wire [1:0] _WTEMP_671;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_4825 (
        .y(_WTEMP_671),
        .in(_T_525)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_4826 (
        .y(_T_526),
        .sel(_T_523),
        .a(2'h2),
        .b(_WTEMP_671)
    );
    wire [1:0] _T_527;
    MUX_UNSIGNED #(.width(2)) u_mux_4827 (
        .y(_T_527),
        .sel(_T_521),
        .a(2'h3),
        .b(_T_526)
    );
    wire [1:0] _T_528;
    MUX_UNSIGNED #(.width(2)) u_mux_4828 (
        .y(_T_528),
        .sel(_T_513),
        .a(_T_520),
        .b(_T_527)
    );
    wire [2:0] _T_529;
    CAT #(.width_a(1), .width_b(2)) cat_4829 (
        .y(_T_529),
        .a(_T_513),
        .b(_T_528)
    );
    wire [3:0] _T_530;
    BITS #(.width(8), .high(7), .low(4)) bits_4830 (
        .y(_T_530),
        .in(_T_507)
    );
    wire [3:0] _T_531;
    BITS #(.width(8), .high(3), .low(0)) bits_4831 (
        .y(_T_531),
        .in(_T_507)
    );
    wire _T_533;
    wire [3:0] _WTEMP_672;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_4832 (
        .y(_WTEMP_672),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_4833 (
        .y(_T_533),
        .a(_T_530),
        .b(_WTEMP_672)
    );
    wire _T_534;
    BITS #(.width(4), .high(3), .low(3)) bits_4834 (
        .y(_T_534),
        .in(_T_530)
    );
    wire _T_536;
    BITS #(.width(4), .high(2), .low(2)) bits_4835 (
        .y(_T_536),
        .in(_T_530)
    );
    wire _T_538;
    BITS #(.width(4), .high(1), .low(1)) bits_4836 (
        .y(_T_538),
        .in(_T_530)
    );
    wire [1:0] _T_539;
    wire [1:0] _WTEMP_673;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_4837 (
        .y(_WTEMP_673),
        .in(_T_538)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_4838 (
        .y(_T_539),
        .sel(_T_536),
        .a(2'h2),
        .b(_WTEMP_673)
    );
    wire [1:0] _T_540;
    MUX_UNSIGNED #(.width(2)) u_mux_4839 (
        .y(_T_540),
        .sel(_T_534),
        .a(2'h3),
        .b(_T_539)
    );
    wire _T_541;
    BITS #(.width(4), .high(3), .low(3)) bits_4840 (
        .y(_T_541),
        .in(_T_531)
    );
    wire _T_543;
    BITS #(.width(4), .high(2), .low(2)) bits_4841 (
        .y(_T_543),
        .in(_T_531)
    );
    wire _T_545;
    BITS #(.width(4), .high(1), .low(1)) bits_4842 (
        .y(_T_545),
        .in(_T_531)
    );
    wire [1:0] _T_546;
    wire [1:0] _WTEMP_674;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_4843 (
        .y(_WTEMP_674),
        .in(_T_545)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_4844 (
        .y(_T_546),
        .sel(_T_543),
        .a(2'h2),
        .b(_WTEMP_674)
    );
    wire [1:0] _T_547;
    MUX_UNSIGNED #(.width(2)) u_mux_4845 (
        .y(_T_547),
        .sel(_T_541),
        .a(2'h3),
        .b(_T_546)
    );
    wire [1:0] _T_548;
    MUX_UNSIGNED #(.width(2)) u_mux_4846 (
        .y(_T_548),
        .sel(_T_533),
        .a(_T_540),
        .b(_T_547)
    );
    wire [2:0] _T_549;
    CAT #(.width_a(1), .width_b(2)) cat_4847 (
        .y(_T_549),
        .a(_T_533),
        .b(_T_548)
    );
    wire [2:0] _T_550;
    MUX_UNSIGNED #(.width(3)) u_mux_4848 (
        .y(_T_550),
        .sel(_T_509),
        .a(_T_529),
        .b(_T_549)
    );
    wire [3:0] _T_551;
    CAT #(.width_a(1), .width_b(3)) cat_4849 (
        .y(_T_551),
        .a(_T_509),
        .b(_T_550)
    );
    wire [3:0] _T_552;
    MUX_UNSIGNED #(.width(4)) u_mux_4850 (
        .y(_T_552),
        .sel(_T_459),
        .a(_T_505),
        .b(_T_551)
    );
    wire [4:0] _T_553;
    CAT #(.width_a(1), .width_b(4)) cat_4851 (
        .y(_T_553),
        .a(_T_459),
        .b(_T_552)
    );
    wire [15:0] _T_554;
    BITS #(.width(32), .high(31), .low(16)) bits_4852 (
        .y(_T_554),
        .in(_T_453)
    );
    wire [15:0] _T_555;
    BITS #(.width(32), .high(15), .low(0)) bits_4853 (
        .y(_T_555),
        .in(_T_453)
    );
    wire _T_557;
    wire [15:0] _WTEMP_675;
    PAD_UNSIGNED #(.width(1), .n(16)) u_pad_4854 (
        .y(_WTEMP_675),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(16)) u_neq_4855 (
        .y(_T_557),
        .a(_T_554),
        .b(_WTEMP_675)
    );
    wire [7:0] _T_558;
    BITS #(.width(16), .high(15), .low(8)) bits_4856 (
        .y(_T_558),
        .in(_T_554)
    );
    wire [7:0] _T_559;
    BITS #(.width(16), .high(7), .low(0)) bits_4857 (
        .y(_T_559),
        .in(_T_554)
    );
    wire _T_561;
    wire [7:0] _WTEMP_676;
    PAD_UNSIGNED #(.width(1), .n(8)) u_pad_4858 (
        .y(_WTEMP_676),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(8)) u_neq_4859 (
        .y(_T_561),
        .a(_T_558),
        .b(_WTEMP_676)
    );
    wire [3:0] _T_562;
    BITS #(.width(8), .high(7), .low(4)) bits_4860 (
        .y(_T_562),
        .in(_T_558)
    );
    wire [3:0] _T_563;
    BITS #(.width(8), .high(3), .low(0)) bits_4861 (
        .y(_T_563),
        .in(_T_558)
    );
    wire _T_565;
    wire [3:0] _WTEMP_677;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_4862 (
        .y(_WTEMP_677),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_4863 (
        .y(_T_565),
        .a(_T_562),
        .b(_WTEMP_677)
    );
    wire _T_566;
    BITS #(.width(4), .high(3), .low(3)) bits_4864 (
        .y(_T_566),
        .in(_T_562)
    );
    wire _T_568;
    BITS #(.width(4), .high(2), .low(2)) bits_4865 (
        .y(_T_568),
        .in(_T_562)
    );
    wire _T_570;
    BITS #(.width(4), .high(1), .low(1)) bits_4866 (
        .y(_T_570),
        .in(_T_562)
    );
    wire [1:0] _T_571;
    wire [1:0] _WTEMP_678;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_4867 (
        .y(_WTEMP_678),
        .in(_T_570)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_4868 (
        .y(_T_571),
        .sel(_T_568),
        .a(2'h2),
        .b(_WTEMP_678)
    );
    wire [1:0] _T_572;
    MUX_UNSIGNED #(.width(2)) u_mux_4869 (
        .y(_T_572),
        .sel(_T_566),
        .a(2'h3),
        .b(_T_571)
    );
    wire _T_573;
    BITS #(.width(4), .high(3), .low(3)) bits_4870 (
        .y(_T_573),
        .in(_T_563)
    );
    wire _T_575;
    BITS #(.width(4), .high(2), .low(2)) bits_4871 (
        .y(_T_575),
        .in(_T_563)
    );
    wire _T_577;
    BITS #(.width(4), .high(1), .low(1)) bits_4872 (
        .y(_T_577),
        .in(_T_563)
    );
    wire [1:0] _T_578;
    wire [1:0] _WTEMP_679;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_4873 (
        .y(_WTEMP_679),
        .in(_T_577)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_4874 (
        .y(_T_578),
        .sel(_T_575),
        .a(2'h2),
        .b(_WTEMP_679)
    );
    wire [1:0] _T_579;
    MUX_UNSIGNED #(.width(2)) u_mux_4875 (
        .y(_T_579),
        .sel(_T_573),
        .a(2'h3),
        .b(_T_578)
    );
    wire [1:0] _T_580;
    MUX_UNSIGNED #(.width(2)) u_mux_4876 (
        .y(_T_580),
        .sel(_T_565),
        .a(_T_572),
        .b(_T_579)
    );
    wire [2:0] _T_581;
    CAT #(.width_a(1), .width_b(2)) cat_4877 (
        .y(_T_581),
        .a(_T_565),
        .b(_T_580)
    );
    wire [3:0] _T_582;
    BITS #(.width(8), .high(7), .low(4)) bits_4878 (
        .y(_T_582),
        .in(_T_559)
    );
    wire [3:0] _T_583;
    BITS #(.width(8), .high(3), .low(0)) bits_4879 (
        .y(_T_583),
        .in(_T_559)
    );
    wire _T_585;
    wire [3:0] _WTEMP_680;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_4880 (
        .y(_WTEMP_680),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_4881 (
        .y(_T_585),
        .a(_T_582),
        .b(_WTEMP_680)
    );
    wire _T_586;
    BITS #(.width(4), .high(3), .low(3)) bits_4882 (
        .y(_T_586),
        .in(_T_582)
    );
    wire _T_588;
    BITS #(.width(4), .high(2), .low(2)) bits_4883 (
        .y(_T_588),
        .in(_T_582)
    );
    wire _T_590;
    BITS #(.width(4), .high(1), .low(1)) bits_4884 (
        .y(_T_590),
        .in(_T_582)
    );
    wire [1:0] _T_591;
    wire [1:0] _WTEMP_681;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_4885 (
        .y(_WTEMP_681),
        .in(_T_590)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_4886 (
        .y(_T_591),
        .sel(_T_588),
        .a(2'h2),
        .b(_WTEMP_681)
    );
    wire [1:0] _T_592;
    MUX_UNSIGNED #(.width(2)) u_mux_4887 (
        .y(_T_592),
        .sel(_T_586),
        .a(2'h3),
        .b(_T_591)
    );
    wire _T_593;
    BITS #(.width(4), .high(3), .low(3)) bits_4888 (
        .y(_T_593),
        .in(_T_583)
    );
    wire _T_595;
    BITS #(.width(4), .high(2), .low(2)) bits_4889 (
        .y(_T_595),
        .in(_T_583)
    );
    wire _T_597;
    BITS #(.width(4), .high(1), .low(1)) bits_4890 (
        .y(_T_597),
        .in(_T_583)
    );
    wire [1:0] _T_598;
    wire [1:0] _WTEMP_682;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_4891 (
        .y(_WTEMP_682),
        .in(_T_597)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_4892 (
        .y(_T_598),
        .sel(_T_595),
        .a(2'h2),
        .b(_WTEMP_682)
    );
    wire [1:0] _T_599;
    MUX_UNSIGNED #(.width(2)) u_mux_4893 (
        .y(_T_599),
        .sel(_T_593),
        .a(2'h3),
        .b(_T_598)
    );
    wire [1:0] _T_600;
    MUX_UNSIGNED #(.width(2)) u_mux_4894 (
        .y(_T_600),
        .sel(_T_585),
        .a(_T_592),
        .b(_T_599)
    );
    wire [2:0] _T_601;
    CAT #(.width_a(1), .width_b(2)) cat_4895 (
        .y(_T_601),
        .a(_T_585),
        .b(_T_600)
    );
    wire [2:0] _T_602;
    MUX_UNSIGNED #(.width(3)) u_mux_4896 (
        .y(_T_602),
        .sel(_T_561),
        .a(_T_581),
        .b(_T_601)
    );
    wire [3:0] _T_603;
    CAT #(.width_a(1), .width_b(3)) cat_4897 (
        .y(_T_603),
        .a(_T_561),
        .b(_T_602)
    );
    wire [7:0] _T_604;
    BITS #(.width(16), .high(15), .low(8)) bits_4898 (
        .y(_T_604),
        .in(_T_555)
    );
    wire [7:0] _T_605;
    BITS #(.width(16), .high(7), .low(0)) bits_4899 (
        .y(_T_605),
        .in(_T_555)
    );
    wire _T_607;
    wire [7:0] _WTEMP_683;
    PAD_UNSIGNED #(.width(1), .n(8)) u_pad_4900 (
        .y(_WTEMP_683),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(8)) u_neq_4901 (
        .y(_T_607),
        .a(_T_604),
        .b(_WTEMP_683)
    );
    wire [3:0] _T_608;
    BITS #(.width(8), .high(7), .low(4)) bits_4902 (
        .y(_T_608),
        .in(_T_604)
    );
    wire [3:0] _T_609;
    BITS #(.width(8), .high(3), .low(0)) bits_4903 (
        .y(_T_609),
        .in(_T_604)
    );
    wire _T_611;
    wire [3:0] _WTEMP_684;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_4904 (
        .y(_WTEMP_684),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_4905 (
        .y(_T_611),
        .a(_T_608),
        .b(_WTEMP_684)
    );
    wire _T_612;
    BITS #(.width(4), .high(3), .low(3)) bits_4906 (
        .y(_T_612),
        .in(_T_608)
    );
    wire _T_614;
    BITS #(.width(4), .high(2), .low(2)) bits_4907 (
        .y(_T_614),
        .in(_T_608)
    );
    wire _T_616;
    BITS #(.width(4), .high(1), .low(1)) bits_4908 (
        .y(_T_616),
        .in(_T_608)
    );
    wire [1:0] _T_617;
    wire [1:0] _WTEMP_685;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_4909 (
        .y(_WTEMP_685),
        .in(_T_616)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_4910 (
        .y(_T_617),
        .sel(_T_614),
        .a(2'h2),
        .b(_WTEMP_685)
    );
    wire [1:0] _T_618;
    MUX_UNSIGNED #(.width(2)) u_mux_4911 (
        .y(_T_618),
        .sel(_T_612),
        .a(2'h3),
        .b(_T_617)
    );
    wire _T_619;
    BITS #(.width(4), .high(3), .low(3)) bits_4912 (
        .y(_T_619),
        .in(_T_609)
    );
    wire _T_621;
    BITS #(.width(4), .high(2), .low(2)) bits_4913 (
        .y(_T_621),
        .in(_T_609)
    );
    wire _T_623;
    BITS #(.width(4), .high(1), .low(1)) bits_4914 (
        .y(_T_623),
        .in(_T_609)
    );
    wire [1:0] _T_624;
    wire [1:0] _WTEMP_686;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_4915 (
        .y(_WTEMP_686),
        .in(_T_623)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_4916 (
        .y(_T_624),
        .sel(_T_621),
        .a(2'h2),
        .b(_WTEMP_686)
    );
    wire [1:0] _T_625;
    MUX_UNSIGNED #(.width(2)) u_mux_4917 (
        .y(_T_625),
        .sel(_T_619),
        .a(2'h3),
        .b(_T_624)
    );
    wire [1:0] _T_626;
    MUX_UNSIGNED #(.width(2)) u_mux_4918 (
        .y(_T_626),
        .sel(_T_611),
        .a(_T_618),
        .b(_T_625)
    );
    wire [2:0] _T_627;
    CAT #(.width_a(1), .width_b(2)) cat_4919 (
        .y(_T_627),
        .a(_T_611),
        .b(_T_626)
    );
    wire [3:0] _T_628;
    BITS #(.width(8), .high(7), .low(4)) bits_4920 (
        .y(_T_628),
        .in(_T_605)
    );
    wire [3:0] _T_629;
    BITS #(.width(8), .high(3), .low(0)) bits_4921 (
        .y(_T_629),
        .in(_T_605)
    );
    wire _T_631;
    wire [3:0] _WTEMP_687;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_4922 (
        .y(_WTEMP_687),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_4923 (
        .y(_T_631),
        .a(_T_628),
        .b(_WTEMP_687)
    );
    wire _T_632;
    BITS #(.width(4), .high(3), .low(3)) bits_4924 (
        .y(_T_632),
        .in(_T_628)
    );
    wire _T_634;
    BITS #(.width(4), .high(2), .low(2)) bits_4925 (
        .y(_T_634),
        .in(_T_628)
    );
    wire _T_636;
    BITS #(.width(4), .high(1), .low(1)) bits_4926 (
        .y(_T_636),
        .in(_T_628)
    );
    wire [1:0] _T_637;
    wire [1:0] _WTEMP_688;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_4927 (
        .y(_WTEMP_688),
        .in(_T_636)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_4928 (
        .y(_T_637),
        .sel(_T_634),
        .a(2'h2),
        .b(_WTEMP_688)
    );
    wire [1:0] _T_638;
    MUX_UNSIGNED #(.width(2)) u_mux_4929 (
        .y(_T_638),
        .sel(_T_632),
        .a(2'h3),
        .b(_T_637)
    );
    wire _T_639;
    BITS #(.width(4), .high(3), .low(3)) bits_4930 (
        .y(_T_639),
        .in(_T_629)
    );
    wire _T_641;
    BITS #(.width(4), .high(2), .low(2)) bits_4931 (
        .y(_T_641),
        .in(_T_629)
    );
    wire _T_643;
    BITS #(.width(4), .high(1), .low(1)) bits_4932 (
        .y(_T_643),
        .in(_T_629)
    );
    wire [1:0] _T_644;
    wire [1:0] _WTEMP_689;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_4933 (
        .y(_WTEMP_689),
        .in(_T_643)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_4934 (
        .y(_T_644),
        .sel(_T_641),
        .a(2'h2),
        .b(_WTEMP_689)
    );
    wire [1:0] _T_645;
    MUX_UNSIGNED #(.width(2)) u_mux_4935 (
        .y(_T_645),
        .sel(_T_639),
        .a(2'h3),
        .b(_T_644)
    );
    wire [1:0] _T_646;
    MUX_UNSIGNED #(.width(2)) u_mux_4936 (
        .y(_T_646),
        .sel(_T_631),
        .a(_T_638),
        .b(_T_645)
    );
    wire [2:0] _T_647;
    CAT #(.width_a(1), .width_b(2)) cat_4937 (
        .y(_T_647),
        .a(_T_631),
        .b(_T_646)
    );
    wire [2:0] _T_648;
    MUX_UNSIGNED #(.width(3)) u_mux_4938 (
        .y(_T_648),
        .sel(_T_607),
        .a(_T_627),
        .b(_T_647)
    );
    wire [3:0] _T_649;
    CAT #(.width_a(1), .width_b(3)) cat_4939 (
        .y(_T_649),
        .a(_T_607),
        .b(_T_648)
    );
    wire [3:0] _T_650;
    MUX_UNSIGNED #(.width(4)) u_mux_4940 (
        .y(_T_650),
        .sel(_T_557),
        .a(_T_603),
        .b(_T_649)
    );
    wire [4:0] _T_651;
    CAT #(.width_a(1), .width_b(4)) cat_4941 (
        .y(_T_651),
        .a(_T_557),
        .b(_T_650)
    );
    wire [4:0] _T_652;
    MUX_UNSIGNED #(.width(5)) u_mux_4942 (
        .y(_T_652),
        .sel(_T_455),
        .a(_T_553),
        .b(_T_651)
    );
    wire [5:0] _T_653;
    CAT #(.width_a(1), .width_b(5)) cat_4943 (
        .y(_T_653),
        .a(_T_455),
        .b(_T_652)
    );
    wire [6:0] _T_655;
    ADD_UNSIGNED #(.width(6)) u_add_4944 (
        .y(_T_655),
        .a(6'h3F),
        .b(_T_450)
    );
    wire [5:0] _T_656;
    TAIL #(.width(7), .n(1)) tail_4945 (
        .y(_T_656),
        .in(_T_655)
    );
    wire [6:0] _T_657;
    SUB_UNSIGNED #(.width(6)) u_sub_4946 (
        .y(_T_657),
        .a(_T_656),
        .b(_T_653)
    );
    wire [6:0] _T_658;
    ASUINT #(.width(7)) asuint_4947 (
        .y(_T_658),
        .in(_T_657)
    );
    wire [5:0] _T_659;
    TAIL #(.width(7), .n(1)) tail_4948 (
        .y(_T_659),
        .in(_T_658)
    );
    wire _T_660;
    GT_UNSIGNED #(.width(6)) u_gt_4949 (
        .y(_T_660),
        .a(_T_450),
        .b(_T_653)
    );
    wire _T_662;
    wire [6:0] _WTEMP_690;
    PAD_UNSIGNED #(.width(1), .n(7)) u_pad_4950 (
        .y(_WTEMP_690),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(7)) u_eq_4951 (
        .y(_T_662),
        .a(_count__q),
        .b(_WTEMP_690)
    );
    wire _T_664;
    EQ_UNSIGNED #(.width(1)) u_eq_4952 (
        .y(_T_664),
        .a(_T_247),
        .b(1'h0)
    );
    wire _T_665;
    BITWISEAND #(.width(1)) bitwiseand_4953 (
        .y(_T_665),
        .a(_T_662),
        .b(_T_664)
    );
    wire _T_667;
    wire [5:0] _WTEMP_691;
    PAD_UNSIGNED #(.width(1), .n(6)) u_pad_4954 (
        .y(_WTEMP_691),
        .in(1'h1)
    );
    GEQ_UNSIGNED #(.width(6)) u_geq_4955 (
        .y(_T_667),
        .a(_T_659),
        .b(_WTEMP_691)
    );
    wire _T_668;
    BITWISEOR #(.width(1)) bitwiseor_4956 (
        .y(_T_668),
        .a(_T_667),
        .b(_T_660)
    );
    wire _T_669;
    BITWISEAND #(.width(1)) bitwiseand_4957 (
        .y(_T_669),
        .a(_T_665),
        .b(_T_668)
    );
    wire [5:0] _T_671;
    MUX_UNSIGNED #(.width(6)) u_mux_4958 (
        .y(_T_671),
        .sel(_T_660),
        .a(6'h3F),
        .b(_T_659)
    );
    wire [5:0] _T_672;
    SHR_UNSIGNED #(.width(6), .n(0)) u_shr_4959 (
        .y(_T_672),
        .in(_T_671)
    );
    wire [5:0] _T_673;
    SHL_UNSIGNED #(.width(6), .n(0)) u_shl_4960 (
        .y(_T_673),
        .in(_T_672)
    );
    wire [63:0] _T_674;
    BITS #(.width(130), .high(63), .low(0)) bits_4961 (
        .y(_T_674),
        .in(_remainder__q)
    );
    wire [126:0] _T_675;
    DSHL_UNSIGNED #(.width_in(64), .width_n(6)) u_dshl_4962 (
        .y(_T_675),
        .in(_T_674),
        .n(_T_673)
    );
    wire _T_677;
    EQ_UNSIGNED #(.width(1)) u_eq_4963 (
        .y(_T_677),
        .a(_isHi__q),
        .b(1'h0)
    );
    wire _T_678;
    BITWISEAND #(.width(1)) bitwiseand_4964 (
        .y(_T_678),
        .a(_T_247),
        .b(_T_677)
    );
    wire [6:0] _node_351;
    wire [6:0] _WTEMP_692;
    PAD_UNSIGNED #(.width(6), .n(7)) u_pad_4965 (
        .y(_WTEMP_692),
        .in(_T_672)
    );
    MUX_UNSIGNED #(.width(7)) u_mux_4966 (
        .y(_node_351),
        .sel(_T_669),
        .a(_WTEMP_692),
        .b(_T_241)
    );
    wire [6:0] _node_352;
    MUX_UNSIGNED #(.width(7)) u_mux_4967 (
        .y(_node_352),
        .sel(_T_161),
        .a(_T_217),
        .b(_count__q)
    );
    wire _node_353;
    MUX_UNSIGNED #(.width(1)) u_mux_4968 (
        .y(_node_353),
        .sel(_T_678),
        .a(1'h0),
        .b(_neg_out__q)
    );
    wire [128:0] _node_354;
    wire [128:0] _WTEMP_693;
    PAD_UNSIGNED #(.width(127), .n(129)) u_pad_4969 (
        .y(_WTEMP_693),
        .in(_T_675)
    );
    MUX_UNSIGNED #(.width(129)) u_mux_4970 (
        .y(_node_354),
        .sel(_T_669),
        .a(_WTEMP_693),
        .b(_T_234)
    );
    wire [129:0] _node_355;
    MUX_UNSIGNED #(.width(130)) u_mux_4971 (
        .y(_node_355),
        .sel(_T_161),
        .a(_T_214),
        .b(_node_347)
    );
    wire [2:0] _node_356;
    MUX_UNSIGNED #(.width(3)) u_mux_4972 (
        .y(_node_356),
        .sel(_T_236),
        .a(_T_238),
        .b(_node_350)
    );
    wire [2:0] _node_357;
    MUX_UNSIGNED #(.width(3)) u_mux_4973 (
        .y(_node_357),
        .sel(_T_161),
        .a(_node_348),
        .b(_node_349)
    );
    wire _T_680;
    BITWISEAND #(.width(1)) bitwiseand_4974 (
        .y(_T_680),
        .a(io_resp_ready),
        .b(io_resp_valid)
    );
    wire _T_681;
    BITWISEOR #(.width(1)) bitwiseor_4975 (
        .y(_T_681),
        .a(_T_680),
        .b(io_kill)
    );
    wire [2:0] _node_358;
    MUX_UNSIGNED #(.width(3)) u_mux_4976 (
        .y(_node_358),
        .sel(_T_225),
        .a(_node_356),
        .b(_node_357)
    );
    wire _T_682;
    BITWISEAND #(.width(1)) bitwiseand_4977 (
        .y(_T_682),
        .a(io_req_ready),
        .b(io_req_valid)
    );
    wire _T_684;
    EQ_UNSIGNED #(.width(1)) u_eq_4978 (
        .y(_T_684),
        .a(cmdMul),
        .b(1'h0)
    );
    wire _T_685;
    BITWISEAND #(.width(1)) bitwiseand_4979 (
        .y(_T_685),
        .a(rhs_sign),
        .b(_T_684)
    );
    wire _T_686;
    BITWISEOR #(.width(1)) bitwiseor_4980 (
        .y(_T_686),
        .a(lhs_sign),
        .b(_T_685)
    );
    wire [2:0] _T_687;
    MUX_UNSIGNED #(.width(3)) u_mux_4981 (
        .y(_T_687),
        .sel(_T_686),
        .a(3'h1),
        .b(3'h2)
    );
    wire _T_690;
    EQ_UNSIGNED #(.width(1)) u_eq_4982 (
        .y(_T_690),
        .a(cmdMul),
        .b(1'h0)
    );
    wire _T_691;
    NEQ_UNSIGNED #(.width(1)) u_neq_4983 (
        .y(_T_691),
        .a(lhs_sign),
        .b(rhs_sign)
    );
    wire _T_692;
    MUX_UNSIGNED #(.width(1)) u_mux_4984 (
        .y(_T_692),
        .sel(cmdHi),
        .a(lhs_sign),
        .b(_T_691)
    );
    wire _T_693;
    BITWISEAND #(.width(1)) bitwiseand_4985 (
        .y(_T_693),
        .a(_T_690),
        .b(_T_692)
    );
    wire [64:0] _T_694;
    CAT #(.width_a(1), .width_b(64)) cat_4986 (
        .y(_T_694),
        .a(rhs_sign),
        .b(rhs_in)
    );
    wire [6:0] _node_359;
    MUX_UNSIGNED #(.width(7)) u_mux_4987 (
        .y(_node_359),
        .sel(_T_225),
        .a(_node_351),
        .b(_node_352)
    );
    wire [64:0] _node_360;
    MUX_UNSIGNED #(.width(65)) u_mux_4988 (
        .y(_node_360),
        .sel(_T_151),
        .a(_node_340),
        .b(_divisor__q)
    );
    wire _node_361;
    MUX_UNSIGNED #(.width(1)) u_mux_4989 (
        .y(_node_361),
        .sel(_T_225),
        .a(_node_353),
        .b(_neg_out__q)
    );
    wire [129:0] _node_362;
    wire [129:0] _WTEMP_694;
    PAD_UNSIGNED #(.width(129), .n(130)) u_pad_4990 (
        .y(_WTEMP_694),
        .in(_node_354)
    );
    MUX_UNSIGNED #(.width(130)) u_mux_4991 (
        .y(_node_362),
        .sel(_T_225),
        .a(_WTEMP_694),
        .b(_node_355)
    );
    wire [2:0] _node_363;
    MUX_UNSIGNED #(.width(3)) u_mux_4992 (
        .y(_node_363),
        .sel(_T_681),
        .a(3'h0),
        .b(_node_358)
    );
    wire _T_697;
    EQ_UNSIGNED #(.width(1)) u_eq_4993 (
        .y(_T_697),
        .a(_req_dw__q),
        .b(1'h0)
    );
    wire _T_698;
    BITWISEAND #(.width(1)) bitwiseand_4994 (
        .y(_T_698),
        .a(1'h1),
        .b(_T_697)
    );
    wire _T_699;
    BITS #(.width(130), .high(31), .low(31)) bits_4995 (
        .y(_T_699),
        .in(_remainder__q)
    );
    wire _T_700;
    BITS #(.width(1), .high(0), .low(0)) bits_4996 (
        .y(_T_700),
        .in(_T_699)
    );
    wire [31:0] _T_703;
    MUX_UNSIGNED #(.width(32)) u_mux_4997 (
        .y(_T_703),
        .sel(_T_700),
        .a(32'hFFFFFFFF),
        .b(32'h0)
    );
    wire [31:0] _T_704;
    BITS #(.width(130), .high(31), .low(0)) bits_4998 (
        .y(_T_704),
        .in(_remainder__q)
    );
    wire [63:0] _T_705;
    CAT #(.width_a(32), .width_b(32)) cat_4999 (
        .y(_T_705),
        .a(_T_703),
        .b(_T_704)
    );
    wire [63:0] _T_706;
    BITS #(.width(130), .high(63), .low(0)) bits_5000 (
        .y(_T_706),
        .in(_remainder__q)
    );
    wire [63:0] _T_707;
    MUX_UNSIGNED #(.width(64)) u_mux_5001 (
        .y(_T_707),
        .sel(_T_698),
        .a(_T_705),
        .b(_T_706)
    );
    wire _T_708;
    EQ_UNSIGNED #(.width(3)) u_eq_5002 (
        .y(_T_708),
        .a(_state__q),
        .b(3'h5)
    );
    wire _T_709;
    EQ_UNSIGNED #(.width(3)) u_eq_5003 (
        .y(_T_709),
        .a(_state__q),
        .b(3'h0)
    );
    wire [6:0] _WTEMP_695;
    PAD_UNSIGNED #(.width(1), .n(7)) u_pad_5004 (
        .y(_WTEMP_695),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(7)) u_mux_5005 (
        .y(_count__d),
        .sel(_T_682),
        .a(_WTEMP_695),
        .b(_node_359)
    );
    MUX_UNSIGNED #(.width(65)) u_mux_5006 (
        .y(_divisor__d),
        .sel(_T_682),
        .a(_T_694),
        .b(_node_360)
    );
    assign io_req_ready = _T_709;
    assign io_resp_bits_data = _T_707;
    assign io_resp_bits_tag = _req_tag__q;
    assign io_resp_valid = _T_708;
    MUX_UNSIGNED #(.width(1)) u_mux_5007 (
        .y(_isHi__d),
        .sel(_T_682),
        .a(cmdHi),
        .b(_isHi__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_5008 (
        .y(_isMul__d),
        .sel(_T_682),
        .a(cmdMul),
        .b(_isMul__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_5009 (
        .y(_neg_out__d),
        .sel(_T_682),
        .a(_T_693),
        .b(_node_361)
    );
    wire [129:0] _WTEMP_696;
    PAD_UNSIGNED #(.width(64), .n(130)) u_pad_5010 (
        .y(_WTEMP_696),
        .in(lhs_in)
    );
    MUX_UNSIGNED #(.width(130)) u_mux_5011 (
        .y(_remainder__d),
        .sel(_T_682),
        .a(_WTEMP_696),
        .b(_node_362)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_5012 (
        .y(_req_dw__d),
        .sel(_T_682),
        .a(io_req_bits_dw),
        .b(_req_dw__q)
    );
    MUX_UNSIGNED #(.width(4)) u_mux_5013 (
        .y(_req_fn__d),
        .sel(_T_682),
        .a(io_req_bits_fn),
        .b(_req_fn__q)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_5014 (
        .y(_req_in1__d),
        .sel(_T_682),
        .a(io_req_bits_in1),
        .b(_req_in1__q)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_5015 (
        .y(_req_in2__d),
        .sel(_T_682),
        .a(io_req_bits_in2),
        .b(_req_in2__q)
    );
    MUX_UNSIGNED #(.width(5)) u_mux_5016 (
        .y(_req_tag__d),
        .sel(_T_682),
        .a(io_req_bits_tag),
        .b(_req_tag__q)
    );
    MUX_UNSIGNED #(.width(3)) u_mux_5017 (
        .y(_WTEMP_614),
        .sel(_T_682),
        .a(_T_687),
        .b(_node_363)
    );
endmodule //MulDiv
module MUL2_SIGNED(y, a, b);
    parameter width_a = 4;
    parameter width_b = 4;
    output [width_a+width_b-1:0] y;
    input [width_a-1:0] a;
    input [width_b-1:0] b;
    assign y = $signed(a) * $signed(b);
endmodule // MUL2_SIGNED
module MUL2_UNSIGNED(y, a, b);
    parameter width_a = 4;
    parameter width_b = 4;
    output [width_a+width_b-1:0] y;
    input [width_a-1:0] a;
    input [width_b-1:0] b;
    assign y = a * b;
endmodule // MUL2_UNSIGNED
module NEQ_SIGNED(y, a, b);
    parameter width = 4;
    output y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = $signed(a) != $signed(b);
endmodule // NEQ_SIGNED
module EQ_SIGNED(y, a, b);
    parameter width = 4;
    output y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = $signed(a) == $signed(b);
endmodule // EQ_SIGNED
