module FPU(
    input clock,
    input reset,
    input [31:0] io_inst,
    input [63:0] io_fromint_data,
    input [2:0] io_fcsr_rm,
    output io_fcsr_flags_valid,
    output [4:0] io_fcsr_flags_bits,
    output [63:0] io_store_data,
    output [63:0] io_toint_data,
    input io_dmem_resp_val,
    input [2:0] io_dmem_resp_type,
    input [4:0] io_dmem_resp_tag,
    input [63:0] io_dmem_resp_data,
    input io_valid,
    output io_fcsr_rdy,
    output io_nack_mem,
    output io_illegal_rm,
    input io_killx,
    input io_killm,
    output [4:0] io_dec_cmd,
    output io_dec_ldst,
    output io_dec_wen,
    output io_dec_ren1,
    output io_dec_ren2,
    output io_dec_ren3,
    output io_dec_swap12,
    output io_dec_swap23,
    output io_dec_single,
    output io_dec_fromint,
    output io_dec_toint,
    output io_dec_fastpipe,
    output io_dec_fma,
    output io_dec_div,
    output io_dec_sqrt,
    output io_dec_wflags,
    output io_sboard_set,
    output io_sboard_clr,
    output [4:0] io_sboard_clra,
    output io_cp_req_ready,
    input io_cp_req_valid,
    input [4:0] io_cp_req_bits_cmd,
    input io_cp_req_bits_ldst,
    input io_cp_req_bits_wen,
    input io_cp_req_bits_ren1,
    input io_cp_req_bits_ren2,
    input io_cp_req_bits_ren3,
    input io_cp_req_bits_swap12,
    input io_cp_req_bits_swap23,
    input io_cp_req_bits_single,
    input io_cp_req_bits_fromint,
    input io_cp_req_bits_toint,
    input io_cp_req_bits_fastpipe,
    input io_cp_req_bits_fma,
    input io_cp_req_bits_div,
    input io_cp_req_bits_sqrt,
    input io_cp_req_bits_wflags,
    input [2:0] io_cp_req_bits_rm,
    input [1:0] io_cp_req_bits_typ,
    input [64:0] io_cp_req_bits_in1,
    input [64:0] io_cp_req_bits_in2,
    input [64:0] io_cp_req_bits_in3,
    input io_cp_resp_ready,
    output io_cp_resp_valid,
    output [64:0] io_cp_resp_bits_data,
    output [4:0] io_cp_resp_bits_exc
);
    wire _ex_reg_valid__q;
    wire _ex_reg_valid__d;
    DFF_POSCLK #(.width(1)) ex_reg_valid (
        .q(_ex_reg_valid__q),
        .d(_ex_reg_valid__d),
        .clk(clock)
    );
    wire _WTEMP_0;
    MUX_UNSIGNED #(.width(1)) u_mux_1 (
        .y(_ex_reg_valid__d),
        .sel(reset),
        .a(1'h0),
        .b(_WTEMP_0)
    );
    wire req_valid;
    BITWISEOR #(.width(1)) bitwiseor_2 (
        .y(req_valid),
        .a(_ex_reg_valid__q),
        .b(io_cp_req_valid)
    );
    wire [31:0] _ex_reg_inst__q;
    wire [31:0] _ex_reg_inst__d;
    DFF_POSCLK #(.width(32)) ex_reg_inst (
        .q(_ex_reg_inst__q),
        .d(_ex_reg_inst__d),
        .clk(clock)
    );
    wire ex_cp_valid;
    BITWISEAND #(.width(1)) bitwiseand_3 (
        .y(ex_cp_valid),
        .a(io_cp_req_ready),
        .b(io_cp_req_valid)
    );
    wire _T_215;
    EQ_UNSIGNED #(.width(1)) u_eq_4 (
        .y(_T_215),
        .a(io_killx),
        .b(1'h0)
    );
    wire _T_216;
    BITWISEAND #(.width(1)) bitwiseand_5 (
        .y(_T_216),
        .a(_ex_reg_valid__q),
        .b(_T_215)
    );
    wire _T_217;
    BITWISEOR #(.width(1)) bitwiseor_6 (
        .y(_T_217),
        .a(_T_216),
        .b(ex_cp_valid)
    );
    wire _mem_reg_valid__q;
    wire _mem_reg_valid__d;
    DFF_POSCLK #(.width(1)) mem_reg_valid (
        .q(_mem_reg_valid__q),
        .d(_mem_reg_valid__d),
        .clk(clock)
    );
    wire _WTEMP_1;
    MUX_UNSIGNED #(.width(1)) u_mux_7 (
        .y(_mem_reg_valid__d),
        .sel(reset),
        .a(1'h0),
        .b(_WTEMP_1)
    );
    wire [31:0] _mem_reg_inst__q;
    wire [31:0] _mem_reg_inst__d;
    DFF_POSCLK #(.width(32)) mem_reg_inst (
        .q(_mem_reg_inst__q),
        .d(_mem_reg_inst__d),
        .clk(clock)
    );
    wire _mem_cp_valid__q;
    wire _mem_cp_valid__d;
    DFF_POSCLK #(.width(1)) mem_cp_valid (
        .q(_mem_cp_valid__q),
        .d(_mem_cp_valid__d),
        .clk(clock)
    );
    wire _WTEMP_2;
    MUX_UNSIGNED #(.width(1)) u_mux_8 (
        .y(_mem_cp_valid__d),
        .sel(reset),
        .a(1'h0),
        .b(_WTEMP_2)
    );
    wire _T_221;
    BITWISEOR #(.width(1)) bitwiseor_9 (
        .y(_T_221),
        .a(io_killm),
        .b(io_nack_mem)
    );
    wire _T_223;
    EQ_UNSIGNED #(.width(1)) u_eq_10 (
        .y(_T_223),
        .a(_mem_cp_valid__q),
        .b(1'h0)
    );
    wire killm;
    BITWISEAND #(.width(1)) bitwiseand_11 (
        .y(killm),
        .a(_T_221),
        .b(_T_223)
    );
    wire _T_225;
    EQ_UNSIGNED #(.width(1)) u_eq_12 (
        .y(_T_225),
        .a(killm),
        .b(1'h0)
    );
    wire _T_226;
    BITWISEOR #(.width(1)) bitwiseor_13 (
        .y(_T_226),
        .a(_T_225),
        .b(_mem_cp_valid__q)
    );
    wire _T_227;
    BITWISEAND #(.width(1)) bitwiseand_14 (
        .y(_T_227),
        .a(_mem_reg_valid__q),
        .b(_T_226)
    );
    wire _wb_reg_valid__q;
    wire _wb_reg_valid__d;
    DFF_POSCLK #(.width(1)) wb_reg_valid (
        .q(_wb_reg_valid__q),
        .d(_wb_reg_valid__d),
        .clk(clock)
    );
    wire _WTEMP_3;
    MUX_UNSIGNED #(.width(1)) u_mux_15 (
        .y(_wb_reg_valid__d),
        .sel(reset),
        .a(1'h0),
        .b(_WTEMP_3)
    );
    wire _wb_cp_valid__q;
    wire _wb_cp_valid__d;
    DFF_POSCLK #(.width(1)) wb_cp_valid (
        .q(_wb_cp_valid__q),
        .d(_wb_cp_valid__d),
        .clk(clock)
    );
    wire _WTEMP_4;
    MUX_UNSIGNED #(.width(1)) u_mux_16 (
        .y(_wb_cp_valid__d),
        .sel(reset),
        .a(1'h0),
        .b(_WTEMP_4)
    );
    wire _fp_decoder__clock;
    wire _fp_decoder__reset;
    wire [31:0] _fp_decoder__io_inst;
    wire [4:0] _fp_decoder__io_sigs_cmd;
    wire _fp_decoder__io_sigs_ldst;
    wire _fp_decoder__io_sigs_wen;
    wire _fp_decoder__io_sigs_ren1;
    wire _fp_decoder__io_sigs_ren2;
    wire _fp_decoder__io_sigs_ren3;
    wire _fp_decoder__io_sigs_swap12;
    wire _fp_decoder__io_sigs_swap23;
    wire _fp_decoder__io_sigs_single;
    wire _fp_decoder__io_sigs_fromint;
    wire _fp_decoder__io_sigs_toint;
    wire _fp_decoder__io_sigs_fastpipe;
    wire _fp_decoder__io_sigs_fma;
    wire _fp_decoder__io_sigs_div;
    wire _fp_decoder__io_sigs_sqrt;
    wire _fp_decoder__io_sigs_wflags;
    FPUDecoder fp_decoder (
        .clock(_fp_decoder__clock),
        .reset(_fp_decoder__reset),
        .io_inst(_fp_decoder__io_inst),
        .io_sigs_cmd(_fp_decoder__io_sigs_cmd),
        .io_sigs_ldst(_fp_decoder__io_sigs_ldst),
        .io_sigs_wen(_fp_decoder__io_sigs_wen),
        .io_sigs_ren1(_fp_decoder__io_sigs_ren1),
        .io_sigs_ren2(_fp_decoder__io_sigs_ren2),
        .io_sigs_ren3(_fp_decoder__io_sigs_ren3),
        .io_sigs_swap12(_fp_decoder__io_sigs_swap12),
        .io_sigs_swap23(_fp_decoder__io_sigs_swap23),
        .io_sigs_single(_fp_decoder__io_sigs_single),
        .io_sigs_fromint(_fp_decoder__io_sigs_fromint),
        .io_sigs_toint(_fp_decoder__io_sigs_toint),
        .io_sigs_fastpipe(_fp_decoder__io_sigs_fastpipe),
        .io_sigs_fma(_fp_decoder__io_sigs_fma),
        .io_sigs_div(_fp_decoder__io_sigs_div),
        .io_sigs_sqrt(_fp_decoder__io_sigs_sqrt),
        .io_sigs_wflags(_fp_decoder__io_sigs_wflags)
    );
    wire [4:0] cp_ctrl_cmd;
    wire cp_ctrl_ldst;
    wire cp_ctrl_wen;
    wire cp_ctrl_ren1;
    wire cp_ctrl_ren2;
    wire cp_ctrl_ren3;
    wire cp_ctrl_swap12;
    wire cp_ctrl_swap23;
    wire cp_ctrl_single;
    wire cp_ctrl_fromint;
    wire cp_ctrl_toint;
    wire cp_ctrl_fastpipe;
    wire cp_ctrl_fma;
    wire cp_ctrl_div;
    wire cp_ctrl_sqrt;
    wire cp_ctrl_wflags;
    wire [4:0] __T_282_cmd__q;
    wire [4:0] __T_282_cmd__d;
    DFF_POSCLK #(.width(5)) _T_282_cmd (
        .q(__T_282_cmd__q),
        .d(__T_282_cmd__d),
        .clk(clock)
    );
    wire __T_282_ldst__q;
    wire __T_282_ldst__d;
    DFF_POSCLK #(.width(1)) _T_282_ldst (
        .q(__T_282_ldst__q),
        .d(__T_282_ldst__d),
        .clk(clock)
    );
    wire __T_282_wen__q;
    wire __T_282_wen__d;
    DFF_POSCLK #(.width(1)) _T_282_wen (
        .q(__T_282_wen__q),
        .d(__T_282_wen__d),
        .clk(clock)
    );
    wire __T_282_ren1__q;
    wire __T_282_ren1__d;
    DFF_POSCLK #(.width(1)) _T_282_ren1 (
        .q(__T_282_ren1__q),
        .d(__T_282_ren1__d),
        .clk(clock)
    );
    wire __T_282_ren2__q;
    wire __T_282_ren2__d;
    DFF_POSCLK #(.width(1)) _T_282_ren2 (
        .q(__T_282_ren2__q),
        .d(__T_282_ren2__d),
        .clk(clock)
    );
    wire __T_282_ren3__q;
    wire __T_282_ren3__d;
    DFF_POSCLK #(.width(1)) _T_282_ren3 (
        .q(__T_282_ren3__q),
        .d(__T_282_ren3__d),
        .clk(clock)
    );
    wire __T_282_swap12__q;
    wire __T_282_swap12__d;
    DFF_POSCLK #(.width(1)) _T_282_swap12 (
        .q(__T_282_swap12__q),
        .d(__T_282_swap12__d),
        .clk(clock)
    );
    wire __T_282_swap23__q;
    wire __T_282_swap23__d;
    DFF_POSCLK #(.width(1)) _T_282_swap23 (
        .q(__T_282_swap23__q),
        .d(__T_282_swap23__d),
        .clk(clock)
    );
    wire __T_282_single__q;
    wire __T_282_single__d;
    DFF_POSCLK #(.width(1)) _T_282_single (
        .q(__T_282_single__q),
        .d(__T_282_single__d),
        .clk(clock)
    );
    wire __T_282_fromint__q;
    wire __T_282_fromint__d;
    DFF_POSCLK #(.width(1)) _T_282_fromint (
        .q(__T_282_fromint__q),
        .d(__T_282_fromint__d),
        .clk(clock)
    );
    wire __T_282_toint__q;
    wire __T_282_toint__d;
    DFF_POSCLK #(.width(1)) _T_282_toint (
        .q(__T_282_toint__q),
        .d(__T_282_toint__d),
        .clk(clock)
    );
    wire __T_282_fastpipe__q;
    wire __T_282_fastpipe__d;
    DFF_POSCLK #(.width(1)) _T_282_fastpipe (
        .q(__T_282_fastpipe__q),
        .d(__T_282_fastpipe__d),
        .clk(clock)
    );
    wire __T_282_fma__q;
    wire __T_282_fma__d;
    DFF_POSCLK #(.width(1)) _T_282_fma (
        .q(__T_282_fma__q),
        .d(__T_282_fma__d),
        .clk(clock)
    );
    wire __T_282_div__q;
    wire __T_282_div__d;
    DFF_POSCLK #(.width(1)) _T_282_div (
        .q(__T_282_div__q),
        .d(__T_282_div__d),
        .clk(clock)
    );
    wire __T_282_sqrt__q;
    wire __T_282_sqrt__d;
    DFF_POSCLK #(.width(1)) _T_282_sqrt (
        .q(__T_282_sqrt__q),
        .d(__T_282_sqrt__d),
        .clk(clock)
    );
    wire __T_282_wflags__q;
    wire __T_282_wflags__d;
    DFF_POSCLK #(.width(1)) _T_282_wflags (
        .q(__T_282_wflags__q),
        .d(__T_282_wflags__d),
        .clk(clock)
    );
    wire [4:0] ex_ctrl_cmd;
    MUX_UNSIGNED #(.width(5)) u_mux_122 (
        .y(ex_ctrl_cmd),
        .sel(ex_cp_valid),
        .a(cp_ctrl_cmd),
        .b(__T_282_cmd__q)
    );
    wire ex_ctrl_ldst;
    MUX_UNSIGNED #(.width(1)) u_mux_123 (
        .y(ex_ctrl_ldst),
        .sel(ex_cp_valid),
        .a(cp_ctrl_ldst),
        .b(__T_282_ldst__q)
    );
    wire ex_ctrl_wen;
    MUX_UNSIGNED #(.width(1)) u_mux_124 (
        .y(ex_ctrl_wen),
        .sel(ex_cp_valid),
        .a(cp_ctrl_wen),
        .b(__T_282_wen__q)
    );
    wire ex_ctrl_ren1;
    MUX_UNSIGNED #(.width(1)) u_mux_125 (
        .y(ex_ctrl_ren1),
        .sel(ex_cp_valid),
        .a(cp_ctrl_ren1),
        .b(__T_282_ren1__q)
    );
    wire ex_ctrl_ren2;
    MUX_UNSIGNED #(.width(1)) u_mux_126 (
        .y(ex_ctrl_ren2),
        .sel(ex_cp_valid),
        .a(cp_ctrl_ren2),
        .b(__T_282_ren2__q)
    );
    wire ex_ctrl_ren3;
    MUX_UNSIGNED #(.width(1)) u_mux_127 (
        .y(ex_ctrl_ren3),
        .sel(ex_cp_valid),
        .a(cp_ctrl_ren3),
        .b(__T_282_ren3__q)
    );
    wire ex_ctrl_swap12;
    MUX_UNSIGNED #(.width(1)) u_mux_128 (
        .y(ex_ctrl_swap12),
        .sel(ex_cp_valid),
        .a(cp_ctrl_swap12),
        .b(__T_282_swap12__q)
    );
    wire ex_ctrl_swap23;
    MUX_UNSIGNED #(.width(1)) u_mux_129 (
        .y(ex_ctrl_swap23),
        .sel(ex_cp_valid),
        .a(cp_ctrl_swap23),
        .b(__T_282_swap23__q)
    );
    wire ex_ctrl_single;
    MUX_UNSIGNED #(.width(1)) u_mux_130 (
        .y(ex_ctrl_single),
        .sel(ex_cp_valid),
        .a(cp_ctrl_single),
        .b(__T_282_single__q)
    );
    wire ex_ctrl_fromint;
    MUX_UNSIGNED #(.width(1)) u_mux_131 (
        .y(ex_ctrl_fromint),
        .sel(ex_cp_valid),
        .a(cp_ctrl_fromint),
        .b(__T_282_fromint__q)
    );
    wire ex_ctrl_toint;
    MUX_UNSIGNED #(.width(1)) u_mux_132 (
        .y(ex_ctrl_toint),
        .sel(ex_cp_valid),
        .a(cp_ctrl_toint),
        .b(__T_282_toint__q)
    );
    wire ex_ctrl_fastpipe;
    MUX_UNSIGNED #(.width(1)) u_mux_133 (
        .y(ex_ctrl_fastpipe),
        .sel(ex_cp_valid),
        .a(cp_ctrl_fastpipe),
        .b(__T_282_fastpipe__q)
    );
    wire ex_ctrl_fma;
    MUX_UNSIGNED #(.width(1)) u_mux_134 (
        .y(ex_ctrl_fma),
        .sel(ex_cp_valid),
        .a(cp_ctrl_fma),
        .b(__T_282_fma__q)
    );
    wire ex_ctrl_div;
    MUX_UNSIGNED #(.width(1)) u_mux_135 (
        .y(ex_ctrl_div),
        .sel(ex_cp_valid),
        .a(cp_ctrl_div),
        .b(__T_282_div__q)
    );
    wire ex_ctrl_sqrt;
    MUX_UNSIGNED #(.width(1)) u_mux_136 (
        .y(ex_ctrl_sqrt),
        .sel(ex_cp_valid),
        .a(cp_ctrl_sqrt),
        .b(__T_282_sqrt__q)
    );
    wire ex_ctrl_wflags;
    MUX_UNSIGNED #(.width(1)) u_mux_137 (
        .y(ex_ctrl_wflags),
        .sel(ex_cp_valid),
        .a(cp_ctrl_wflags),
        .b(__T_282_wflags__q)
    );
    wire [4:0] _mem_ctrl_cmd__q;
    wire [4:0] _mem_ctrl_cmd__d;
    DFF_POSCLK #(.width(5)) mem_ctrl_cmd (
        .q(_mem_ctrl_cmd__q),
        .d(_mem_ctrl_cmd__d),
        .clk(clock)
    );
    wire _mem_ctrl_ldst__q;
    wire _mem_ctrl_ldst__d;
    DFF_POSCLK #(.width(1)) mem_ctrl_ldst (
        .q(_mem_ctrl_ldst__q),
        .d(_mem_ctrl_ldst__d),
        .clk(clock)
    );
    wire _mem_ctrl_wen__q;
    wire _mem_ctrl_wen__d;
    DFF_POSCLK #(.width(1)) mem_ctrl_wen (
        .q(_mem_ctrl_wen__q),
        .d(_mem_ctrl_wen__d),
        .clk(clock)
    );
    wire _mem_ctrl_ren1__q;
    wire _mem_ctrl_ren1__d;
    DFF_POSCLK #(.width(1)) mem_ctrl_ren1 (
        .q(_mem_ctrl_ren1__q),
        .d(_mem_ctrl_ren1__d),
        .clk(clock)
    );
    wire _mem_ctrl_ren2__q;
    wire _mem_ctrl_ren2__d;
    DFF_POSCLK #(.width(1)) mem_ctrl_ren2 (
        .q(_mem_ctrl_ren2__q),
        .d(_mem_ctrl_ren2__d),
        .clk(clock)
    );
    wire _mem_ctrl_ren3__q;
    wire _mem_ctrl_ren3__d;
    DFF_POSCLK #(.width(1)) mem_ctrl_ren3 (
        .q(_mem_ctrl_ren3__q),
        .d(_mem_ctrl_ren3__d),
        .clk(clock)
    );
    wire _mem_ctrl_swap12__q;
    wire _mem_ctrl_swap12__d;
    DFF_POSCLK #(.width(1)) mem_ctrl_swap12 (
        .q(_mem_ctrl_swap12__q),
        .d(_mem_ctrl_swap12__d),
        .clk(clock)
    );
    wire _mem_ctrl_swap23__q;
    wire _mem_ctrl_swap23__d;
    DFF_POSCLK #(.width(1)) mem_ctrl_swap23 (
        .q(_mem_ctrl_swap23__q),
        .d(_mem_ctrl_swap23__d),
        .clk(clock)
    );
    wire _mem_ctrl_single__q;
    wire _mem_ctrl_single__d;
    DFF_POSCLK #(.width(1)) mem_ctrl_single (
        .q(_mem_ctrl_single__q),
        .d(_mem_ctrl_single__d),
        .clk(clock)
    );
    wire _mem_ctrl_fromint__q;
    wire _mem_ctrl_fromint__d;
    DFF_POSCLK #(.width(1)) mem_ctrl_fromint (
        .q(_mem_ctrl_fromint__q),
        .d(_mem_ctrl_fromint__d),
        .clk(clock)
    );
    wire _mem_ctrl_toint__q;
    wire _mem_ctrl_toint__d;
    DFF_POSCLK #(.width(1)) mem_ctrl_toint (
        .q(_mem_ctrl_toint__q),
        .d(_mem_ctrl_toint__d),
        .clk(clock)
    );
    wire _mem_ctrl_fastpipe__q;
    wire _mem_ctrl_fastpipe__d;
    DFF_POSCLK #(.width(1)) mem_ctrl_fastpipe (
        .q(_mem_ctrl_fastpipe__q),
        .d(_mem_ctrl_fastpipe__d),
        .clk(clock)
    );
    wire _mem_ctrl_fma__q;
    wire _mem_ctrl_fma__d;
    DFF_POSCLK #(.width(1)) mem_ctrl_fma (
        .q(_mem_ctrl_fma__q),
        .d(_mem_ctrl_fma__d),
        .clk(clock)
    );
    wire _mem_ctrl_div__q;
    wire _mem_ctrl_div__d;
    DFF_POSCLK #(.width(1)) mem_ctrl_div (
        .q(_mem_ctrl_div__q),
        .d(_mem_ctrl_div__d),
        .clk(clock)
    );
    wire _mem_ctrl_sqrt__q;
    wire _mem_ctrl_sqrt__d;
    DFF_POSCLK #(.width(1)) mem_ctrl_sqrt (
        .q(_mem_ctrl_sqrt__q),
        .d(_mem_ctrl_sqrt__d),
        .clk(clock)
    );
    wire _mem_ctrl_wflags__q;
    wire _mem_ctrl_wflags__d;
    DFF_POSCLK #(.width(1)) mem_ctrl_wflags (
        .q(_mem_ctrl_wflags__q),
        .d(_mem_ctrl_wflags__d),
        .clk(clock)
    );
    wire [4:0] _wb_ctrl_cmd__q;
    wire [4:0] _wb_ctrl_cmd__d;
    DFF_POSCLK #(.width(5)) wb_ctrl_cmd (
        .q(_wb_ctrl_cmd__q),
        .d(_wb_ctrl_cmd__d),
        .clk(clock)
    );
    wire _wb_ctrl_ldst__q;
    wire _wb_ctrl_ldst__d;
    DFF_POSCLK #(.width(1)) wb_ctrl_ldst (
        .q(_wb_ctrl_ldst__q),
        .d(_wb_ctrl_ldst__d),
        .clk(clock)
    );
    wire _wb_ctrl_wen__q;
    wire _wb_ctrl_wen__d;
    DFF_POSCLK #(.width(1)) wb_ctrl_wen (
        .q(_wb_ctrl_wen__q),
        .d(_wb_ctrl_wen__d),
        .clk(clock)
    );
    wire _wb_ctrl_ren1__q;
    wire _wb_ctrl_ren1__d;
    DFF_POSCLK #(.width(1)) wb_ctrl_ren1 (
        .q(_wb_ctrl_ren1__q),
        .d(_wb_ctrl_ren1__d),
        .clk(clock)
    );
    wire _wb_ctrl_ren2__q;
    wire _wb_ctrl_ren2__d;
    DFF_POSCLK #(.width(1)) wb_ctrl_ren2 (
        .q(_wb_ctrl_ren2__q),
        .d(_wb_ctrl_ren2__d),
        .clk(clock)
    );
    wire _wb_ctrl_ren3__q;
    wire _wb_ctrl_ren3__d;
    DFF_POSCLK #(.width(1)) wb_ctrl_ren3 (
        .q(_wb_ctrl_ren3__q),
        .d(_wb_ctrl_ren3__d),
        .clk(clock)
    );
    wire _wb_ctrl_swap12__q;
    wire _wb_ctrl_swap12__d;
    DFF_POSCLK #(.width(1)) wb_ctrl_swap12 (
        .q(_wb_ctrl_swap12__q),
        .d(_wb_ctrl_swap12__d),
        .clk(clock)
    );
    wire _wb_ctrl_swap23__q;
    wire _wb_ctrl_swap23__d;
    DFF_POSCLK #(.width(1)) wb_ctrl_swap23 (
        .q(_wb_ctrl_swap23__q),
        .d(_wb_ctrl_swap23__d),
        .clk(clock)
    );
    wire _wb_ctrl_single__q;
    wire _wb_ctrl_single__d;
    DFF_POSCLK #(.width(1)) wb_ctrl_single (
        .q(_wb_ctrl_single__q),
        .d(_wb_ctrl_single__d),
        .clk(clock)
    );
    wire _wb_ctrl_fromint__q;
    wire _wb_ctrl_fromint__d;
    DFF_POSCLK #(.width(1)) wb_ctrl_fromint (
        .q(_wb_ctrl_fromint__q),
        .d(_wb_ctrl_fromint__d),
        .clk(clock)
    );
    wire _wb_ctrl_toint__q;
    wire _wb_ctrl_toint__d;
    DFF_POSCLK #(.width(1)) wb_ctrl_toint (
        .q(_wb_ctrl_toint__q),
        .d(_wb_ctrl_toint__d),
        .clk(clock)
    );
    wire _wb_ctrl_fastpipe__q;
    wire _wb_ctrl_fastpipe__d;
    DFF_POSCLK #(.width(1)) wb_ctrl_fastpipe (
        .q(_wb_ctrl_fastpipe__q),
        .d(_wb_ctrl_fastpipe__d),
        .clk(clock)
    );
    wire _wb_ctrl_fma__q;
    wire _wb_ctrl_fma__d;
    DFF_POSCLK #(.width(1)) wb_ctrl_fma (
        .q(_wb_ctrl_fma__q),
        .d(_wb_ctrl_fma__d),
        .clk(clock)
    );
    wire _wb_ctrl_div__q;
    wire _wb_ctrl_div__d;
    DFF_POSCLK #(.width(1)) wb_ctrl_div (
        .q(_wb_ctrl_div__q),
        .d(_wb_ctrl_div__d),
        .clk(clock)
    );
    wire _wb_ctrl_sqrt__q;
    wire _wb_ctrl_sqrt__d;
    DFF_POSCLK #(.width(1)) wb_ctrl_sqrt (
        .q(_wb_ctrl_sqrt__q),
        .d(_wb_ctrl_sqrt__d),
        .clk(clock)
    );
    wire _wb_ctrl_wflags__q;
    wire _wb_ctrl_wflags__d;
    DFF_POSCLK #(.width(1)) wb_ctrl_wflags (
        .q(_wb_ctrl_wflags__q),
        .d(_wb_ctrl_wflags__d),
        .clk(clock)
    );
    wire _load_wb__q;
    wire _load_wb__d;
    DFF_POSCLK #(.width(1)) load_wb (
        .q(_load_wb__q),
        .d(_load_wb__d),
        .clk(clock)
    );
    wire _T_381;
    BITS #(.width(3), .high(0), .low(0)) bits_138 (
        .y(_T_381),
        .in(io_dmem_resp_type)
    );
    wire _T_383;
    EQ_UNSIGNED #(.width(1)) u_eq_139 (
        .y(_T_383),
        .a(_T_381),
        .b(1'h0)
    );
    wire _load_wb_single__q;
    wire _load_wb_single__d;
    DFF_POSCLK #(.width(1)) load_wb_single (
        .q(_load_wb_single__q),
        .d(_load_wb_single__d),
        .clk(clock)
    );
    wire [63:0] _load_wb_data__q;
    wire [63:0] _load_wb_data__d;
    DFF_POSCLK #(.width(64)) load_wb_data (
        .q(_load_wb_data__q),
        .d(_load_wb_data__d),
        .clk(clock)
    );
    wire [4:0] _load_wb_tag__q;
    wire [4:0] _load_wb_tag__d;
    DFF_POSCLK #(.width(5)) load_wb_tag (
        .q(_load_wb_tag__q),
        .d(_load_wb_tag__d),
        .clk(clock)
    );
    wire _T_387;
    BITS #(.width(64), .high(31), .low(31)) bits_140 (
        .y(_T_387),
        .in(_load_wb_data__q)
    );
    wire [7:0] _T_388;
    BITS #(.width(64), .high(30), .low(23)) bits_141 (
        .y(_T_388),
        .in(_load_wb_data__q)
    );
    wire [22:0] _T_389;
    BITS #(.width(64), .high(22), .low(0)) bits_142 (
        .y(_T_389),
        .in(_load_wb_data__q)
    );
    wire _T_391;
    wire [7:0] _WTEMP_5;
    PAD_UNSIGNED #(.width(1), .n(8)) u_pad_143 (
        .y(_WTEMP_5),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(8)) u_eq_144 (
        .y(_T_391),
        .a(_T_388),
        .b(_WTEMP_5)
    );
    wire _T_393;
    wire [22:0] _WTEMP_6;
    PAD_UNSIGNED #(.width(1), .n(23)) u_pad_145 (
        .y(_WTEMP_6),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(23)) u_eq_146 (
        .y(_T_393),
        .a(_T_389),
        .b(_WTEMP_6)
    );
    wire _T_394;
    BITWISEAND #(.width(1)) bitwiseand_147 (
        .y(_T_394),
        .a(_T_391),
        .b(_T_393)
    );
    wire [31:0] _T_395;
    SHL_UNSIGNED #(.width(23), .n(9)) u_shl_148 (
        .y(_T_395),
        .in(_T_389)
    );
    wire [15:0] _T_396;
    BITS #(.width(32), .high(31), .low(16)) bits_149 (
        .y(_T_396),
        .in(_T_395)
    );
    wire [15:0] _T_397;
    BITS #(.width(32), .high(15), .low(0)) bits_150 (
        .y(_T_397),
        .in(_T_395)
    );
    wire _T_399;
    wire [15:0] _WTEMP_7;
    PAD_UNSIGNED #(.width(1), .n(16)) u_pad_151 (
        .y(_WTEMP_7),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(16)) u_neq_152 (
        .y(_T_399),
        .a(_T_396),
        .b(_WTEMP_7)
    );
    wire [7:0] _T_400;
    BITS #(.width(16), .high(15), .low(8)) bits_153 (
        .y(_T_400),
        .in(_T_396)
    );
    wire [7:0] _T_401;
    BITS #(.width(16), .high(7), .low(0)) bits_154 (
        .y(_T_401),
        .in(_T_396)
    );
    wire _T_403;
    wire [7:0] _WTEMP_8;
    PAD_UNSIGNED #(.width(1), .n(8)) u_pad_155 (
        .y(_WTEMP_8),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(8)) u_neq_156 (
        .y(_T_403),
        .a(_T_400),
        .b(_WTEMP_8)
    );
    wire [3:0] _T_404;
    BITS #(.width(8), .high(7), .low(4)) bits_157 (
        .y(_T_404),
        .in(_T_400)
    );
    wire [3:0] _T_405;
    BITS #(.width(8), .high(3), .low(0)) bits_158 (
        .y(_T_405),
        .in(_T_400)
    );
    wire _T_407;
    wire [3:0] _WTEMP_9;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_159 (
        .y(_WTEMP_9),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_160 (
        .y(_T_407),
        .a(_T_404),
        .b(_WTEMP_9)
    );
    wire _T_408;
    BITS #(.width(4), .high(3), .low(3)) bits_161 (
        .y(_T_408),
        .in(_T_404)
    );
    wire _T_410;
    BITS #(.width(4), .high(2), .low(2)) bits_162 (
        .y(_T_410),
        .in(_T_404)
    );
    wire _T_412;
    BITS #(.width(4), .high(1), .low(1)) bits_163 (
        .y(_T_412),
        .in(_T_404)
    );
    wire [1:0] _T_413;
    wire [1:0] _WTEMP_10;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_164 (
        .y(_WTEMP_10),
        .in(_T_412)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_165 (
        .y(_T_413),
        .sel(_T_410),
        .a(2'h2),
        .b(_WTEMP_10)
    );
    wire [1:0] _T_414;
    MUX_UNSIGNED #(.width(2)) u_mux_166 (
        .y(_T_414),
        .sel(_T_408),
        .a(2'h3),
        .b(_T_413)
    );
    wire _T_415;
    BITS #(.width(4), .high(3), .low(3)) bits_167 (
        .y(_T_415),
        .in(_T_405)
    );
    wire _T_417;
    BITS #(.width(4), .high(2), .low(2)) bits_168 (
        .y(_T_417),
        .in(_T_405)
    );
    wire _T_419;
    BITS #(.width(4), .high(1), .low(1)) bits_169 (
        .y(_T_419),
        .in(_T_405)
    );
    wire [1:0] _T_420;
    wire [1:0] _WTEMP_11;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_170 (
        .y(_WTEMP_11),
        .in(_T_419)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_171 (
        .y(_T_420),
        .sel(_T_417),
        .a(2'h2),
        .b(_WTEMP_11)
    );
    wire [1:0] _T_421;
    MUX_UNSIGNED #(.width(2)) u_mux_172 (
        .y(_T_421),
        .sel(_T_415),
        .a(2'h3),
        .b(_T_420)
    );
    wire [1:0] _T_422;
    MUX_UNSIGNED #(.width(2)) u_mux_173 (
        .y(_T_422),
        .sel(_T_407),
        .a(_T_414),
        .b(_T_421)
    );
    wire [2:0] _T_423;
    CAT #(.width_a(1), .width_b(2)) cat_174 (
        .y(_T_423),
        .a(_T_407),
        .b(_T_422)
    );
    wire [3:0] _T_424;
    BITS #(.width(8), .high(7), .low(4)) bits_175 (
        .y(_T_424),
        .in(_T_401)
    );
    wire [3:0] _T_425;
    BITS #(.width(8), .high(3), .low(0)) bits_176 (
        .y(_T_425),
        .in(_T_401)
    );
    wire _T_427;
    wire [3:0] _WTEMP_12;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_177 (
        .y(_WTEMP_12),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_178 (
        .y(_T_427),
        .a(_T_424),
        .b(_WTEMP_12)
    );
    wire _T_428;
    BITS #(.width(4), .high(3), .low(3)) bits_179 (
        .y(_T_428),
        .in(_T_424)
    );
    wire _T_430;
    BITS #(.width(4), .high(2), .low(2)) bits_180 (
        .y(_T_430),
        .in(_T_424)
    );
    wire _T_432;
    BITS #(.width(4), .high(1), .low(1)) bits_181 (
        .y(_T_432),
        .in(_T_424)
    );
    wire [1:0] _T_433;
    wire [1:0] _WTEMP_13;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_182 (
        .y(_WTEMP_13),
        .in(_T_432)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_183 (
        .y(_T_433),
        .sel(_T_430),
        .a(2'h2),
        .b(_WTEMP_13)
    );
    wire [1:0] _T_434;
    MUX_UNSIGNED #(.width(2)) u_mux_184 (
        .y(_T_434),
        .sel(_T_428),
        .a(2'h3),
        .b(_T_433)
    );
    wire _T_435;
    BITS #(.width(4), .high(3), .low(3)) bits_185 (
        .y(_T_435),
        .in(_T_425)
    );
    wire _T_437;
    BITS #(.width(4), .high(2), .low(2)) bits_186 (
        .y(_T_437),
        .in(_T_425)
    );
    wire _T_439;
    BITS #(.width(4), .high(1), .low(1)) bits_187 (
        .y(_T_439),
        .in(_T_425)
    );
    wire [1:0] _T_440;
    wire [1:0] _WTEMP_14;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_188 (
        .y(_WTEMP_14),
        .in(_T_439)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_189 (
        .y(_T_440),
        .sel(_T_437),
        .a(2'h2),
        .b(_WTEMP_14)
    );
    wire [1:0] _T_441;
    MUX_UNSIGNED #(.width(2)) u_mux_190 (
        .y(_T_441),
        .sel(_T_435),
        .a(2'h3),
        .b(_T_440)
    );
    wire [1:0] _T_442;
    MUX_UNSIGNED #(.width(2)) u_mux_191 (
        .y(_T_442),
        .sel(_T_427),
        .a(_T_434),
        .b(_T_441)
    );
    wire [2:0] _T_443;
    CAT #(.width_a(1), .width_b(2)) cat_192 (
        .y(_T_443),
        .a(_T_427),
        .b(_T_442)
    );
    wire [2:0] _T_444;
    MUX_UNSIGNED #(.width(3)) u_mux_193 (
        .y(_T_444),
        .sel(_T_403),
        .a(_T_423),
        .b(_T_443)
    );
    wire [3:0] _T_445;
    CAT #(.width_a(1), .width_b(3)) cat_194 (
        .y(_T_445),
        .a(_T_403),
        .b(_T_444)
    );
    wire [7:0] _T_446;
    BITS #(.width(16), .high(15), .low(8)) bits_195 (
        .y(_T_446),
        .in(_T_397)
    );
    wire [7:0] _T_447;
    BITS #(.width(16), .high(7), .low(0)) bits_196 (
        .y(_T_447),
        .in(_T_397)
    );
    wire _T_449;
    wire [7:0] _WTEMP_15;
    PAD_UNSIGNED #(.width(1), .n(8)) u_pad_197 (
        .y(_WTEMP_15),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(8)) u_neq_198 (
        .y(_T_449),
        .a(_T_446),
        .b(_WTEMP_15)
    );
    wire [3:0] _T_450;
    BITS #(.width(8), .high(7), .low(4)) bits_199 (
        .y(_T_450),
        .in(_T_446)
    );
    wire [3:0] _T_451;
    BITS #(.width(8), .high(3), .low(0)) bits_200 (
        .y(_T_451),
        .in(_T_446)
    );
    wire _T_453;
    wire [3:0] _WTEMP_16;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_201 (
        .y(_WTEMP_16),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_202 (
        .y(_T_453),
        .a(_T_450),
        .b(_WTEMP_16)
    );
    wire _T_454;
    BITS #(.width(4), .high(3), .low(3)) bits_203 (
        .y(_T_454),
        .in(_T_450)
    );
    wire _T_456;
    BITS #(.width(4), .high(2), .low(2)) bits_204 (
        .y(_T_456),
        .in(_T_450)
    );
    wire _T_458;
    BITS #(.width(4), .high(1), .low(1)) bits_205 (
        .y(_T_458),
        .in(_T_450)
    );
    wire [1:0] _T_459;
    wire [1:0] _WTEMP_17;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_206 (
        .y(_WTEMP_17),
        .in(_T_458)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_207 (
        .y(_T_459),
        .sel(_T_456),
        .a(2'h2),
        .b(_WTEMP_17)
    );
    wire [1:0] _T_460;
    MUX_UNSIGNED #(.width(2)) u_mux_208 (
        .y(_T_460),
        .sel(_T_454),
        .a(2'h3),
        .b(_T_459)
    );
    wire _T_461;
    BITS #(.width(4), .high(3), .low(3)) bits_209 (
        .y(_T_461),
        .in(_T_451)
    );
    wire _T_463;
    BITS #(.width(4), .high(2), .low(2)) bits_210 (
        .y(_T_463),
        .in(_T_451)
    );
    wire _T_465;
    BITS #(.width(4), .high(1), .low(1)) bits_211 (
        .y(_T_465),
        .in(_T_451)
    );
    wire [1:0] _T_466;
    wire [1:0] _WTEMP_18;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_212 (
        .y(_WTEMP_18),
        .in(_T_465)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_213 (
        .y(_T_466),
        .sel(_T_463),
        .a(2'h2),
        .b(_WTEMP_18)
    );
    wire [1:0] _T_467;
    MUX_UNSIGNED #(.width(2)) u_mux_214 (
        .y(_T_467),
        .sel(_T_461),
        .a(2'h3),
        .b(_T_466)
    );
    wire [1:0] _T_468;
    MUX_UNSIGNED #(.width(2)) u_mux_215 (
        .y(_T_468),
        .sel(_T_453),
        .a(_T_460),
        .b(_T_467)
    );
    wire [2:0] _T_469;
    CAT #(.width_a(1), .width_b(2)) cat_216 (
        .y(_T_469),
        .a(_T_453),
        .b(_T_468)
    );
    wire [3:0] _T_470;
    BITS #(.width(8), .high(7), .low(4)) bits_217 (
        .y(_T_470),
        .in(_T_447)
    );
    wire [3:0] _T_471;
    BITS #(.width(8), .high(3), .low(0)) bits_218 (
        .y(_T_471),
        .in(_T_447)
    );
    wire _T_473;
    wire [3:0] _WTEMP_19;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_219 (
        .y(_WTEMP_19),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_220 (
        .y(_T_473),
        .a(_T_470),
        .b(_WTEMP_19)
    );
    wire _T_474;
    BITS #(.width(4), .high(3), .low(3)) bits_221 (
        .y(_T_474),
        .in(_T_470)
    );
    wire _T_476;
    BITS #(.width(4), .high(2), .low(2)) bits_222 (
        .y(_T_476),
        .in(_T_470)
    );
    wire _T_478;
    BITS #(.width(4), .high(1), .low(1)) bits_223 (
        .y(_T_478),
        .in(_T_470)
    );
    wire [1:0] _T_479;
    wire [1:0] _WTEMP_20;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_224 (
        .y(_WTEMP_20),
        .in(_T_478)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_225 (
        .y(_T_479),
        .sel(_T_476),
        .a(2'h2),
        .b(_WTEMP_20)
    );
    wire [1:0] _T_480;
    MUX_UNSIGNED #(.width(2)) u_mux_226 (
        .y(_T_480),
        .sel(_T_474),
        .a(2'h3),
        .b(_T_479)
    );
    wire _T_481;
    BITS #(.width(4), .high(3), .low(3)) bits_227 (
        .y(_T_481),
        .in(_T_471)
    );
    wire _T_483;
    BITS #(.width(4), .high(2), .low(2)) bits_228 (
        .y(_T_483),
        .in(_T_471)
    );
    wire _T_485;
    BITS #(.width(4), .high(1), .low(1)) bits_229 (
        .y(_T_485),
        .in(_T_471)
    );
    wire [1:0] _T_486;
    wire [1:0] _WTEMP_21;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_230 (
        .y(_WTEMP_21),
        .in(_T_485)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_231 (
        .y(_T_486),
        .sel(_T_483),
        .a(2'h2),
        .b(_WTEMP_21)
    );
    wire [1:0] _T_487;
    MUX_UNSIGNED #(.width(2)) u_mux_232 (
        .y(_T_487),
        .sel(_T_481),
        .a(2'h3),
        .b(_T_486)
    );
    wire [1:0] _T_488;
    MUX_UNSIGNED #(.width(2)) u_mux_233 (
        .y(_T_488),
        .sel(_T_473),
        .a(_T_480),
        .b(_T_487)
    );
    wire [2:0] _T_489;
    CAT #(.width_a(1), .width_b(2)) cat_234 (
        .y(_T_489),
        .a(_T_473),
        .b(_T_488)
    );
    wire [2:0] _T_490;
    MUX_UNSIGNED #(.width(3)) u_mux_235 (
        .y(_T_490),
        .sel(_T_449),
        .a(_T_469),
        .b(_T_489)
    );
    wire [3:0] _T_491;
    CAT #(.width_a(1), .width_b(3)) cat_236 (
        .y(_T_491),
        .a(_T_449),
        .b(_T_490)
    );
    wire [3:0] _T_492;
    MUX_UNSIGNED #(.width(4)) u_mux_237 (
        .y(_T_492),
        .sel(_T_399),
        .a(_T_445),
        .b(_T_491)
    );
    wire [4:0] _T_493;
    CAT #(.width_a(1), .width_b(4)) cat_238 (
        .y(_T_493),
        .a(_T_399),
        .b(_T_492)
    );
    wire [4:0] _T_494;
    BITWISENOT #(.width(5)) bitwisenot_239 (
        .y(_T_494),
        .in(_T_493)
    );
    wire [53:0] _T_495;
    DSHL_UNSIGNED #(.width_in(23), .width_n(5)) u_dshl_240 (
        .y(_T_495),
        .in(_T_389),
        .n(_T_494)
    );
    wire [21:0] _T_496;
    BITS #(.width(54), .high(21), .low(0)) bits_241 (
        .y(_T_496),
        .in(_T_495)
    );
    wire [22:0] _T_498;
    CAT #(.width_a(22), .width_b(1)) cat_242 (
        .y(_T_498),
        .a(_T_496),
        .b(1'h0)
    );
    wire [8:0] _T_503;
    assign _T_503 = 9'h1FF;
    wire [8:0] _T_504;
    wire [8:0] _WTEMP_22;
    PAD_UNSIGNED #(.width(5), .n(9)) u_pad_243 (
        .y(_WTEMP_22),
        .in(_T_494)
    );
    BITWISEXOR #(.width(9)) bitwisexor_244 (
        .y(_T_504),
        .a(_WTEMP_22),
        .b(_T_503)
    );
    wire [8:0] _T_505;
    wire [8:0] _WTEMP_23;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_245 (
        .y(_WTEMP_23),
        .in(_T_388)
    );
    MUX_UNSIGNED #(.width(9)) u_mux_246 (
        .y(_T_505),
        .sel(_T_391),
        .a(_T_504),
        .b(_WTEMP_23)
    );
    wire [1:0] _T_509;
    wire [1:0] _WTEMP_24;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_247 (
        .y(_WTEMP_24),
        .in(1'h1)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_248 (
        .y(_T_509),
        .sel(_T_391),
        .a(2'h2),
        .b(_WTEMP_24)
    );
    wire [7:0] _T_510;
    wire [7:0] _WTEMP_25;
    PAD_UNSIGNED #(.width(2), .n(8)) u_pad_249 (
        .y(_WTEMP_25),
        .in(_T_509)
    );
    BITWISEOR #(.width(8)) bitwiseor_250 (
        .y(_T_510),
        .a(8'h80),
        .b(_WTEMP_25)
    );
    wire [9:0] _T_511;
    wire [8:0] _WTEMP_26;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_251 (
        .y(_WTEMP_26),
        .in(_T_510)
    );
    ADD_UNSIGNED #(.width(9)) u_add_252 (
        .y(_T_511),
        .a(_T_505),
        .b(_WTEMP_26)
    );
    wire [8:0] _T_512;
    TAIL #(.width(10), .n(1)) tail_253 (
        .y(_T_512),
        .in(_T_511)
    );
    wire [1:0] _T_513;
    BITS #(.width(9), .high(8), .low(7)) bits_254 (
        .y(_T_513),
        .in(_T_512)
    );
    wire _T_515;
    EQ_UNSIGNED #(.width(2)) u_eq_255 (
        .y(_T_515),
        .a(_T_513),
        .b(2'h3)
    );
    wire _T_517;
    EQ_UNSIGNED #(.width(1)) u_eq_256 (
        .y(_T_517),
        .a(_T_393),
        .b(1'h0)
    );
    wire _T_518;
    BITWISEAND #(.width(1)) bitwiseand_257 (
        .y(_T_518),
        .a(_T_515),
        .b(_T_517)
    );
    wire _T_519;
    BITS #(.width(1), .high(0), .low(0)) bits_258 (
        .y(_T_519),
        .in(_T_394)
    );
    wire [2:0] _T_522;
    MUX_UNSIGNED #(.width(3)) u_mux_259 (
        .y(_T_522),
        .sel(_T_519),
        .a(3'h7),
        .b(3'h0)
    );
    wire [8:0] _T_523;
    SHL_UNSIGNED #(.width(3), .n(6)) u_shl_260 (
        .y(_T_523),
        .in(_T_522)
    );
    wire [8:0] _T_524;
    BITWISENOT #(.width(9)) bitwisenot_261 (
        .y(_T_524),
        .in(_T_523)
    );
    wire [8:0] _T_525;
    BITWISEAND #(.width(9)) bitwiseand_262 (
        .y(_T_525),
        .a(_T_512),
        .b(_T_524)
    );
    wire [6:0] _T_526;
    SHL_UNSIGNED #(.width(1), .n(6)) u_shl_263 (
        .y(_T_526),
        .in(_T_518)
    );
    wire [8:0] _T_527;
    wire [8:0] _WTEMP_27;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_264 (
        .y(_WTEMP_27),
        .in(_T_526)
    );
    BITWISEOR #(.width(9)) bitwiseor_265 (
        .y(_T_527),
        .a(_T_525),
        .b(_WTEMP_27)
    );
    wire [22:0] _T_528;
    MUX_UNSIGNED #(.width(23)) u_mux_266 (
        .y(_T_528),
        .sel(_T_391),
        .a(_T_498),
        .b(_T_389)
    );
    wire [9:0] _T_529;
    CAT #(.width_a(1), .width_b(9)) cat_267 (
        .y(_T_529),
        .a(_T_387),
        .b(_T_527)
    );
    wire [32:0] rec_s;
    CAT #(.width_a(10), .width_b(23)) cat_268 (
        .y(rec_s),
        .a(_T_529),
        .b(_T_528)
    );
    wire _T_530;
    BITS #(.width(64), .high(63), .low(63)) bits_269 (
        .y(_T_530),
        .in(_load_wb_data__q)
    );
    wire [10:0] _T_531;
    BITS #(.width(64), .high(62), .low(52)) bits_270 (
        .y(_T_531),
        .in(_load_wb_data__q)
    );
    wire [51:0] _T_532;
    BITS #(.width(64), .high(51), .low(0)) bits_271 (
        .y(_T_532),
        .in(_load_wb_data__q)
    );
    wire _T_534;
    wire [10:0] _WTEMP_28;
    PAD_UNSIGNED #(.width(1), .n(11)) u_pad_272 (
        .y(_WTEMP_28),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(11)) u_eq_273 (
        .y(_T_534),
        .a(_T_531),
        .b(_WTEMP_28)
    );
    wire _T_536;
    wire [51:0] _WTEMP_29;
    PAD_UNSIGNED #(.width(1), .n(52)) u_pad_274 (
        .y(_WTEMP_29),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(52)) u_eq_275 (
        .y(_T_536),
        .a(_T_532),
        .b(_WTEMP_29)
    );
    wire _T_537;
    BITWISEAND #(.width(1)) bitwiseand_276 (
        .y(_T_537),
        .a(_T_534),
        .b(_T_536)
    );
    wire [63:0] _T_538;
    SHL_UNSIGNED #(.width(52), .n(12)) u_shl_277 (
        .y(_T_538),
        .in(_T_532)
    );
    wire [31:0] _T_539;
    BITS #(.width(64), .high(63), .low(32)) bits_278 (
        .y(_T_539),
        .in(_T_538)
    );
    wire [31:0] _T_540;
    BITS #(.width(64), .high(31), .low(0)) bits_279 (
        .y(_T_540),
        .in(_T_538)
    );
    wire _T_542;
    wire [31:0] _WTEMP_30;
    PAD_UNSIGNED #(.width(1), .n(32)) u_pad_280 (
        .y(_WTEMP_30),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(32)) u_neq_281 (
        .y(_T_542),
        .a(_T_539),
        .b(_WTEMP_30)
    );
    wire [15:0] _T_543;
    BITS #(.width(32), .high(31), .low(16)) bits_282 (
        .y(_T_543),
        .in(_T_539)
    );
    wire [15:0] _T_544;
    BITS #(.width(32), .high(15), .low(0)) bits_283 (
        .y(_T_544),
        .in(_T_539)
    );
    wire _T_546;
    wire [15:0] _WTEMP_31;
    PAD_UNSIGNED #(.width(1), .n(16)) u_pad_284 (
        .y(_WTEMP_31),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(16)) u_neq_285 (
        .y(_T_546),
        .a(_T_543),
        .b(_WTEMP_31)
    );
    wire [7:0] _T_547;
    BITS #(.width(16), .high(15), .low(8)) bits_286 (
        .y(_T_547),
        .in(_T_543)
    );
    wire [7:0] _T_548;
    BITS #(.width(16), .high(7), .low(0)) bits_287 (
        .y(_T_548),
        .in(_T_543)
    );
    wire _T_550;
    wire [7:0] _WTEMP_32;
    PAD_UNSIGNED #(.width(1), .n(8)) u_pad_288 (
        .y(_WTEMP_32),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(8)) u_neq_289 (
        .y(_T_550),
        .a(_T_547),
        .b(_WTEMP_32)
    );
    wire [3:0] _T_551;
    BITS #(.width(8), .high(7), .low(4)) bits_290 (
        .y(_T_551),
        .in(_T_547)
    );
    wire [3:0] _T_552;
    BITS #(.width(8), .high(3), .low(0)) bits_291 (
        .y(_T_552),
        .in(_T_547)
    );
    wire _T_554;
    wire [3:0] _WTEMP_33;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_292 (
        .y(_WTEMP_33),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_293 (
        .y(_T_554),
        .a(_T_551),
        .b(_WTEMP_33)
    );
    wire _T_555;
    BITS #(.width(4), .high(3), .low(3)) bits_294 (
        .y(_T_555),
        .in(_T_551)
    );
    wire _T_557;
    BITS #(.width(4), .high(2), .low(2)) bits_295 (
        .y(_T_557),
        .in(_T_551)
    );
    wire _T_559;
    BITS #(.width(4), .high(1), .low(1)) bits_296 (
        .y(_T_559),
        .in(_T_551)
    );
    wire [1:0] _T_560;
    wire [1:0] _WTEMP_34;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_297 (
        .y(_WTEMP_34),
        .in(_T_559)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_298 (
        .y(_T_560),
        .sel(_T_557),
        .a(2'h2),
        .b(_WTEMP_34)
    );
    wire [1:0] _T_561;
    MUX_UNSIGNED #(.width(2)) u_mux_299 (
        .y(_T_561),
        .sel(_T_555),
        .a(2'h3),
        .b(_T_560)
    );
    wire _T_562;
    BITS #(.width(4), .high(3), .low(3)) bits_300 (
        .y(_T_562),
        .in(_T_552)
    );
    wire _T_564;
    BITS #(.width(4), .high(2), .low(2)) bits_301 (
        .y(_T_564),
        .in(_T_552)
    );
    wire _T_566;
    BITS #(.width(4), .high(1), .low(1)) bits_302 (
        .y(_T_566),
        .in(_T_552)
    );
    wire [1:0] _T_567;
    wire [1:0] _WTEMP_35;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_303 (
        .y(_WTEMP_35),
        .in(_T_566)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_304 (
        .y(_T_567),
        .sel(_T_564),
        .a(2'h2),
        .b(_WTEMP_35)
    );
    wire [1:0] _T_568;
    MUX_UNSIGNED #(.width(2)) u_mux_305 (
        .y(_T_568),
        .sel(_T_562),
        .a(2'h3),
        .b(_T_567)
    );
    wire [1:0] _T_569;
    MUX_UNSIGNED #(.width(2)) u_mux_306 (
        .y(_T_569),
        .sel(_T_554),
        .a(_T_561),
        .b(_T_568)
    );
    wire [2:0] _T_570;
    CAT #(.width_a(1), .width_b(2)) cat_307 (
        .y(_T_570),
        .a(_T_554),
        .b(_T_569)
    );
    wire [3:0] _T_571;
    BITS #(.width(8), .high(7), .low(4)) bits_308 (
        .y(_T_571),
        .in(_T_548)
    );
    wire [3:0] _T_572;
    BITS #(.width(8), .high(3), .low(0)) bits_309 (
        .y(_T_572),
        .in(_T_548)
    );
    wire _T_574;
    wire [3:0] _WTEMP_36;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_310 (
        .y(_WTEMP_36),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_311 (
        .y(_T_574),
        .a(_T_571),
        .b(_WTEMP_36)
    );
    wire _T_575;
    BITS #(.width(4), .high(3), .low(3)) bits_312 (
        .y(_T_575),
        .in(_T_571)
    );
    wire _T_577;
    BITS #(.width(4), .high(2), .low(2)) bits_313 (
        .y(_T_577),
        .in(_T_571)
    );
    wire _T_579;
    BITS #(.width(4), .high(1), .low(1)) bits_314 (
        .y(_T_579),
        .in(_T_571)
    );
    wire [1:0] _T_580;
    wire [1:0] _WTEMP_37;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_315 (
        .y(_WTEMP_37),
        .in(_T_579)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_316 (
        .y(_T_580),
        .sel(_T_577),
        .a(2'h2),
        .b(_WTEMP_37)
    );
    wire [1:0] _T_581;
    MUX_UNSIGNED #(.width(2)) u_mux_317 (
        .y(_T_581),
        .sel(_T_575),
        .a(2'h3),
        .b(_T_580)
    );
    wire _T_582;
    BITS #(.width(4), .high(3), .low(3)) bits_318 (
        .y(_T_582),
        .in(_T_572)
    );
    wire _T_584;
    BITS #(.width(4), .high(2), .low(2)) bits_319 (
        .y(_T_584),
        .in(_T_572)
    );
    wire _T_586;
    BITS #(.width(4), .high(1), .low(1)) bits_320 (
        .y(_T_586),
        .in(_T_572)
    );
    wire [1:0] _T_587;
    wire [1:0] _WTEMP_38;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_321 (
        .y(_WTEMP_38),
        .in(_T_586)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_322 (
        .y(_T_587),
        .sel(_T_584),
        .a(2'h2),
        .b(_WTEMP_38)
    );
    wire [1:0] _T_588;
    MUX_UNSIGNED #(.width(2)) u_mux_323 (
        .y(_T_588),
        .sel(_T_582),
        .a(2'h3),
        .b(_T_587)
    );
    wire [1:0] _T_589;
    MUX_UNSIGNED #(.width(2)) u_mux_324 (
        .y(_T_589),
        .sel(_T_574),
        .a(_T_581),
        .b(_T_588)
    );
    wire [2:0] _T_590;
    CAT #(.width_a(1), .width_b(2)) cat_325 (
        .y(_T_590),
        .a(_T_574),
        .b(_T_589)
    );
    wire [2:0] _T_591;
    MUX_UNSIGNED #(.width(3)) u_mux_326 (
        .y(_T_591),
        .sel(_T_550),
        .a(_T_570),
        .b(_T_590)
    );
    wire [3:0] _T_592;
    CAT #(.width_a(1), .width_b(3)) cat_327 (
        .y(_T_592),
        .a(_T_550),
        .b(_T_591)
    );
    wire [7:0] _T_593;
    BITS #(.width(16), .high(15), .low(8)) bits_328 (
        .y(_T_593),
        .in(_T_544)
    );
    wire [7:0] _T_594;
    BITS #(.width(16), .high(7), .low(0)) bits_329 (
        .y(_T_594),
        .in(_T_544)
    );
    wire _T_596;
    wire [7:0] _WTEMP_39;
    PAD_UNSIGNED #(.width(1), .n(8)) u_pad_330 (
        .y(_WTEMP_39),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(8)) u_neq_331 (
        .y(_T_596),
        .a(_T_593),
        .b(_WTEMP_39)
    );
    wire [3:0] _T_597;
    BITS #(.width(8), .high(7), .low(4)) bits_332 (
        .y(_T_597),
        .in(_T_593)
    );
    wire [3:0] _T_598;
    BITS #(.width(8), .high(3), .low(0)) bits_333 (
        .y(_T_598),
        .in(_T_593)
    );
    wire _T_600;
    wire [3:0] _WTEMP_40;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_334 (
        .y(_WTEMP_40),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_335 (
        .y(_T_600),
        .a(_T_597),
        .b(_WTEMP_40)
    );
    wire _T_601;
    BITS #(.width(4), .high(3), .low(3)) bits_336 (
        .y(_T_601),
        .in(_T_597)
    );
    wire _T_603;
    BITS #(.width(4), .high(2), .low(2)) bits_337 (
        .y(_T_603),
        .in(_T_597)
    );
    wire _T_605;
    BITS #(.width(4), .high(1), .low(1)) bits_338 (
        .y(_T_605),
        .in(_T_597)
    );
    wire [1:0] _T_606;
    wire [1:0] _WTEMP_41;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_339 (
        .y(_WTEMP_41),
        .in(_T_605)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_340 (
        .y(_T_606),
        .sel(_T_603),
        .a(2'h2),
        .b(_WTEMP_41)
    );
    wire [1:0] _T_607;
    MUX_UNSIGNED #(.width(2)) u_mux_341 (
        .y(_T_607),
        .sel(_T_601),
        .a(2'h3),
        .b(_T_606)
    );
    wire _T_608;
    BITS #(.width(4), .high(3), .low(3)) bits_342 (
        .y(_T_608),
        .in(_T_598)
    );
    wire _T_610;
    BITS #(.width(4), .high(2), .low(2)) bits_343 (
        .y(_T_610),
        .in(_T_598)
    );
    wire _T_612;
    BITS #(.width(4), .high(1), .low(1)) bits_344 (
        .y(_T_612),
        .in(_T_598)
    );
    wire [1:0] _T_613;
    wire [1:0] _WTEMP_42;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_345 (
        .y(_WTEMP_42),
        .in(_T_612)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_346 (
        .y(_T_613),
        .sel(_T_610),
        .a(2'h2),
        .b(_WTEMP_42)
    );
    wire [1:0] _T_614;
    MUX_UNSIGNED #(.width(2)) u_mux_347 (
        .y(_T_614),
        .sel(_T_608),
        .a(2'h3),
        .b(_T_613)
    );
    wire [1:0] _T_615;
    MUX_UNSIGNED #(.width(2)) u_mux_348 (
        .y(_T_615),
        .sel(_T_600),
        .a(_T_607),
        .b(_T_614)
    );
    wire [2:0] _T_616;
    CAT #(.width_a(1), .width_b(2)) cat_349 (
        .y(_T_616),
        .a(_T_600),
        .b(_T_615)
    );
    wire [3:0] _T_617;
    BITS #(.width(8), .high(7), .low(4)) bits_350 (
        .y(_T_617),
        .in(_T_594)
    );
    wire [3:0] _T_618;
    BITS #(.width(8), .high(3), .low(0)) bits_351 (
        .y(_T_618),
        .in(_T_594)
    );
    wire _T_620;
    wire [3:0] _WTEMP_43;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_352 (
        .y(_WTEMP_43),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_353 (
        .y(_T_620),
        .a(_T_617),
        .b(_WTEMP_43)
    );
    wire _T_621;
    BITS #(.width(4), .high(3), .low(3)) bits_354 (
        .y(_T_621),
        .in(_T_617)
    );
    wire _T_623;
    BITS #(.width(4), .high(2), .low(2)) bits_355 (
        .y(_T_623),
        .in(_T_617)
    );
    wire _T_625;
    BITS #(.width(4), .high(1), .low(1)) bits_356 (
        .y(_T_625),
        .in(_T_617)
    );
    wire [1:0] _T_626;
    wire [1:0] _WTEMP_44;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_357 (
        .y(_WTEMP_44),
        .in(_T_625)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_358 (
        .y(_T_626),
        .sel(_T_623),
        .a(2'h2),
        .b(_WTEMP_44)
    );
    wire [1:0] _T_627;
    MUX_UNSIGNED #(.width(2)) u_mux_359 (
        .y(_T_627),
        .sel(_T_621),
        .a(2'h3),
        .b(_T_626)
    );
    wire _T_628;
    BITS #(.width(4), .high(3), .low(3)) bits_360 (
        .y(_T_628),
        .in(_T_618)
    );
    wire _T_630;
    BITS #(.width(4), .high(2), .low(2)) bits_361 (
        .y(_T_630),
        .in(_T_618)
    );
    wire _T_632;
    BITS #(.width(4), .high(1), .low(1)) bits_362 (
        .y(_T_632),
        .in(_T_618)
    );
    wire [1:0] _T_633;
    wire [1:0] _WTEMP_45;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_363 (
        .y(_WTEMP_45),
        .in(_T_632)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_364 (
        .y(_T_633),
        .sel(_T_630),
        .a(2'h2),
        .b(_WTEMP_45)
    );
    wire [1:0] _T_634;
    MUX_UNSIGNED #(.width(2)) u_mux_365 (
        .y(_T_634),
        .sel(_T_628),
        .a(2'h3),
        .b(_T_633)
    );
    wire [1:0] _T_635;
    MUX_UNSIGNED #(.width(2)) u_mux_366 (
        .y(_T_635),
        .sel(_T_620),
        .a(_T_627),
        .b(_T_634)
    );
    wire [2:0] _T_636;
    CAT #(.width_a(1), .width_b(2)) cat_367 (
        .y(_T_636),
        .a(_T_620),
        .b(_T_635)
    );
    wire [2:0] _T_637;
    MUX_UNSIGNED #(.width(3)) u_mux_368 (
        .y(_T_637),
        .sel(_T_596),
        .a(_T_616),
        .b(_T_636)
    );
    wire [3:0] _T_638;
    CAT #(.width_a(1), .width_b(3)) cat_369 (
        .y(_T_638),
        .a(_T_596),
        .b(_T_637)
    );
    wire [3:0] _T_639;
    MUX_UNSIGNED #(.width(4)) u_mux_370 (
        .y(_T_639),
        .sel(_T_546),
        .a(_T_592),
        .b(_T_638)
    );
    wire [4:0] _T_640;
    CAT #(.width_a(1), .width_b(4)) cat_371 (
        .y(_T_640),
        .a(_T_546),
        .b(_T_639)
    );
    wire [15:0] _T_641;
    BITS #(.width(32), .high(31), .low(16)) bits_372 (
        .y(_T_641),
        .in(_T_540)
    );
    wire [15:0] _T_642;
    BITS #(.width(32), .high(15), .low(0)) bits_373 (
        .y(_T_642),
        .in(_T_540)
    );
    wire _T_644;
    wire [15:0] _WTEMP_46;
    PAD_UNSIGNED #(.width(1), .n(16)) u_pad_374 (
        .y(_WTEMP_46),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(16)) u_neq_375 (
        .y(_T_644),
        .a(_T_641),
        .b(_WTEMP_46)
    );
    wire [7:0] _T_645;
    BITS #(.width(16), .high(15), .low(8)) bits_376 (
        .y(_T_645),
        .in(_T_641)
    );
    wire [7:0] _T_646;
    BITS #(.width(16), .high(7), .low(0)) bits_377 (
        .y(_T_646),
        .in(_T_641)
    );
    wire _T_648;
    wire [7:0] _WTEMP_47;
    PAD_UNSIGNED #(.width(1), .n(8)) u_pad_378 (
        .y(_WTEMP_47),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(8)) u_neq_379 (
        .y(_T_648),
        .a(_T_645),
        .b(_WTEMP_47)
    );
    wire [3:0] _T_649;
    BITS #(.width(8), .high(7), .low(4)) bits_380 (
        .y(_T_649),
        .in(_T_645)
    );
    wire [3:0] _T_650;
    BITS #(.width(8), .high(3), .low(0)) bits_381 (
        .y(_T_650),
        .in(_T_645)
    );
    wire _T_652;
    wire [3:0] _WTEMP_48;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_382 (
        .y(_WTEMP_48),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_383 (
        .y(_T_652),
        .a(_T_649),
        .b(_WTEMP_48)
    );
    wire _T_653;
    BITS #(.width(4), .high(3), .low(3)) bits_384 (
        .y(_T_653),
        .in(_T_649)
    );
    wire _T_655;
    BITS #(.width(4), .high(2), .low(2)) bits_385 (
        .y(_T_655),
        .in(_T_649)
    );
    wire _T_657;
    BITS #(.width(4), .high(1), .low(1)) bits_386 (
        .y(_T_657),
        .in(_T_649)
    );
    wire [1:0] _T_658;
    wire [1:0] _WTEMP_49;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_387 (
        .y(_WTEMP_49),
        .in(_T_657)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_388 (
        .y(_T_658),
        .sel(_T_655),
        .a(2'h2),
        .b(_WTEMP_49)
    );
    wire [1:0] _T_659;
    MUX_UNSIGNED #(.width(2)) u_mux_389 (
        .y(_T_659),
        .sel(_T_653),
        .a(2'h3),
        .b(_T_658)
    );
    wire _T_660;
    BITS #(.width(4), .high(3), .low(3)) bits_390 (
        .y(_T_660),
        .in(_T_650)
    );
    wire _T_662;
    BITS #(.width(4), .high(2), .low(2)) bits_391 (
        .y(_T_662),
        .in(_T_650)
    );
    wire _T_664;
    BITS #(.width(4), .high(1), .low(1)) bits_392 (
        .y(_T_664),
        .in(_T_650)
    );
    wire [1:0] _T_665;
    wire [1:0] _WTEMP_50;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_393 (
        .y(_WTEMP_50),
        .in(_T_664)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_394 (
        .y(_T_665),
        .sel(_T_662),
        .a(2'h2),
        .b(_WTEMP_50)
    );
    wire [1:0] _T_666;
    MUX_UNSIGNED #(.width(2)) u_mux_395 (
        .y(_T_666),
        .sel(_T_660),
        .a(2'h3),
        .b(_T_665)
    );
    wire [1:0] _T_667;
    MUX_UNSIGNED #(.width(2)) u_mux_396 (
        .y(_T_667),
        .sel(_T_652),
        .a(_T_659),
        .b(_T_666)
    );
    wire [2:0] _T_668;
    CAT #(.width_a(1), .width_b(2)) cat_397 (
        .y(_T_668),
        .a(_T_652),
        .b(_T_667)
    );
    wire [3:0] _T_669;
    BITS #(.width(8), .high(7), .low(4)) bits_398 (
        .y(_T_669),
        .in(_T_646)
    );
    wire [3:0] _T_670;
    BITS #(.width(8), .high(3), .low(0)) bits_399 (
        .y(_T_670),
        .in(_T_646)
    );
    wire _T_672;
    wire [3:0] _WTEMP_51;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_400 (
        .y(_WTEMP_51),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_401 (
        .y(_T_672),
        .a(_T_669),
        .b(_WTEMP_51)
    );
    wire _T_673;
    BITS #(.width(4), .high(3), .low(3)) bits_402 (
        .y(_T_673),
        .in(_T_669)
    );
    wire _T_675;
    BITS #(.width(4), .high(2), .low(2)) bits_403 (
        .y(_T_675),
        .in(_T_669)
    );
    wire _T_677;
    BITS #(.width(4), .high(1), .low(1)) bits_404 (
        .y(_T_677),
        .in(_T_669)
    );
    wire [1:0] _T_678;
    wire [1:0] _WTEMP_52;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_405 (
        .y(_WTEMP_52),
        .in(_T_677)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_406 (
        .y(_T_678),
        .sel(_T_675),
        .a(2'h2),
        .b(_WTEMP_52)
    );
    wire [1:0] _T_679;
    MUX_UNSIGNED #(.width(2)) u_mux_407 (
        .y(_T_679),
        .sel(_T_673),
        .a(2'h3),
        .b(_T_678)
    );
    wire _T_680;
    BITS #(.width(4), .high(3), .low(3)) bits_408 (
        .y(_T_680),
        .in(_T_670)
    );
    wire _T_682;
    BITS #(.width(4), .high(2), .low(2)) bits_409 (
        .y(_T_682),
        .in(_T_670)
    );
    wire _T_684;
    BITS #(.width(4), .high(1), .low(1)) bits_410 (
        .y(_T_684),
        .in(_T_670)
    );
    wire [1:0] _T_685;
    wire [1:0] _WTEMP_53;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_411 (
        .y(_WTEMP_53),
        .in(_T_684)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_412 (
        .y(_T_685),
        .sel(_T_682),
        .a(2'h2),
        .b(_WTEMP_53)
    );
    wire [1:0] _T_686;
    MUX_UNSIGNED #(.width(2)) u_mux_413 (
        .y(_T_686),
        .sel(_T_680),
        .a(2'h3),
        .b(_T_685)
    );
    wire [1:0] _T_687;
    MUX_UNSIGNED #(.width(2)) u_mux_414 (
        .y(_T_687),
        .sel(_T_672),
        .a(_T_679),
        .b(_T_686)
    );
    wire [2:0] _T_688;
    CAT #(.width_a(1), .width_b(2)) cat_415 (
        .y(_T_688),
        .a(_T_672),
        .b(_T_687)
    );
    wire [2:0] _T_689;
    MUX_UNSIGNED #(.width(3)) u_mux_416 (
        .y(_T_689),
        .sel(_T_648),
        .a(_T_668),
        .b(_T_688)
    );
    wire [3:0] _T_690;
    CAT #(.width_a(1), .width_b(3)) cat_417 (
        .y(_T_690),
        .a(_T_648),
        .b(_T_689)
    );
    wire [7:0] _T_691;
    BITS #(.width(16), .high(15), .low(8)) bits_418 (
        .y(_T_691),
        .in(_T_642)
    );
    wire [7:0] _T_692;
    BITS #(.width(16), .high(7), .low(0)) bits_419 (
        .y(_T_692),
        .in(_T_642)
    );
    wire _T_694;
    wire [7:0] _WTEMP_54;
    PAD_UNSIGNED #(.width(1), .n(8)) u_pad_420 (
        .y(_WTEMP_54),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(8)) u_neq_421 (
        .y(_T_694),
        .a(_T_691),
        .b(_WTEMP_54)
    );
    wire [3:0] _T_695;
    BITS #(.width(8), .high(7), .low(4)) bits_422 (
        .y(_T_695),
        .in(_T_691)
    );
    wire [3:0] _T_696;
    BITS #(.width(8), .high(3), .low(0)) bits_423 (
        .y(_T_696),
        .in(_T_691)
    );
    wire _T_698;
    wire [3:0] _WTEMP_55;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_424 (
        .y(_WTEMP_55),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_425 (
        .y(_T_698),
        .a(_T_695),
        .b(_WTEMP_55)
    );
    wire _T_699;
    BITS #(.width(4), .high(3), .low(3)) bits_426 (
        .y(_T_699),
        .in(_T_695)
    );
    wire _T_701;
    BITS #(.width(4), .high(2), .low(2)) bits_427 (
        .y(_T_701),
        .in(_T_695)
    );
    wire _T_703;
    BITS #(.width(4), .high(1), .low(1)) bits_428 (
        .y(_T_703),
        .in(_T_695)
    );
    wire [1:0] _T_704;
    wire [1:0] _WTEMP_56;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_429 (
        .y(_WTEMP_56),
        .in(_T_703)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_430 (
        .y(_T_704),
        .sel(_T_701),
        .a(2'h2),
        .b(_WTEMP_56)
    );
    wire [1:0] _T_705;
    MUX_UNSIGNED #(.width(2)) u_mux_431 (
        .y(_T_705),
        .sel(_T_699),
        .a(2'h3),
        .b(_T_704)
    );
    wire _T_706;
    BITS #(.width(4), .high(3), .low(3)) bits_432 (
        .y(_T_706),
        .in(_T_696)
    );
    wire _T_708;
    BITS #(.width(4), .high(2), .low(2)) bits_433 (
        .y(_T_708),
        .in(_T_696)
    );
    wire _T_710;
    BITS #(.width(4), .high(1), .low(1)) bits_434 (
        .y(_T_710),
        .in(_T_696)
    );
    wire [1:0] _T_711;
    wire [1:0] _WTEMP_57;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_435 (
        .y(_WTEMP_57),
        .in(_T_710)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_436 (
        .y(_T_711),
        .sel(_T_708),
        .a(2'h2),
        .b(_WTEMP_57)
    );
    wire [1:0] _T_712;
    MUX_UNSIGNED #(.width(2)) u_mux_437 (
        .y(_T_712),
        .sel(_T_706),
        .a(2'h3),
        .b(_T_711)
    );
    wire [1:0] _T_713;
    MUX_UNSIGNED #(.width(2)) u_mux_438 (
        .y(_T_713),
        .sel(_T_698),
        .a(_T_705),
        .b(_T_712)
    );
    wire [2:0] _T_714;
    CAT #(.width_a(1), .width_b(2)) cat_439 (
        .y(_T_714),
        .a(_T_698),
        .b(_T_713)
    );
    wire [3:0] _T_715;
    BITS #(.width(8), .high(7), .low(4)) bits_440 (
        .y(_T_715),
        .in(_T_692)
    );
    wire [3:0] _T_716;
    BITS #(.width(8), .high(3), .low(0)) bits_441 (
        .y(_T_716),
        .in(_T_692)
    );
    wire _T_718;
    wire [3:0] _WTEMP_58;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_442 (
        .y(_WTEMP_58),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_443 (
        .y(_T_718),
        .a(_T_715),
        .b(_WTEMP_58)
    );
    wire _T_719;
    BITS #(.width(4), .high(3), .low(3)) bits_444 (
        .y(_T_719),
        .in(_T_715)
    );
    wire _T_721;
    BITS #(.width(4), .high(2), .low(2)) bits_445 (
        .y(_T_721),
        .in(_T_715)
    );
    wire _T_723;
    BITS #(.width(4), .high(1), .low(1)) bits_446 (
        .y(_T_723),
        .in(_T_715)
    );
    wire [1:0] _T_724;
    wire [1:0] _WTEMP_59;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_447 (
        .y(_WTEMP_59),
        .in(_T_723)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_448 (
        .y(_T_724),
        .sel(_T_721),
        .a(2'h2),
        .b(_WTEMP_59)
    );
    wire [1:0] _T_725;
    MUX_UNSIGNED #(.width(2)) u_mux_449 (
        .y(_T_725),
        .sel(_T_719),
        .a(2'h3),
        .b(_T_724)
    );
    wire _T_726;
    BITS #(.width(4), .high(3), .low(3)) bits_450 (
        .y(_T_726),
        .in(_T_716)
    );
    wire _T_728;
    BITS #(.width(4), .high(2), .low(2)) bits_451 (
        .y(_T_728),
        .in(_T_716)
    );
    wire _T_730;
    BITS #(.width(4), .high(1), .low(1)) bits_452 (
        .y(_T_730),
        .in(_T_716)
    );
    wire [1:0] _T_731;
    wire [1:0] _WTEMP_60;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_453 (
        .y(_WTEMP_60),
        .in(_T_730)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_454 (
        .y(_T_731),
        .sel(_T_728),
        .a(2'h2),
        .b(_WTEMP_60)
    );
    wire [1:0] _T_732;
    MUX_UNSIGNED #(.width(2)) u_mux_455 (
        .y(_T_732),
        .sel(_T_726),
        .a(2'h3),
        .b(_T_731)
    );
    wire [1:0] _T_733;
    MUX_UNSIGNED #(.width(2)) u_mux_456 (
        .y(_T_733),
        .sel(_T_718),
        .a(_T_725),
        .b(_T_732)
    );
    wire [2:0] _T_734;
    CAT #(.width_a(1), .width_b(2)) cat_457 (
        .y(_T_734),
        .a(_T_718),
        .b(_T_733)
    );
    wire [2:0] _T_735;
    MUX_UNSIGNED #(.width(3)) u_mux_458 (
        .y(_T_735),
        .sel(_T_694),
        .a(_T_714),
        .b(_T_734)
    );
    wire [3:0] _T_736;
    CAT #(.width_a(1), .width_b(3)) cat_459 (
        .y(_T_736),
        .a(_T_694),
        .b(_T_735)
    );
    wire [3:0] _T_737;
    MUX_UNSIGNED #(.width(4)) u_mux_460 (
        .y(_T_737),
        .sel(_T_644),
        .a(_T_690),
        .b(_T_736)
    );
    wire [4:0] _T_738;
    CAT #(.width_a(1), .width_b(4)) cat_461 (
        .y(_T_738),
        .a(_T_644),
        .b(_T_737)
    );
    wire [4:0] _T_739;
    MUX_UNSIGNED #(.width(5)) u_mux_462 (
        .y(_T_739),
        .sel(_T_542),
        .a(_T_640),
        .b(_T_738)
    );
    wire [5:0] _T_740;
    CAT #(.width_a(1), .width_b(5)) cat_463 (
        .y(_T_740),
        .a(_T_542),
        .b(_T_739)
    );
    wire [5:0] _T_741;
    BITWISENOT #(.width(6)) bitwisenot_464 (
        .y(_T_741),
        .in(_T_740)
    );
    wire [114:0] _T_742;
    DSHL_UNSIGNED #(.width_in(52), .width_n(6)) u_dshl_465 (
        .y(_T_742),
        .in(_T_532),
        .n(_T_741)
    );
    wire [50:0] _T_743;
    BITS #(.width(115), .high(50), .low(0)) bits_466 (
        .y(_T_743),
        .in(_T_742)
    );
    wire [51:0] _T_745;
    CAT #(.width_a(51), .width_b(1)) cat_467 (
        .y(_T_745),
        .a(_T_743),
        .b(1'h0)
    );
    wire [11:0] _T_750;
    assign _T_750 = 12'hFFF;
    wire [11:0] _T_751;
    wire [11:0] _WTEMP_61;
    PAD_UNSIGNED #(.width(6), .n(12)) u_pad_468 (
        .y(_WTEMP_61),
        .in(_T_741)
    );
    BITWISEXOR #(.width(12)) bitwisexor_469 (
        .y(_T_751),
        .a(_WTEMP_61),
        .b(_T_750)
    );
    wire [11:0] _T_752;
    wire [11:0] _WTEMP_62;
    PAD_UNSIGNED #(.width(11), .n(12)) u_pad_470 (
        .y(_WTEMP_62),
        .in(_T_531)
    );
    MUX_UNSIGNED #(.width(12)) u_mux_471 (
        .y(_T_752),
        .sel(_T_534),
        .a(_T_751),
        .b(_WTEMP_62)
    );
    wire [1:0] _T_756;
    wire [1:0] _WTEMP_63;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_472 (
        .y(_WTEMP_63),
        .in(1'h1)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_473 (
        .y(_T_756),
        .sel(_T_534),
        .a(2'h2),
        .b(_WTEMP_63)
    );
    wire [10:0] _T_757;
    wire [10:0] _WTEMP_64;
    PAD_UNSIGNED #(.width(2), .n(11)) u_pad_474 (
        .y(_WTEMP_64),
        .in(_T_756)
    );
    BITWISEOR #(.width(11)) bitwiseor_475 (
        .y(_T_757),
        .a(11'h400),
        .b(_WTEMP_64)
    );
    wire [12:0] _T_758;
    wire [11:0] _WTEMP_65;
    PAD_UNSIGNED #(.width(11), .n(12)) u_pad_476 (
        .y(_WTEMP_65),
        .in(_T_757)
    );
    ADD_UNSIGNED #(.width(12)) u_add_477 (
        .y(_T_758),
        .a(_T_752),
        .b(_WTEMP_65)
    );
    wire [11:0] _T_759;
    TAIL #(.width(13), .n(1)) tail_478 (
        .y(_T_759),
        .in(_T_758)
    );
    wire [1:0] _T_760;
    BITS #(.width(12), .high(11), .low(10)) bits_479 (
        .y(_T_760),
        .in(_T_759)
    );
    wire _T_762;
    EQ_UNSIGNED #(.width(2)) u_eq_480 (
        .y(_T_762),
        .a(_T_760),
        .b(2'h3)
    );
    wire _T_764;
    EQ_UNSIGNED #(.width(1)) u_eq_481 (
        .y(_T_764),
        .a(_T_536),
        .b(1'h0)
    );
    wire _T_765;
    BITWISEAND #(.width(1)) bitwiseand_482 (
        .y(_T_765),
        .a(_T_762),
        .b(_T_764)
    );
    wire _T_766;
    BITS #(.width(1), .high(0), .low(0)) bits_483 (
        .y(_T_766),
        .in(_T_537)
    );
    wire [2:0] _T_769;
    MUX_UNSIGNED #(.width(3)) u_mux_484 (
        .y(_T_769),
        .sel(_T_766),
        .a(3'h7),
        .b(3'h0)
    );
    wire [11:0] _T_770;
    SHL_UNSIGNED #(.width(3), .n(9)) u_shl_485 (
        .y(_T_770),
        .in(_T_769)
    );
    wire [11:0] _T_771;
    BITWISENOT #(.width(12)) bitwisenot_486 (
        .y(_T_771),
        .in(_T_770)
    );
    wire [11:0] _T_772;
    BITWISEAND #(.width(12)) bitwiseand_487 (
        .y(_T_772),
        .a(_T_759),
        .b(_T_771)
    );
    wire [9:0] _T_773;
    SHL_UNSIGNED #(.width(1), .n(9)) u_shl_488 (
        .y(_T_773),
        .in(_T_765)
    );
    wire [11:0] _T_774;
    wire [11:0] _WTEMP_66;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_489 (
        .y(_WTEMP_66),
        .in(_T_773)
    );
    BITWISEOR #(.width(12)) bitwiseor_490 (
        .y(_T_774),
        .a(_T_772),
        .b(_WTEMP_66)
    );
    wire [51:0] _T_775;
    MUX_UNSIGNED #(.width(52)) u_mux_491 (
        .y(_T_775),
        .sel(_T_534),
        .a(_T_745),
        .b(_T_532)
    );
    wire [12:0] _T_776;
    CAT #(.width_a(1), .width_b(12)) cat_492 (
        .y(_T_776),
        .a(_T_530),
        .b(_T_774)
    );
    wire [64:0] _T_777;
    CAT #(.width_a(13), .width_b(52)) cat_493 (
        .y(_T_777),
        .a(_T_776),
        .b(_T_775)
    );
    wire [64:0] _T_779;
    wire [64:0] _WTEMP_67;
    PAD_UNSIGNED #(.width(33), .n(65)) u_pad_494 (
        .y(_WTEMP_67),
        .in(rec_s)
    );
    BITWISEOR #(.width(65)) bitwiseor_495 (
        .y(_T_779),
        .a(_WTEMP_67),
        .b(65'hE004000000000000)
    );
    wire [64:0] load_wb_data_recoded;
    MUX_UNSIGNED #(.width(65)) u_mux_496 (
        .y(load_wb_data_recoded),
        .sel(_load_wb_single__q),
        .a(_T_779),
        .b(_T_777)
    );
    wire regfile__T_782_clk;
    wire regfile__T_782_en;
    wire regfile__T_782_mask;
    wire [4:0] regfile__T_782_addr;
    wire [64:0] regfile__T_782_data;
    wire [64:0] regfile__T_849_data;
    wire regfile__T_849_clk;
    wire regfile__T_849_en;
    wire [4:0] regfile__T_849_addr;
    wire [64:0] regfile__T_853_data;
    wire regfile__T_853_clk;
    wire regfile__T_853_en;
    wire [4:0] regfile__T_853_addr;
    wire [64:0] regfile__T_857_data;
    wire regfile__T_857_clk;
    wire regfile__T_857_en;
    wire [4:0] regfile__T_857_addr;
    wire regfile__T_1131_clk;
    wire regfile__T_1131_en;
    wire regfile__T_1131_mask;
    wire [4:0] regfile__T_1131_addr;
    wire [64:0] regfile__T_1131_data;
    wire [194:0] regfile_read_datas;
    wire [2:0] regfile_read_clks;
    wire [2:0] regfile_read_ens;
    wire [14:0] regfile_read_addrs;
    wire [1:0] regfile_write_clks;
    wire [1:0] regfile_write_ens;
    wire [1:0] regfile_write_masks;
    wire [9:0] regfile_write_addrs;
    wire [129:0] regfile_write_datas;
    BITS #(.width(195), .high(64), .low(0)) bits_497 (
        .y(regfile__T_849_data),
        .in(regfile_read_datas)
    );
    BITS #(.width(195), .high(129), .low(65)) bits_498 (
        .y(regfile__T_853_data),
        .in(regfile_read_datas)
    );
    BITS #(.width(195), .high(194), .low(130)) bits_499 (
        .y(regfile__T_857_data),
        .in(regfile_read_datas)
    );
    wire [1:0] _WTEMP_68;
    CAT #(.width_a(1), .width_b(1)) cat_500 (
        .y(_WTEMP_68),
        .a(regfile__T_857_clk),
        .b(regfile__T_853_clk)
    );
    CAT #(.width_a(2), .width_b(1)) cat_501 (
        .y(regfile_read_clks),
        .a(_WTEMP_68),
        .b(regfile__T_849_clk)
    );
    wire [1:0] _WTEMP_69;
    CAT #(.width_a(1), .width_b(1)) cat_502 (
        .y(_WTEMP_69),
        .a(regfile__T_857_en),
        .b(regfile__T_853_en)
    );
    CAT #(.width_a(2), .width_b(1)) cat_503 (
        .y(regfile_read_ens),
        .a(_WTEMP_69),
        .b(regfile__T_849_en)
    );
    wire [9:0] _WTEMP_70;
    CAT #(.width_a(5), .width_b(5)) cat_504 (
        .y(_WTEMP_70),
        .a(regfile__T_857_addr),
        .b(regfile__T_853_addr)
    );
    CAT #(.width_a(10), .width_b(5)) cat_505 (
        .y(regfile_read_addrs),
        .a(_WTEMP_70),
        .b(regfile__T_849_addr)
    );
    CAT #(.width_a(65), .width_b(65)) cat_506 (
        .y(regfile_write_datas),
        .a(regfile__T_1131_data),
        .b(regfile__T_782_data)
    );
    CAT #(.width_a(1), .width_b(1)) cat_507 (
        .y(regfile_write_clks),
        .a(regfile__T_1131_clk),
        .b(regfile__T_782_clk)
    );
    CAT #(.width_a(1), .width_b(1)) cat_508 (
        .y(regfile_write_ens),
        .a(regfile__T_1131_en),
        .b(regfile__T_782_en)
    );
    CAT #(.width_a(5), .width_b(5)) cat_509 (
        .y(regfile_write_addrs),
        .a(regfile__T_1131_addr),
        .b(regfile__T_782_addr)
    );
    CAT #(.width_a(1), .width_b(1)) cat_510 (
        .y(regfile_write_masks),
        .a(regfile__T_1131_mask),
        .b(regfile__T_782_mask)
    );
    MRMWMEM #(.depth(32), .addrbits(5), .width(65), .readernum(3), .writernum(2), .isSyncRead(0)) regfile (
        .read_datas(regfile_read_datas),
        .read_clks(regfile_read_clks),
        .read_ens(regfile_read_ens),
        .read_addrs(regfile_read_addrs),
        .write_clks(regfile_write_clks),
        .write_ens(regfile_write_ens),
        .write_masks(regfile_write_masks),
        .write_addrs(regfile_write_addrs),
        .write_datas(regfile_write_datas)
    );
    assign regfile__T_782_addr = _load_wb_tag__q;
    assign regfile__T_782_en = _load_wb__q;
    assign regfile__T_782_clk = clock;
    assign regfile__T_782_mask = 1'h1;
    wire [4:0] _ex_ra1__q;
    wire [4:0] _ex_ra1__d;
    DFF_POSCLK #(.width(5)) ex_ra1 (
        .q(_ex_ra1__q),
        .d(_ex_ra1__d),
        .clk(clock)
    );
    wire [4:0] _ex_ra2__q;
    wire [4:0] _ex_ra2__d;
    DFF_POSCLK #(.width(5)) ex_ra2 (
        .q(_ex_ra2__q),
        .d(_ex_ra2__d),
        .clk(clock)
    );
    wire [4:0] _ex_ra3__q;
    wire [4:0] _ex_ra3__d;
    DFF_POSCLK #(.width(5)) ex_ra3 (
        .q(_ex_ra3__q),
        .d(_ex_ra3__d),
        .clk(clock)
    );
    wire _T_787;
    EQ_UNSIGNED #(.width(1)) u_eq_511 (
        .y(_T_787),
        .a(_fp_decoder__io_sigs_swap12),
        .b(1'h0)
    );
    wire [4:0] _T_788;
    BITS #(.width(32), .high(19), .low(15)) bits_512 (
        .y(_T_788),
        .in(io_inst)
    );
    wire [4:0] _T_789;
    BITS #(.width(32), .high(19), .low(15)) bits_513 (
        .y(_T_789),
        .in(io_inst)
    );
    wire [4:0] _node_0;
    MUX_UNSIGNED #(.width(5)) u_mux_514 (
        .y(_node_0),
        .sel(_T_787),
        .a(_T_788),
        .b(_ex_ra1__q)
    );
    wire [4:0] _node_1;
    MUX_UNSIGNED #(.width(5)) u_mux_515 (
        .y(_node_1),
        .sel(_fp_decoder__io_sigs_swap12),
        .a(_T_789),
        .b(_ex_ra2__q)
    );
    wire [4:0] _T_790;
    BITS #(.width(32), .high(24), .low(20)) bits_516 (
        .y(_T_790),
        .in(io_inst)
    );
    wire [4:0] _node_2;
    MUX_UNSIGNED #(.width(5)) u_mux_517 (
        .y(_node_2),
        .sel(_fp_decoder__io_sigs_ren1),
        .a(_node_0),
        .b(_ex_ra1__q)
    );
    wire [4:0] _T_791;
    BITS #(.width(32), .high(24), .low(20)) bits_518 (
        .y(_T_791),
        .in(io_inst)
    );
    wire _T_793;
    EQ_UNSIGNED #(.width(1)) u_eq_519 (
        .y(_T_793),
        .a(_fp_decoder__io_sigs_swap12),
        .b(1'h0)
    );
    wire _T_795;
    EQ_UNSIGNED #(.width(1)) u_eq_520 (
        .y(_T_795),
        .a(_fp_decoder__io_sigs_swap23),
        .b(1'h0)
    );
    wire _T_796;
    BITWISEAND #(.width(1)) bitwiseand_521 (
        .y(_T_796),
        .a(_T_793),
        .b(_T_795)
    );
    wire [4:0] _T_797;
    BITS #(.width(32), .high(24), .low(20)) bits_522 (
        .y(_T_797),
        .in(io_inst)
    );
    wire [4:0] _node_3;
    MUX_UNSIGNED #(.width(5)) u_mux_523 (
        .y(_node_3),
        .sel(_fp_decoder__io_sigs_ren1),
        .a(_node_1),
        .b(_ex_ra2__q)
    );
    wire [4:0] _node_4;
    MUX_UNSIGNED #(.width(5)) u_mux_524 (
        .y(_node_4),
        .sel(_fp_decoder__io_sigs_swap12),
        .a(_T_790),
        .b(_node_2)
    );
    wire [4:0] _node_5;
    MUX_UNSIGNED #(.width(5)) u_mux_525 (
        .y(_node_5),
        .sel(_fp_decoder__io_sigs_ren1),
        .a(_node_0),
        .b(_ex_ra1__q)
    );
    wire [4:0] _node_6;
    MUX_UNSIGNED #(.width(5)) u_mux_526 (
        .y(_node_6),
        .sel(_T_796),
        .a(_T_797),
        .b(_node_3)
    );
    wire [4:0] _node_7;
    MUX_UNSIGNED #(.width(5)) u_mux_527 (
        .y(_node_7),
        .sel(_fp_decoder__io_sigs_ren1),
        .a(_node_1),
        .b(_ex_ra2__q)
    );
    wire [4:0] _node_8;
    MUX_UNSIGNED #(.width(5)) u_mux_528 (
        .y(_node_8),
        .sel(_fp_decoder__io_sigs_swap23),
        .a(_T_791),
        .b(_ex_ra3__q)
    );
    wire [4:0] _T_798;
    BITS #(.width(32), .high(31), .low(27)) bits_529 (
        .y(_T_798),
        .in(io_inst)
    );
    wire [4:0] _node_9;
    MUX_UNSIGNED #(.width(5)) u_mux_530 (
        .y(_node_9),
        .sel(_fp_decoder__io_sigs_ren2),
        .a(_node_8),
        .b(_ex_ra3__q)
    );
    wire [4:0] _node_10;
    MUX_UNSIGNED #(.width(5)) u_mux_531 (
        .y(_node_10),
        .sel(_fp_decoder__io_sigs_ren2),
        .a(_node_4),
        .b(_node_5)
    );
    wire [4:0] _node_11;
    MUX_UNSIGNED #(.width(5)) u_mux_532 (
        .y(_node_11),
        .sel(_fp_decoder__io_sigs_ren2),
        .a(_node_6),
        .b(_node_7)
    );
    wire [4:0] _node_12;
    MUX_UNSIGNED #(.width(5)) u_mux_533 (
        .y(_node_12),
        .sel(_fp_decoder__io_sigs_ren3),
        .a(_T_798),
        .b(_node_9)
    );
    wire [2:0] _T_799;
    BITS #(.width(32), .high(14), .low(12)) bits_534 (
        .y(_T_799),
        .in(_ex_reg_inst__q)
    );
    wire _T_801;
    EQ_UNSIGNED #(.width(3)) u_eq_535 (
        .y(_T_801),
        .a(_T_799),
        .b(3'h7)
    );
    wire [2:0] _T_802;
    BITS #(.width(32), .high(14), .low(12)) bits_536 (
        .y(_T_802),
        .in(_ex_reg_inst__q)
    );
    wire [2:0] ex_rm;
    MUX_UNSIGNED #(.width(3)) u_mux_537 (
        .y(ex_rm),
        .sel(_T_801),
        .a(io_fcsr_rm),
        .b(_T_802)
    );
    wire [4:0] req_cmd;
    wire req_ldst;
    wire req_wen;
    wire req_ren1;
    wire req_ren2;
    wire req_ren3;
    wire req_swap12;
    wire req_swap23;
    wire req_single;
    wire req_fromint;
    wire req_toint;
    wire req_fastpipe;
    wire req_fma;
    wire req_div;
    wire req_sqrt;
    wire req_wflags;
    wire [2:0] req_rm;
    wire [1:0] req_typ;
    wire [64:0] req_in1;
    wire [64:0] req_in2;
    wire [64:0] req_in3;
    wire [4:0] _T_847;
    BITWISEOR #(.width(5)) bitwiseor_538 (
        .y(_T_847),
        .a(_ex_ra1__q),
        .b(5'h0)
    );
    wire [4:0] _T_848;
    BITS #(.width(5), .high(4), .low(0)) bits_539 (
        .y(_T_848),
        .in(_T_847)
    );
    assign regfile__T_849_addr = _T_848;
    assign regfile__T_849_en = 1'h1;
    assign regfile__T_849_clk = clock;
    wire [4:0] _T_851;
    BITWISEOR #(.width(5)) bitwiseor_540 (
        .y(_T_851),
        .a(_ex_ra2__q),
        .b(5'h0)
    );
    wire [4:0] _T_852;
    BITS #(.width(5), .high(4), .low(0)) bits_541 (
        .y(_T_852),
        .in(_T_851)
    );
    assign regfile__T_853_addr = _T_852;
    assign regfile__T_853_en = 1'h1;
    assign regfile__T_853_clk = clock;
    wire [4:0] _T_855;
    BITWISEOR #(.width(5)) bitwiseor_542 (
        .y(_T_855),
        .a(_ex_ra3__q),
        .b(5'h0)
    );
    wire [4:0] _T_856;
    BITS #(.width(5), .high(4), .low(0)) bits_543 (
        .y(_T_856),
        .in(_T_855)
    );
    assign regfile__T_857_addr = _T_856;
    assign regfile__T_857_en = 1'h1;
    assign regfile__T_857_clk = clock;
    wire [1:0] _T_858;
    BITS #(.width(32), .high(21), .low(20)) bits_544 (
        .y(_T_858),
        .in(_ex_reg_inst__q)
    );
    wire [64:0] _node_13;
    MUX_UNSIGNED #(.width(65)) u_mux_545 (
        .y(_node_13),
        .sel(io_cp_req_bits_swap23),
        .a(io_cp_req_bits_in3),
        .b(io_cp_req_bits_in2)
    );
    wire [64:0] _node_14;
    MUX_UNSIGNED #(.width(65)) u_mux_546 (
        .y(_node_14),
        .sel(io_cp_req_bits_swap23),
        .a(io_cp_req_bits_in2),
        .b(io_cp_req_bits_in3)
    );
    wire _sfma__clock;
    wire _sfma__reset;
    wire _sfma__io_in_valid;
    wire [4:0] _sfma__io_in_bits_cmd;
    wire _sfma__io_in_bits_ldst;
    wire _sfma__io_in_bits_wen;
    wire _sfma__io_in_bits_ren1;
    wire _sfma__io_in_bits_ren2;
    wire _sfma__io_in_bits_ren3;
    wire _sfma__io_in_bits_swap12;
    wire _sfma__io_in_bits_swap23;
    wire _sfma__io_in_bits_single;
    wire _sfma__io_in_bits_fromint;
    wire _sfma__io_in_bits_toint;
    wire _sfma__io_in_bits_fastpipe;
    wire _sfma__io_in_bits_fma;
    wire _sfma__io_in_bits_div;
    wire _sfma__io_in_bits_sqrt;
    wire _sfma__io_in_bits_wflags;
    wire [2:0] _sfma__io_in_bits_rm;
    wire [1:0] _sfma__io_in_bits_typ;
    wire [64:0] _sfma__io_in_bits_in1;
    wire [64:0] _sfma__io_in_bits_in2;
    wire [64:0] _sfma__io_in_bits_in3;
    wire _sfma__io_out_valid;
    wire [64:0] _sfma__io_out_bits_data;
    wire [4:0] _sfma__io_out_bits_exc;
    FPUFMAPipe sfma (
        .clock(_sfma__clock),
        .reset(_sfma__reset),
        .io_in_valid(_sfma__io_in_valid),
        .io_in_bits_cmd(_sfma__io_in_bits_cmd),
        .io_in_bits_ldst(_sfma__io_in_bits_ldst),
        .io_in_bits_wen(_sfma__io_in_bits_wen),
        .io_in_bits_ren1(_sfma__io_in_bits_ren1),
        .io_in_bits_ren2(_sfma__io_in_bits_ren2),
        .io_in_bits_ren3(_sfma__io_in_bits_ren3),
        .io_in_bits_swap12(_sfma__io_in_bits_swap12),
        .io_in_bits_swap23(_sfma__io_in_bits_swap23),
        .io_in_bits_single(_sfma__io_in_bits_single),
        .io_in_bits_fromint(_sfma__io_in_bits_fromint),
        .io_in_bits_toint(_sfma__io_in_bits_toint),
        .io_in_bits_fastpipe(_sfma__io_in_bits_fastpipe),
        .io_in_bits_fma(_sfma__io_in_bits_fma),
        .io_in_bits_div(_sfma__io_in_bits_div),
        .io_in_bits_sqrt(_sfma__io_in_bits_sqrt),
        .io_in_bits_wflags(_sfma__io_in_bits_wflags),
        .io_in_bits_rm(_sfma__io_in_bits_rm),
        .io_in_bits_typ(_sfma__io_in_bits_typ),
        .io_in_bits_in1(_sfma__io_in_bits_in1),
        .io_in_bits_in2(_sfma__io_in_bits_in2),
        .io_in_bits_in3(_sfma__io_in_bits_in3),
        .io_out_valid(_sfma__io_out_valid),
        .io_out_bits_data(_sfma__io_out_bits_data),
        .io_out_bits_exc(_sfma__io_out_bits_exc)
    );
    wire _T_859;
    BITWISEAND #(.width(1)) bitwiseand_1455 (
        .y(_T_859),
        .a(req_valid),
        .b(ex_ctrl_fma)
    );
    wire _T_860;
    BITWISEAND #(.width(1)) bitwiseand_1456 (
        .y(_T_860),
        .a(_T_859),
        .b(ex_ctrl_single)
    );
    wire _fpiu__clock;
    wire _fpiu__reset;
    wire _fpiu__io_in_valid;
    wire [4:0] _fpiu__io_in_bits_cmd;
    wire _fpiu__io_in_bits_ldst;
    wire _fpiu__io_in_bits_wen;
    wire _fpiu__io_in_bits_ren1;
    wire _fpiu__io_in_bits_ren2;
    wire _fpiu__io_in_bits_ren3;
    wire _fpiu__io_in_bits_swap12;
    wire _fpiu__io_in_bits_swap23;
    wire _fpiu__io_in_bits_single;
    wire _fpiu__io_in_bits_fromint;
    wire _fpiu__io_in_bits_toint;
    wire _fpiu__io_in_bits_fastpipe;
    wire _fpiu__io_in_bits_fma;
    wire _fpiu__io_in_bits_div;
    wire _fpiu__io_in_bits_sqrt;
    wire _fpiu__io_in_bits_wflags;
    wire [2:0] _fpiu__io_in_bits_rm;
    wire [1:0] _fpiu__io_in_bits_typ;
    wire [64:0] _fpiu__io_in_bits_in1;
    wire [64:0] _fpiu__io_in_bits_in2;
    wire [64:0] _fpiu__io_in_bits_in3;
    wire [4:0] _fpiu__io_as_double_cmd;
    wire _fpiu__io_as_double_ldst;
    wire _fpiu__io_as_double_wen;
    wire _fpiu__io_as_double_ren1;
    wire _fpiu__io_as_double_ren2;
    wire _fpiu__io_as_double_ren3;
    wire _fpiu__io_as_double_swap12;
    wire _fpiu__io_as_double_swap23;
    wire _fpiu__io_as_double_single;
    wire _fpiu__io_as_double_fromint;
    wire _fpiu__io_as_double_toint;
    wire _fpiu__io_as_double_fastpipe;
    wire _fpiu__io_as_double_fma;
    wire _fpiu__io_as_double_div;
    wire _fpiu__io_as_double_sqrt;
    wire _fpiu__io_as_double_wflags;
    wire [2:0] _fpiu__io_as_double_rm;
    wire [1:0] _fpiu__io_as_double_typ;
    wire [64:0] _fpiu__io_as_double_in1;
    wire [64:0] _fpiu__io_as_double_in2;
    wire [64:0] _fpiu__io_as_double_in3;
    wire _fpiu__io_out_valid;
    wire _fpiu__io_out_bits_lt;
    wire [63:0] _fpiu__io_out_bits_store;
    wire [63:0] _fpiu__io_out_bits_toint;
    wire [4:0] _fpiu__io_out_bits_exc;
    FPToInt fpiu (
        .clock(_fpiu__clock),
        .reset(_fpiu__reset),
        .io_in_valid(_fpiu__io_in_valid),
        .io_in_bits_cmd(_fpiu__io_in_bits_cmd),
        .io_in_bits_ldst(_fpiu__io_in_bits_ldst),
        .io_in_bits_wen(_fpiu__io_in_bits_wen),
        .io_in_bits_ren1(_fpiu__io_in_bits_ren1),
        .io_in_bits_ren2(_fpiu__io_in_bits_ren2),
        .io_in_bits_ren3(_fpiu__io_in_bits_ren3),
        .io_in_bits_swap12(_fpiu__io_in_bits_swap12),
        .io_in_bits_swap23(_fpiu__io_in_bits_swap23),
        .io_in_bits_single(_fpiu__io_in_bits_single),
        .io_in_bits_fromint(_fpiu__io_in_bits_fromint),
        .io_in_bits_toint(_fpiu__io_in_bits_toint),
        .io_in_bits_fastpipe(_fpiu__io_in_bits_fastpipe),
        .io_in_bits_fma(_fpiu__io_in_bits_fma),
        .io_in_bits_div(_fpiu__io_in_bits_div),
        .io_in_bits_sqrt(_fpiu__io_in_bits_sqrt),
        .io_in_bits_wflags(_fpiu__io_in_bits_wflags),
        .io_in_bits_rm(_fpiu__io_in_bits_rm),
        .io_in_bits_typ(_fpiu__io_in_bits_typ),
        .io_in_bits_in1(_fpiu__io_in_bits_in1),
        .io_in_bits_in2(_fpiu__io_in_bits_in2),
        .io_in_bits_in3(_fpiu__io_in_bits_in3),
        .io_as_double_cmd(_fpiu__io_as_double_cmd),
        .io_as_double_ldst(_fpiu__io_as_double_ldst),
        .io_as_double_wen(_fpiu__io_as_double_wen),
        .io_as_double_ren1(_fpiu__io_as_double_ren1),
        .io_as_double_ren2(_fpiu__io_as_double_ren2),
        .io_as_double_ren3(_fpiu__io_as_double_ren3),
        .io_as_double_swap12(_fpiu__io_as_double_swap12),
        .io_as_double_swap23(_fpiu__io_as_double_swap23),
        .io_as_double_single(_fpiu__io_as_double_single),
        .io_as_double_fromint(_fpiu__io_as_double_fromint),
        .io_as_double_toint(_fpiu__io_as_double_toint),
        .io_as_double_fastpipe(_fpiu__io_as_double_fastpipe),
        .io_as_double_fma(_fpiu__io_as_double_fma),
        .io_as_double_div(_fpiu__io_as_double_div),
        .io_as_double_sqrt(_fpiu__io_as_double_sqrt),
        .io_as_double_wflags(_fpiu__io_as_double_wflags),
        .io_as_double_rm(_fpiu__io_as_double_rm),
        .io_as_double_typ(_fpiu__io_as_double_typ),
        .io_as_double_in1(_fpiu__io_as_double_in1),
        .io_as_double_in2(_fpiu__io_as_double_in2),
        .io_as_double_in3(_fpiu__io_as_double_in3),
        .io_out_valid(_fpiu__io_out_valid),
        .io_out_bits_lt(_fpiu__io_out_bits_lt),
        .io_out_bits_store(_fpiu__io_out_bits_store),
        .io_out_bits_toint(_fpiu__io_out_bits_toint),
        .io_out_bits_exc(_fpiu__io_out_bits_exc)
    );
    wire _T_861;
    BITWISEOR #(.width(1)) bitwiseor_2136 (
        .y(_T_861),
        .a(ex_ctrl_toint),
        .b(ex_ctrl_div)
    );
    wire _T_862;
    BITWISEOR #(.width(1)) bitwiseor_2137 (
        .y(_T_862),
        .a(_T_861),
        .b(ex_ctrl_sqrt)
    );
    wire [4:0] _T_865;
    wire [4:0] _WTEMP_274;
    PAD_UNSIGNED #(.width(4), .n(5)) u_pad_2138 (
        .y(_WTEMP_274),
        .in(4'hD)
    );
    BITWISEAND #(.width(5)) bitwiseand_2139 (
        .y(_T_865),
        .a(ex_ctrl_cmd),
        .b(_WTEMP_274)
    );
    wire _T_866;
    wire [4:0] _WTEMP_275;
    PAD_UNSIGNED #(.width(3), .n(5)) u_pad_2140 (
        .y(_WTEMP_275),
        .in(3'h5)
    );
    EQ_UNSIGNED #(.width(5)) u_eq_2141 (
        .y(_T_866),
        .a(_WTEMP_275),
        .b(_T_865)
    );
    wire _T_867;
    BITWISEOR #(.width(1)) bitwiseor_2142 (
        .y(_T_867),
        .a(_T_862),
        .b(_T_866)
    );
    wire _T_868;
    BITWISEAND #(.width(1)) bitwiseand_2143 (
        .y(_T_868),
        .a(req_valid),
        .b(_T_867)
    );
    wire _T_869;
    BITWISEAND #(.width(1)) bitwiseand_2144 (
        .y(_T_869),
        .a(_fpiu__io_out_valid),
        .b(_mem_cp_valid__q)
    );
    wire _T_870;
    BITWISEAND #(.width(1)) bitwiseand_2145 (
        .y(_T_870),
        .a(_T_869),
        .b(_mem_ctrl_toint__q)
    );
    wire _ifpu__clock;
    wire _ifpu__reset;
    wire _ifpu__io_in_valid;
    wire [4:0] _ifpu__io_in_bits_cmd;
    wire _ifpu__io_in_bits_ldst;
    wire _ifpu__io_in_bits_wen;
    wire _ifpu__io_in_bits_ren1;
    wire _ifpu__io_in_bits_ren2;
    wire _ifpu__io_in_bits_ren3;
    wire _ifpu__io_in_bits_swap12;
    wire _ifpu__io_in_bits_swap23;
    wire _ifpu__io_in_bits_single;
    wire _ifpu__io_in_bits_fromint;
    wire _ifpu__io_in_bits_toint;
    wire _ifpu__io_in_bits_fastpipe;
    wire _ifpu__io_in_bits_fma;
    wire _ifpu__io_in_bits_div;
    wire _ifpu__io_in_bits_sqrt;
    wire _ifpu__io_in_bits_wflags;
    wire [2:0] _ifpu__io_in_bits_rm;
    wire [1:0] _ifpu__io_in_bits_typ;
    wire [64:0] _ifpu__io_in_bits_in1;
    wire [64:0] _ifpu__io_in_bits_in2;
    wire [64:0] _ifpu__io_in_bits_in3;
    wire _ifpu__io_out_valid;
    wire [64:0] _ifpu__io_out_bits_data;
    wire [4:0] _ifpu__io_out_bits_exc;
    IntToFP ifpu (
        .clock(_ifpu__clock),
        .reset(_ifpu__reset),
        .io_in_valid(_ifpu__io_in_valid),
        .io_in_bits_cmd(_ifpu__io_in_bits_cmd),
        .io_in_bits_ldst(_ifpu__io_in_bits_ldst),
        .io_in_bits_wen(_ifpu__io_in_bits_wen),
        .io_in_bits_ren1(_ifpu__io_in_bits_ren1),
        .io_in_bits_ren2(_ifpu__io_in_bits_ren2),
        .io_in_bits_ren3(_ifpu__io_in_bits_ren3),
        .io_in_bits_swap12(_ifpu__io_in_bits_swap12),
        .io_in_bits_swap23(_ifpu__io_in_bits_swap23),
        .io_in_bits_single(_ifpu__io_in_bits_single),
        .io_in_bits_fromint(_ifpu__io_in_bits_fromint),
        .io_in_bits_toint(_ifpu__io_in_bits_toint),
        .io_in_bits_fastpipe(_ifpu__io_in_bits_fastpipe),
        .io_in_bits_fma(_ifpu__io_in_bits_fma),
        .io_in_bits_div(_ifpu__io_in_bits_div),
        .io_in_bits_sqrt(_ifpu__io_in_bits_sqrt),
        .io_in_bits_wflags(_ifpu__io_in_bits_wflags),
        .io_in_bits_rm(_ifpu__io_in_bits_rm),
        .io_in_bits_typ(_ifpu__io_in_bits_typ),
        .io_in_bits_in1(_ifpu__io_in_bits_in1),
        .io_in_bits_in2(_ifpu__io_in_bits_in2),
        .io_in_bits_in3(_ifpu__io_in_bits_in3),
        .io_out_valid(_ifpu__io_out_valid),
        .io_out_bits_data(_ifpu__io_out_bits_data),
        .io_out_bits_exc(_ifpu__io_out_bits_exc)
    );
    wire _T_872;
    BITWISEAND #(.width(1)) bitwiseand_3054 (
        .y(_T_872),
        .a(req_valid),
        .b(ex_ctrl_fromint)
    );
    wire [64:0] _T_873;
    wire [64:0] _WTEMP_422;
    PAD_UNSIGNED #(.width(64), .n(65)) u_pad_3055 (
        .y(_WTEMP_422),
        .in(io_fromint_data)
    );
    MUX_UNSIGNED #(.width(65)) u_mux_3056 (
        .y(_T_873),
        .sel(ex_cp_valid),
        .a(io_cp_req_bits_in1),
        .b(_WTEMP_422)
    );
    wire _fpmu__clock;
    wire _fpmu__reset;
    wire _fpmu__io_in_valid;
    wire [4:0] _fpmu__io_in_bits_cmd;
    wire _fpmu__io_in_bits_ldst;
    wire _fpmu__io_in_bits_wen;
    wire _fpmu__io_in_bits_ren1;
    wire _fpmu__io_in_bits_ren2;
    wire _fpmu__io_in_bits_ren3;
    wire _fpmu__io_in_bits_swap12;
    wire _fpmu__io_in_bits_swap23;
    wire _fpmu__io_in_bits_single;
    wire _fpmu__io_in_bits_fromint;
    wire _fpmu__io_in_bits_toint;
    wire _fpmu__io_in_bits_fastpipe;
    wire _fpmu__io_in_bits_fma;
    wire _fpmu__io_in_bits_div;
    wire _fpmu__io_in_bits_sqrt;
    wire _fpmu__io_in_bits_wflags;
    wire [2:0] _fpmu__io_in_bits_rm;
    wire [1:0] _fpmu__io_in_bits_typ;
    wire [64:0] _fpmu__io_in_bits_in1;
    wire [64:0] _fpmu__io_in_bits_in2;
    wire [64:0] _fpmu__io_in_bits_in3;
    wire _fpmu__io_out_valid;
    wire [64:0] _fpmu__io_out_bits_data;
    wire [4:0] _fpmu__io_out_bits_exc;
    wire _fpmu__io_lt;
    FPToFP fpmu (
        .clock(_fpmu__clock),
        .reset(_fpmu__reset),
        .io_in_valid(_fpmu__io_in_valid),
        .io_in_bits_cmd(_fpmu__io_in_bits_cmd),
        .io_in_bits_ldst(_fpmu__io_in_bits_ldst),
        .io_in_bits_wen(_fpmu__io_in_bits_wen),
        .io_in_bits_ren1(_fpmu__io_in_bits_ren1),
        .io_in_bits_ren2(_fpmu__io_in_bits_ren2),
        .io_in_bits_ren3(_fpmu__io_in_bits_ren3),
        .io_in_bits_swap12(_fpmu__io_in_bits_swap12),
        .io_in_bits_swap23(_fpmu__io_in_bits_swap23),
        .io_in_bits_single(_fpmu__io_in_bits_single),
        .io_in_bits_fromint(_fpmu__io_in_bits_fromint),
        .io_in_bits_toint(_fpmu__io_in_bits_toint),
        .io_in_bits_fastpipe(_fpmu__io_in_bits_fastpipe),
        .io_in_bits_fma(_fpmu__io_in_bits_fma),
        .io_in_bits_div(_fpmu__io_in_bits_div),
        .io_in_bits_sqrt(_fpmu__io_in_bits_sqrt),
        .io_in_bits_wflags(_fpmu__io_in_bits_wflags),
        .io_in_bits_rm(_fpmu__io_in_bits_rm),
        .io_in_bits_typ(_fpmu__io_in_bits_typ),
        .io_in_bits_in1(_fpmu__io_in_bits_in1),
        .io_in_bits_in2(_fpmu__io_in_bits_in2),
        .io_in_bits_in3(_fpmu__io_in_bits_in3),
        .io_out_valid(_fpmu__io_out_valid),
        .io_out_bits_data(_fpmu__io_out_bits_data),
        .io_out_bits_exc(_fpmu__io_out_bits_exc),
        .io_lt(_fpmu__io_lt)
    );
    wire _T_874;
    BITWISEAND #(.width(1)) bitwiseand_3477 (
        .y(_T_874),
        .a(req_valid),
        .b(ex_ctrl_fastpipe)
    );
    wire _divSqrt_wen__q;
    wire _divSqrt_wen__d;
    DFF_POSCLK #(.width(1)) divSqrt_wen (
        .q(_divSqrt_wen__q),
        .d(_divSqrt_wen__d),
        .clk(clock)
    );
    wire divSqrt_inReady;
    wire [4:0] _divSqrt_waddr__q;
    wire [4:0] _divSqrt_waddr__d;
    DFF_POSCLK #(.width(5)) divSqrt_waddr (
        .q(_divSqrt_waddr__q),
        .d(_divSqrt_waddr__d),
        .clk(clock)
    );
    wire _divSqrt_single__q;
    wire _divSqrt_single__d;
    DFF_POSCLK #(.width(1)) divSqrt_single (
        .q(_divSqrt_single__q),
        .d(_divSqrt_single__d),
        .clk(clock)
    );
    wire [64:0] divSqrt_wdata;
    wire [4:0] divSqrt_flags;
    wire _divSqrt_in_flight__q;
    wire _divSqrt_in_flight__d;
    DFF_POSCLK #(.width(1)) divSqrt_in_flight (
        .q(_divSqrt_in_flight__q),
        .d(_divSqrt_in_flight__d),
        .clk(clock)
    );
    wire _WTEMP_477;
    MUX_UNSIGNED #(.width(1)) u_mux_3478 (
        .y(_divSqrt_in_flight__d),
        .sel(reset),
        .a(1'h0),
        .b(_WTEMP_477)
    );
    wire _divSqrt_killed__q;
    wire _divSqrt_killed__d;
    DFF_POSCLK #(.width(1)) divSqrt_killed (
        .q(_divSqrt_killed__q),
        .d(_divSqrt_killed__d),
        .clk(clock)
    );
    wire _FPUFMAPipe__clock;
    wire _FPUFMAPipe__reset;
    wire _FPUFMAPipe__io_in_valid;
    wire [4:0] _FPUFMAPipe__io_in_bits_cmd;
    wire _FPUFMAPipe__io_in_bits_ldst;
    wire _FPUFMAPipe__io_in_bits_wen;
    wire _FPUFMAPipe__io_in_bits_ren1;
    wire _FPUFMAPipe__io_in_bits_ren2;
    wire _FPUFMAPipe__io_in_bits_ren3;
    wire _FPUFMAPipe__io_in_bits_swap12;
    wire _FPUFMAPipe__io_in_bits_swap23;
    wire _FPUFMAPipe__io_in_bits_single;
    wire _FPUFMAPipe__io_in_bits_fromint;
    wire _FPUFMAPipe__io_in_bits_toint;
    wire _FPUFMAPipe__io_in_bits_fastpipe;
    wire _FPUFMAPipe__io_in_bits_fma;
    wire _FPUFMAPipe__io_in_bits_div;
    wire _FPUFMAPipe__io_in_bits_sqrt;
    wire _FPUFMAPipe__io_in_bits_wflags;
    wire [2:0] _FPUFMAPipe__io_in_bits_rm;
    wire [1:0] _FPUFMAPipe__io_in_bits_typ;
    wire [64:0] _FPUFMAPipe__io_in_bits_in1;
    wire [64:0] _FPUFMAPipe__io_in_bits_in2;
    wire [64:0] _FPUFMAPipe__io_in_bits_in3;
    wire _FPUFMAPipe__io_out_valid;
    wire [64:0] _FPUFMAPipe__io_out_bits_data;
    wire [4:0] _FPUFMAPipe__io_out_bits_exc;
    FPUFMAPipe_1 FPUFMAPipe (
        .clock(_FPUFMAPipe__clock),
        .reset(_FPUFMAPipe__reset),
        .io_in_valid(_FPUFMAPipe__io_in_valid),
        .io_in_bits_cmd(_FPUFMAPipe__io_in_bits_cmd),
        .io_in_bits_ldst(_FPUFMAPipe__io_in_bits_ldst),
        .io_in_bits_wen(_FPUFMAPipe__io_in_bits_wen),
        .io_in_bits_ren1(_FPUFMAPipe__io_in_bits_ren1),
        .io_in_bits_ren2(_FPUFMAPipe__io_in_bits_ren2),
        .io_in_bits_ren3(_FPUFMAPipe__io_in_bits_ren3),
        .io_in_bits_swap12(_FPUFMAPipe__io_in_bits_swap12),
        .io_in_bits_swap23(_FPUFMAPipe__io_in_bits_swap23),
        .io_in_bits_single(_FPUFMAPipe__io_in_bits_single),
        .io_in_bits_fromint(_FPUFMAPipe__io_in_bits_fromint),
        .io_in_bits_toint(_FPUFMAPipe__io_in_bits_toint),
        .io_in_bits_fastpipe(_FPUFMAPipe__io_in_bits_fastpipe),
        .io_in_bits_fma(_FPUFMAPipe__io_in_bits_fma),
        .io_in_bits_div(_FPUFMAPipe__io_in_bits_div),
        .io_in_bits_sqrt(_FPUFMAPipe__io_in_bits_sqrt),
        .io_in_bits_wflags(_FPUFMAPipe__io_in_bits_wflags),
        .io_in_bits_rm(_FPUFMAPipe__io_in_bits_rm),
        .io_in_bits_typ(_FPUFMAPipe__io_in_bits_typ),
        .io_in_bits_in1(_FPUFMAPipe__io_in_bits_in1),
        .io_in_bits_in2(_FPUFMAPipe__io_in_bits_in2),
        .io_in_bits_in3(_FPUFMAPipe__io_in_bits_in3),
        .io_out_valid(_FPUFMAPipe__io_out_valid),
        .io_out_bits_data(_FPUFMAPipe__io_out_bits_data),
        .io_out_bits_exc(_FPUFMAPipe__io_out_bits_exc)
    );
    wire _T_883;
    BITWISEAND #(.width(1)) bitwiseand_4694 (
        .y(_T_883),
        .a(req_valid),
        .b(ex_ctrl_fma)
    );
    wire _T_885;
    EQ_UNSIGNED #(.width(1)) u_eq_4695 (
        .y(_T_885),
        .a(ex_ctrl_single),
        .b(1'h0)
    );
    wire _T_886;
    BITWISEAND #(.width(1)) bitwiseand_4696 (
        .y(_T_886),
        .a(_T_883),
        .b(_T_885)
    );
    wire _T_889;
    MUX_UNSIGNED #(.width(1)) u_mux_4697 (
        .y(_T_889),
        .sel(_mem_ctrl_fastpipe__q),
        .a(1'h1),
        .b(1'h0)
    );
    wire _T_892;
    MUX_UNSIGNED #(.width(1)) u_mux_4698 (
        .y(_T_892),
        .sel(_mem_ctrl_fromint__q),
        .a(1'h1),
        .b(1'h0)
    );
    wire _T_893;
    BITWISEAND #(.width(1)) bitwiseand_4699 (
        .y(_T_893),
        .a(_mem_ctrl_fma__q),
        .b(_mem_ctrl_single__q)
    );
    wire [1:0] _T_896;
    wire [1:0] _WTEMP_646;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_4700 (
        .y(_WTEMP_646),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_4701 (
        .y(_T_896),
        .sel(_T_893),
        .a(2'h2),
        .b(_WTEMP_646)
    );
    wire _T_898;
    EQ_UNSIGNED #(.width(1)) u_eq_4702 (
        .y(_T_898),
        .a(_mem_ctrl_single__q),
        .b(1'h0)
    );
    wire _T_899;
    BITWISEAND #(.width(1)) bitwiseand_4703 (
        .y(_T_899),
        .a(_mem_ctrl_fma__q),
        .b(_T_898)
    );
    wire [2:0] _T_902;
    wire [2:0] _WTEMP_647;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_4704 (
        .y(_WTEMP_647),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(3)) u_mux_4705 (
        .y(_T_902),
        .sel(_T_899),
        .a(3'h4),
        .b(_WTEMP_647)
    );
    wire _T_903;
    BITWISEOR #(.width(1)) bitwiseor_4706 (
        .y(_T_903),
        .a(_T_889),
        .b(_T_892)
    );
    wire [1:0] _T_904;
    wire [1:0] _WTEMP_648;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_4707 (
        .y(_WTEMP_648),
        .in(_T_903)
    );
    BITWISEOR #(.width(2)) bitwiseor_4708 (
        .y(_T_904),
        .a(_WTEMP_648),
        .b(_T_896)
    );
    wire [2:0] memLatencyMask;
    wire [2:0] _WTEMP_649;
    PAD_UNSIGNED #(.width(2), .n(3)) u_pad_4709 (
        .y(_WTEMP_649),
        .in(_T_904)
    );
    BITWISEOR #(.width(3)) bitwiseor_4710 (
        .y(memLatencyMask),
        .a(_WTEMP_649),
        .b(_T_902)
    );
    wire [2:0] _wen__q;
    wire [2:0] _wen__d;
    DFF_POSCLK #(.width(3)) wen (
        .q(_wen__q),
        .d(_wen__d),
        .clk(clock)
    );
    wire [2:0] _WTEMP_650;
    MUX_UNSIGNED #(.width(3)) u_mux_4711 (
        .y(_wen__d),
        .sel(reset),
        .a(3'h0),
        .b(_WTEMP_650)
    );
    wire [4:0] _wbInfo_0_rd__q;
    wire [4:0] _wbInfo_0_rd__d;
    DFF_POSCLK #(.width(5)) wbInfo_0_rd (
        .q(_wbInfo_0_rd__q),
        .d(_wbInfo_0_rd__d),
        .clk(clock)
    );
    wire _wbInfo_0_single__q;
    wire _wbInfo_0_single__d;
    DFF_POSCLK #(.width(1)) wbInfo_0_single (
        .q(_wbInfo_0_single__q),
        .d(_wbInfo_0_single__d),
        .clk(clock)
    );
    wire _wbInfo_0_cp__q;
    wire _wbInfo_0_cp__d;
    DFF_POSCLK #(.width(1)) wbInfo_0_cp (
        .q(_wbInfo_0_cp__q),
        .d(_wbInfo_0_cp__d),
        .clk(clock)
    );
    wire [1:0] _wbInfo_0_pipeid__q;
    wire [1:0] _wbInfo_0_pipeid__d;
    DFF_POSCLK #(.width(2)) wbInfo_0_pipeid (
        .q(_wbInfo_0_pipeid__q),
        .d(_wbInfo_0_pipeid__d),
        .clk(clock)
    );
    wire [4:0] _wbInfo_1_rd__q;
    wire [4:0] _wbInfo_1_rd__d;
    DFF_POSCLK #(.width(5)) wbInfo_1_rd (
        .q(_wbInfo_1_rd__q),
        .d(_wbInfo_1_rd__d),
        .clk(clock)
    );
    wire _wbInfo_1_single__q;
    wire _wbInfo_1_single__d;
    DFF_POSCLK #(.width(1)) wbInfo_1_single (
        .q(_wbInfo_1_single__q),
        .d(_wbInfo_1_single__d),
        .clk(clock)
    );
    wire _wbInfo_1_cp__q;
    wire _wbInfo_1_cp__d;
    DFF_POSCLK #(.width(1)) wbInfo_1_cp (
        .q(_wbInfo_1_cp__q),
        .d(_wbInfo_1_cp__d),
        .clk(clock)
    );
    wire [1:0] _wbInfo_1_pipeid__q;
    wire [1:0] _wbInfo_1_pipeid__d;
    DFF_POSCLK #(.width(2)) wbInfo_1_pipeid (
        .q(_wbInfo_1_pipeid__q),
        .d(_wbInfo_1_pipeid__d),
        .clk(clock)
    );
    wire [4:0] _wbInfo_2_rd__q;
    wire [4:0] _wbInfo_2_rd__d;
    DFF_POSCLK #(.width(5)) wbInfo_2_rd (
        .q(_wbInfo_2_rd__q),
        .d(_wbInfo_2_rd__d),
        .clk(clock)
    );
    wire _wbInfo_2_single__q;
    wire _wbInfo_2_single__d;
    DFF_POSCLK #(.width(1)) wbInfo_2_single (
        .q(_wbInfo_2_single__q),
        .d(_wbInfo_2_single__d),
        .clk(clock)
    );
    wire _wbInfo_2_cp__q;
    wire _wbInfo_2_cp__d;
    DFF_POSCLK #(.width(1)) wbInfo_2_cp (
        .q(_wbInfo_2_cp__q),
        .d(_wbInfo_2_cp__d),
        .clk(clock)
    );
    wire [1:0] _wbInfo_2_pipeid__q;
    wire [1:0] _wbInfo_2_pipeid__d;
    DFF_POSCLK #(.width(2)) wbInfo_2_pipeid (
        .q(_wbInfo_2_pipeid__q),
        .d(_wbInfo_2_pipeid__d),
        .clk(clock)
    );
    wire _T_966;
    BITWISEOR #(.width(1)) bitwiseor_4712 (
        .y(_T_966),
        .a(_mem_ctrl_fma__q),
        .b(_mem_ctrl_fastpipe__q)
    );
    wire _T_967;
    BITWISEOR #(.width(1)) bitwiseor_4713 (
        .y(_T_967),
        .a(_T_966),
        .b(_mem_ctrl_fromint__q)
    );
    wire mem_wen;
    BITWISEAND #(.width(1)) bitwiseand_4714 (
        .y(mem_wen),
        .a(_mem_reg_valid__q),
        .b(_T_967)
    );
    wire [1:0] _T_970;
    wire [1:0] _WTEMP_651;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_4715 (
        .y(_WTEMP_651),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_4716 (
        .y(_T_970),
        .sel(ex_ctrl_fastpipe),
        .a(2'h2),
        .b(_WTEMP_651)
    );
    wire [1:0] _T_973;
    wire [1:0] _WTEMP_652;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_4717 (
        .y(_WTEMP_652),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_4718 (
        .y(_T_973),
        .sel(ex_ctrl_fromint),
        .a(2'h2),
        .b(_WTEMP_652)
    );
    wire _T_974;
    BITWISEAND #(.width(1)) bitwiseand_4719 (
        .y(_T_974),
        .a(ex_ctrl_fma),
        .b(ex_ctrl_single)
    );
    wire [2:0] _T_977;
    wire [2:0] _WTEMP_653;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_4720 (
        .y(_WTEMP_653),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(3)) u_mux_4721 (
        .y(_T_977),
        .sel(_T_974),
        .a(3'h4),
        .b(_WTEMP_653)
    );
    wire _T_979;
    EQ_UNSIGNED #(.width(1)) u_eq_4722 (
        .y(_T_979),
        .a(ex_ctrl_single),
        .b(1'h0)
    );
    wire _T_980;
    BITWISEAND #(.width(1)) bitwiseand_4723 (
        .y(_T_980),
        .a(ex_ctrl_fma),
        .b(_T_979)
    );
    wire [3:0] _T_983;
    wire [3:0] _WTEMP_654;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_4724 (
        .y(_WTEMP_654),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(4)) u_mux_4725 (
        .y(_T_983),
        .sel(_T_980),
        .a(4'h8),
        .b(_WTEMP_654)
    );
    wire [1:0] _T_984;
    BITWISEOR #(.width(2)) bitwiseor_4726 (
        .y(_T_984),
        .a(_T_970),
        .b(_T_973)
    );
    wire [2:0] _T_985;
    wire [2:0] _WTEMP_655;
    PAD_UNSIGNED #(.width(2), .n(3)) u_pad_4727 (
        .y(_WTEMP_655),
        .in(_T_984)
    );
    BITWISEOR #(.width(3)) bitwiseor_4728 (
        .y(_T_985),
        .a(_WTEMP_655),
        .b(_T_977)
    );
    wire [3:0] _T_986;
    wire [3:0] _WTEMP_656;
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_4729 (
        .y(_WTEMP_656),
        .in(_T_985)
    );
    BITWISEOR #(.width(4)) bitwiseor_4730 (
        .y(_T_986),
        .a(_WTEMP_656),
        .b(_T_983)
    );
    wire [3:0] _T_987;
    wire [3:0] _WTEMP_657;
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_4731 (
        .y(_WTEMP_657),
        .in(memLatencyMask)
    );
    BITWISEAND #(.width(4)) bitwiseand_4732 (
        .y(_T_987),
        .a(_WTEMP_657),
        .b(_T_986)
    );
    wire _T_989;
    wire [3:0] _WTEMP_658;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_4733 (
        .y(_WTEMP_658),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_4734 (
        .y(_T_989),
        .a(_T_987),
        .b(_WTEMP_658)
    );
    wire _T_990;
    BITWISEAND #(.width(1)) bitwiseand_4735 (
        .y(_T_990),
        .a(mem_wen),
        .b(_T_989)
    );
    wire [2:0] _T_993;
    wire [2:0] _WTEMP_659;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_4736 (
        .y(_WTEMP_659),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(3)) u_mux_4737 (
        .y(_T_993),
        .sel(ex_ctrl_fastpipe),
        .a(3'h4),
        .b(_WTEMP_659)
    );
    wire [2:0] _T_996;
    wire [2:0] _WTEMP_660;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_4738 (
        .y(_WTEMP_660),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(3)) u_mux_4739 (
        .y(_T_996),
        .sel(ex_ctrl_fromint),
        .a(3'h4),
        .b(_WTEMP_660)
    );
    wire _T_997;
    BITWISEAND #(.width(1)) bitwiseand_4740 (
        .y(_T_997),
        .a(ex_ctrl_fma),
        .b(ex_ctrl_single)
    );
    wire [3:0] _T_1000;
    wire [3:0] _WTEMP_661;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_4741 (
        .y(_WTEMP_661),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(4)) u_mux_4742 (
        .y(_T_1000),
        .sel(_T_997),
        .a(4'h8),
        .b(_WTEMP_661)
    );
    wire _T_1002;
    EQ_UNSIGNED #(.width(1)) u_eq_4743 (
        .y(_T_1002),
        .a(ex_ctrl_single),
        .b(1'h0)
    );
    wire _T_1003;
    BITWISEAND #(.width(1)) bitwiseand_4744 (
        .y(_T_1003),
        .a(ex_ctrl_fma),
        .b(_T_1002)
    );
    wire [4:0] _T_1006;
    wire [4:0] _WTEMP_662;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_4745 (
        .y(_WTEMP_662),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(5)) u_mux_4746 (
        .y(_T_1006),
        .sel(_T_1003),
        .a(5'h10),
        .b(_WTEMP_662)
    );
    wire [2:0] _T_1007;
    BITWISEOR #(.width(3)) bitwiseor_4747 (
        .y(_T_1007),
        .a(_T_993),
        .b(_T_996)
    );
    wire [3:0] _T_1008;
    wire [3:0] _WTEMP_663;
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_4748 (
        .y(_WTEMP_663),
        .in(_T_1007)
    );
    BITWISEOR #(.width(4)) bitwiseor_4749 (
        .y(_T_1008),
        .a(_WTEMP_663),
        .b(_T_1000)
    );
    wire [4:0] _T_1009;
    wire [4:0] _WTEMP_664;
    PAD_UNSIGNED #(.width(4), .n(5)) u_pad_4750 (
        .y(_WTEMP_664),
        .in(_T_1008)
    );
    BITWISEOR #(.width(5)) bitwiseor_4751 (
        .y(_T_1009),
        .a(_WTEMP_664),
        .b(_T_1006)
    );
    wire [4:0] _T_1010;
    wire [4:0] _WTEMP_665;
    PAD_UNSIGNED #(.width(3), .n(5)) u_pad_4752 (
        .y(_WTEMP_665),
        .in(_wen__q)
    );
    BITWISEAND #(.width(5)) bitwiseand_4753 (
        .y(_T_1010),
        .a(_WTEMP_665),
        .b(_T_1009)
    );
    wire _T_1012;
    wire [4:0] _WTEMP_666;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_4754 (
        .y(_WTEMP_666),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(5)) u_neq_4755 (
        .y(_T_1012),
        .a(_T_1010),
        .b(_WTEMP_666)
    );
    wire _T_1013;
    BITWISEOR #(.width(1)) bitwiseor_4756 (
        .y(_T_1013),
        .a(_T_990),
        .b(_T_1012)
    );
    wire _write_port_busy__q;
    wire _write_port_busy__d;
    DFF_POSCLK #(.width(1)) write_port_busy (
        .q(_write_port_busy__q),
        .d(_write_port_busy__d),
        .clk(clock)
    );
    wire _T_1015;
    BITS #(.width(3), .high(1), .low(1)) bits_4757 (
        .y(_T_1015),
        .in(_wen__q)
    );
    wire _T_1016;
    BITS #(.width(3), .high(2), .low(2)) bits_4758 (
        .y(_T_1016),
        .in(_wen__q)
    );
    wire [1:0] _T_1017;
    SHR_UNSIGNED #(.width(3), .n(1)) u_shr_4759 (
        .y(_T_1017),
        .in(_wen__q)
    );
    wire _T_1019;
    EQ_UNSIGNED #(.width(1)) u_eq_4760 (
        .y(_T_1019),
        .a(killm),
        .b(1'h0)
    );
    wire [1:0] _T_1020;
    SHR_UNSIGNED #(.width(3), .n(1)) u_shr_4761 (
        .y(_T_1020),
        .in(_wen__q)
    );
    wire [2:0] _T_1021;
    wire [2:0] _WTEMP_667;
    PAD_UNSIGNED #(.width(2), .n(3)) u_pad_4762 (
        .y(_WTEMP_667),
        .in(_T_1020)
    );
    BITWISEOR #(.width(3)) bitwiseor_4763 (
        .y(_T_1021),
        .a(_WTEMP_667),
        .b(memLatencyMask)
    );
    wire _T_1023;
    EQ_UNSIGNED #(.width(1)) u_eq_4764 (
        .y(_T_1023),
        .a(_write_port_busy__q),
        .b(1'h0)
    );
    wire _T_1024;
    BITS #(.width(3), .high(0), .low(0)) bits_4765 (
        .y(_T_1024),
        .in(memLatencyMask)
    );
    wire _T_1025;
    BITWISEAND #(.width(1)) bitwiseand_4766 (
        .y(_T_1025),
        .a(_T_1023),
        .b(_T_1024)
    );
    wire _T_1028;
    assign _T_1028 = 1'h0;
    wire _T_1031;
    MUX_UNSIGNED #(.width(1)) u_mux_4767 (
        .y(_T_1031),
        .sel(_mem_ctrl_fromint__q),
        .a(1'h1),
        .b(1'h0)
    );
    wire _T_1032;
    BITWISEAND #(.width(1)) bitwiseand_4768 (
        .y(_T_1032),
        .a(_mem_ctrl_fma__q),
        .b(_mem_ctrl_single__q)
    );
    wire [1:0] _T_1035;
    wire [1:0] _WTEMP_668;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_4769 (
        .y(_WTEMP_668),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_4770 (
        .y(_T_1035),
        .sel(_T_1032),
        .a(2'h2),
        .b(_WTEMP_668)
    );
    wire _T_1037;
    EQ_UNSIGNED #(.width(1)) u_eq_4771 (
        .y(_T_1037),
        .a(_mem_ctrl_single__q),
        .b(1'h0)
    );
    wire _T_1038;
    BITWISEAND #(.width(1)) bitwiseand_4772 (
        .y(_T_1038),
        .a(_mem_ctrl_fma__q),
        .b(_T_1037)
    );
    wire [1:0] _T_1041;
    wire [1:0] _WTEMP_669;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_4773 (
        .y(_WTEMP_669),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_4774 (
        .y(_T_1041),
        .sel(_T_1038),
        .a(2'h3),
        .b(_WTEMP_669)
    );
    wire _T_1042;
    BITWISEOR #(.width(1)) bitwiseor_4775 (
        .y(_T_1042),
        .a(_T_1028),
        .b(_T_1031)
    );
    wire [1:0] _T_1043;
    wire [1:0] _WTEMP_670;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_4776 (
        .y(_WTEMP_670),
        .in(_T_1042)
    );
    BITWISEOR #(.width(2)) bitwiseor_4777 (
        .y(_T_1043),
        .a(_WTEMP_670),
        .b(_T_1035)
    );
    wire [1:0] _T_1044;
    BITWISEOR #(.width(2)) bitwiseor_4778 (
        .y(_T_1044),
        .a(_T_1043),
        .b(_T_1041)
    );
    wire [4:0] _T_1045;
    BITS #(.width(32), .high(11), .low(7)) bits_4779 (
        .y(_T_1045),
        .in(_mem_reg_inst__q)
    );
    wire _node_40;
    MUX_UNSIGNED #(.width(1)) u_mux_4780 (
        .y(_node_40),
        .sel(_T_1015),
        .a(_wbInfo_1_cp__q),
        .b(_wbInfo_0_cp__q)
    );
    wire [1:0] _node_41;
    MUX_UNSIGNED #(.width(2)) u_mux_4781 (
        .y(_node_41),
        .sel(_T_1015),
        .a(_wbInfo_1_pipeid__q),
        .b(_wbInfo_0_pipeid__q)
    );
    wire [4:0] _node_42;
    MUX_UNSIGNED #(.width(5)) u_mux_4782 (
        .y(_node_42),
        .sel(_T_1015),
        .a(_wbInfo_1_rd__q),
        .b(_wbInfo_0_rd__q)
    );
    wire _node_43;
    MUX_UNSIGNED #(.width(1)) u_mux_4783 (
        .y(_node_43),
        .sel(_T_1015),
        .a(_wbInfo_1_single__q),
        .b(_wbInfo_0_single__q)
    );
    wire _T_1047;
    EQ_UNSIGNED #(.width(1)) u_eq_4784 (
        .y(_T_1047),
        .a(_write_port_busy__q),
        .b(1'h0)
    );
    wire _T_1048;
    BITS #(.width(3), .high(1), .low(1)) bits_4785 (
        .y(_T_1048),
        .in(memLatencyMask)
    );
    wire _T_1049;
    BITWISEAND #(.width(1)) bitwiseand_4786 (
        .y(_T_1049),
        .a(_T_1047),
        .b(_T_1048)
    );
    wire _T_1052;
    assign _T_1052 = 1'h0;
    wire _T_1055;
    MUX_UNSIGNED #(.width(1)) u_mux_4787 (
        .y(_T_1055),
        .sel(_mem_ctrl_fromint__q),
        .a(1'h1),
        .b(1'h0)
    );
    wire _T_1056;
    BITWISEAND #(.width(1)) bitwiseand_4788 (
        .y(_T_1056),
        .a(_mem_ctrl_fma__q),
        .b(_mem_ctrl_single__q)
    );
    wire [1:0] _T_1059;
    wire [1:0] _WTEMP_671;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_4789 (
        .y(_WTEMP_671),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_4790 (
        .y(_T_1059),
        .sel(_T_1056),
        .a(2'h2),
        .b(_WTEMP_671)
    );
    wire _T_1061;
    EQ_UNSIGNED #(.width(1)) u_eq_4791 (
        .y(_T_1061),
        .a(_mem_ctrl_single__q),
        .b(1'h0)
    );
    wire _T_1062;
    BITWISEAND #(.width(1)) bitwiseand_4792 (
        .y(_T_1062),
        .a(_mem_ctrl_fma__q),
        .b(_T_1061)
    );
    wire [1:0] _T_1065;
    wire [1:0] _WTEMP_672;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_4793 (
        .y(_WTEMP_672),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_4794 (
        .y(_T_1065),
        .sel(_T_1062),
        .a(2'h3),
        .b(_WTEMP_672)
    );
    wire _T_1066;
    BITWISEOR #(.width(1)) bitwiseor_4795 (
        .y(_T_1066),
        .a(_T_1052),
        .b(_T_1055)
    );
    wire [1:0] _T_1067;
    wire [1:0] _WTEMP_673;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_4796 (
        .y(_WTEMP_673),
        .in(_T_1066)
    );
    BITWISEOR #(.width(2)) bitwiseor_4797 (
        .y(_T_1067),
        .a(_WTEMP_673),
        .b(_T_1059)
    );
    wire [1:0] _T_1068;
    BITWISEOR #(.width(2)) bitwiseor_4798 (
        .y(_T_1068),
        .a(_T_1067),
        .b(_T_1065)
    );
    wire [4:0] _T_1069;
    BITS #(.width(32), .high(11), .low(7)) bits_4799 (
        .y(_T_1069),
        .in(_mem_reg_inst__q)
    );
    wire _node_44;
    MUX_UNSIGNED #(.width(1)) u_mux_4800 (
        .y(_node_44),
        .sel(_T_1016),
        .a(_wbInfo_2_cp__q),
        .b(_wbInfo_1_cp__q)
    );
    wire [1:0] _node_45;
    MUX_UNSIGNED #(.width(2)) u_mux_4801 (
        .y(_node_45),
        .sel(_T_1016),
        .a(_wbInfo_2_pipeid__q),
        .b(_wbInfo_1_pipeid__q)
    );
    wire [4:0] _node_46;
    MUX_UNSIGNED #(.width(5)) u_mux_4802 (
        .y(_node_46),
        .sel(_T_1016),
        .a(_wbInfo_2_rd__q),
        .b(_wbInfo_1_rd__q)
    );
    wire _node_47;
    MUX_UNSIGNED #(.width(1)) u_mux_4803 (
        .y(_node_47),
        .sel(_T_1016),
        .a(_wbInfo_2_single__q),
        .b(_wbInfo_1_single__q)
    );
    wire _T_1071;
    EQ_UNSIGNED #(.width(1)) u_eq_4804 (
        .y(_T_1071),
        .a(_write_port_busy__q),
        .b(1'h0)
    );
    wire _T_1072;
    BITS #(.width(3), .high(2), .low(2)) bits_4805 (
        .y(_T_1072),
        .in(memLatencyMask)
    );
    wire _T_1073;
    BITWISEAND #(.width(1)) bitwiseand_4806 (
        .y(_T_1073),
        .a(_T_1071),
        .b(_T_1072)
    );
    wire _T_1076;
    assign _T_1076 = 1'h0;
    wire _T_1079;
    MUX_UNSIGNED #(.width(1)) u_mux_4807 (
        .y(_T_1079),
        .sel(_mem_ctrl_fromint__q),
        .a(1'h1),
        .b(1'h0)
    );
    wire _T_1080;
    BITWISEAND #(.width(1)) bitwiseand_4808 (
        .y(_T_1080),
        .a(_mem_ctrl_fma__q),
        .b(_mem_ctrl_single__q)
    );
    wire [1:0] _T_1083;
    wire [1:0] _WTEMP_674;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_4809 (
        .y(_WTEMP_674),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_4810 (
        .y(_T_1083),
        .sel(_T_1080),
        .a(2'h2),
        .b(_WTEMP_674)
    );
    wire _T_1085;
    EQ_UNSIGNED #(.width(1)) u_eq_4811 (
        .y(_T_1085),
        .a(_mem_ctrl_single__q),
        .b(1'h0)
    );
    wire _T_1086;
    BITWISEAND #(.width(1)) bitwiseand_4812 (
        .y(_T_1086),
        .a(_mem_ctrl_fma__q),
        .b(_T_1085)
    );
    wire [1:0] _T_1089;
    wire [1:0] _WTEMP_675;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_4813 (
        .y(_WTEMP_675),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_4814 (
        .y(_T_1089),
        .sel(_T_1086),
        .a(2'h3),
        .b(_WTEMP_675)
    );
    wire _T_1090;
    BITWISEOR #(.width(1)) bitwiseor_4815 (
        .y(_T_1090),
        .a(_T_1076),
        .b(_T_1079)
    );
    wire [1:0] _T_1091;
    wire [1:0] _WTEMP_676;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_4816 (
        .y(_WTEMP_676),
        .in(_T_1090)
    );
    BITWISEOR #(.width(2)) bitwiseor_4817 (
        .y(_T_1091),
        .a(_WTEMP_676),
        .b(_T_1083)
    );
    wire [1:0] _T_1092;
    BITWISEOR #(.width(2)) bitwiseor_4818 (
        .y(_T_1092),
        .a(_T_1091),
        .b(_T_1089)
    );
    wire [4:0] _T_1093;
    BITS #(.width(32), .high(11), .low(7)) bits_4819 (
        .y(_T_1093),
        .in(_mem_reg_inst__q)
    );
    wire _node_48;
    MUX_UNSIGNED #(.width(1)) u_mux_4820 (
        .y(_node_48),
        .sel(_T_1025),
        .a(_mem_cp_valid__q),
        .b(_node_40)
    );
    wire _node_49;
    MUX_UNSIGNED #(.width(1)) u_mux_4821 (
        .y(_node_49),
        .sel(_T_1015),
        .a(_wbInfo_1_cp__q),
        .b(_wbInfo_0_cp__q)
    );
    wire [1:0] _node_50;
    MUX_UNSIGNED #(.width(2)) u_mux_4822 (
        .y(_node_50),
        .sel(_T_1025),
        .a(_T_1044),
        .b(_node_41)
    );
    wire [1:0] _node_51;
    MUX_UNSIGNED #(.width(2)) u_mux_4823 (
        .y(_node_51),
        .sel(_T_1015),
        .a(_wbInfo_1_pipeid__q),
        .b(_wbInfo_0_pipeid__q)
    );
    wire [4:0] _node_52;
    MUX_UNSIGNED #(.width(5)) u_mux_4824 (
        .y(_node_52),
        .sel(_T_1025),
        .a(_T_1045),
        .b(_node_42)
    );
    wire [4:0] _node_53;
    MUX_UNSIGNED #(.width(5)) u_mux_4825 (
        .y(_node_53),
        .sel(_T_1015),
        .a(_wbInfo_1_rd__q),
        .b(_wbInfo_0_rd__q)
    );
    wire _node_54;
    MUX_UNSIGNED #(.width(1)) u_mux_4826 (
        .y(_node_54),
        .sel(_T_1025),
        .a(_mem_ctrl_single__q),
        .b(_node_43)
    );
    wire _node_55;
    MUX_UNSIGNED #(.width(1)) u_mux_4827 (
        .y(_node_55),
        .sel(_T_1015),
        .a(_wbInfo_1_single__q),
        .b(_wbInfo_0_single__q)
    );
    wire _node_56;
    MUX_UNSIGNED #(.width(1)) u_mux_4828 (
        .y(_node_56),
        .sel(_T_1049),
        .a(_mem_cp_valid__q),
        .b(_node_44)
    );
    wire _node_57;
    MUX_UNSIGNED #(.width(1)) u_mux_4829 (
        .y(_node_57),
        .sel(_T_1016),
        .a(_wbInfo_2_cp__q),
        .b(_wbInfo_1_cp__q)
    );
    wire [1:0] _node_58;
    MUX_UNSIGNED #(.width(2)) u_mux_4830 (
        .y(_node_58),
        .sel(_T_1049),
        .a(_T_1068),
        .b(_node_45)
    );
    wire [1:0] _node_59;
    MUX_UNSIGNED #(.width(2)) u_mux_4831 (
        .y(_node_59),
        .sel(_T_1016),
        .a(_wbInfo_2_pipeid__q),
        .b(_wbInfo_1_pipeid__q)
    );
    wire [4:0] _node_60;
    MUX_UNSIGNED #(.width(5)) u_mux_4832 (
        .y(_node_60),
        .sel(_T_1049),
        .a(_T_1069),
        .b(_node_46)
    );
    wire [4:0] _node_61;
    MUX_UNSIGNED #(.width(5)) u_mux_4833 (
        .y(_node_61),
        .sel(_T_1016),
        .a(_wbInfo_2_rd__q),
        .b(_wbInfo_1_rd__q)
    );
    wire _node_62;
    MUX_UNSIGNED #(.width(1)) u_mux_4834 (
        .y(_node_62),
        .sel(_T_1049),
        .a(_mem_ctrl_single__q),
        .b(_node_47)
    );
    wire _node_63;
    MUX_UNSIGNED #(.width(1)) u_mux_4835 (
        .y(_node_63),
        .sel(_T_1016),
        .a(_wbInfo_2_single__q),
        .b(_wbInfo_1_single__q)
    );
    wire _node_64;
    MUX_UNSIGNED #(.width(1)) u_mux_4836 (
        .y(_node_64),
        .sel(_T_1073),
        .a(_mem_cp_valid__q),
        .b(_wbInfo_2_cp__q)
    );
    wire [1:0] _node_65;
    MUX_UNSIGNED #(.width(2)) u_mux_4837 (
        .y(_node_65),
        .sel(_T_1073),
        .a(_T_1092),
        .b(_wbInfo_2_pipeid__q)
    );
    wire [4:0] _node_66;
    MUX_UNSIGNED #(.width(5)) u_mux_4838 (
        .y(_node_66),
        .sel(_T_1073),
        .a(_T_1093),
        .b(_wbInfo_2_rd__q)
    );
    wire _node_67;
    MUX_UNSIGNED #(.width(1)) u_mux_4839 (
        .y(_node_67),
        .sel(_T_1073),
        .a(_mem_ctrl_single__q),
        .b(_wbInfo_2_single__q)
    );
    wire [2:0] _node_68;
    wire [2:0] _WTEMP_677;
    PAD_UNSIGNED #(.width(2), .n(3)) u_pad_4840 (
        .y(_WTEMP_677),
        .in(_T_1017)
    );
    MUX_UNSIGNED #(.width(3)) u_mux_4841 (
        .y(_node_68),
        .sel(_T_1019),
        .a(_T_1021),
        .b(_WTEMP_677)
    );
    wire [4:0] waddr;
    MUX_UNSIGNED #(.width(5)) u_mux_4842 (
        .y(waddr),
        .sel(_divSqrt_wen__q),
        .a(_divSqrt_waddr__q),
        .b(_wbInfo_0_rd__q)
    );
    wire [1:0] _T_1095;
    wire [1:0] _WTEMP_678;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_4843 (
        .y(_WTEMP_678),
        .in(1'h1)
    );
    BITWISEAND #(.width(2)) bitwiseand_4844 (
        .y(_T_1095),
        .a(_wbInfo_0_pipeid__q),
        .b(_WTEMP_678)
    );
    wire _T_1097;
    GEQ_UNSIGNED #(.width(2)) u_geq_4845 (
        .y(_T_1097),
        .a(_wbInfo_0_pipeid__q),
        .b(2'h2)
    );
    wire [1:0] _T_1099;
    assign _T_1099 = 2'h0;
    wire _T_1101;
    wire [1:0] _WTEMP_679;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_4846 (
        .y(_WTEMP_679),
        .in(1'h1)
    );
    GEQ_UNSIGNED #(.width(2)) u_geq_4847 (
        .y(_T_1101),
        .a(_T_1095),
        .b(_WTEMP_679)
    );
    wire [64:0] _T_1102;
    MUX_UNSIGNED #(.width(65)) u_mux_4848 (
        .y(_T_1102),
        .sel(_T_1101),
        .a(_FPUFMAPipe__io_out_bits_data),
        .b(_sfma__io_out_bits_data)
    );
    wire [1:0] _T_1104;
    assign _T_1104 = 2'h0;
    wire _T_1106;
    wire [1:0] _WTEMP_680;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_4849 (
        .y(_WTEMP_680),
        .in(1'h1)
    );
    GEQ_UNSIGNED #(.width(2)) u_geq_4850 (
        .y(_T_1106),
        .a(_T_1095),
        .b(_WTEMP_680)
    );
    wire [64:0] _T_1107;
    MUX_UNSIGNED #(.width(65)) u_mux_4851 (
        .y(_T_1107),
        .sel(_T_1106),
        .a(_ifpu__io_out_bits_data),
        .b(_fpmu__io_out_bits_data)
    );
    wire [64:0] _T_1108;
    MUX_UNSIGNED #(.width(65)) u_mux_4852 (
        .y(_T_1108),
        .sel(_T_1097),
        .a(_T_1102),
        .b(_T_1107)
    );
    wire [64:0] wdata0;
    MUX_UNSIGNED #(.width(65)) u_mux_4853 (
        .y(wdata0),
        .sel(_divSqrt_wen__q),
        .a(divSqrt_wdata),
        .b(_T_1108)
    );
    wire wsingle;
    MUX_UNSIGNED #(.width(1)) u_mux_4854 (
        .y(wsingle),
        .sel(_divSqrt_wen__q),
        .a(_divSqrt_single__q),
        .b(_wbInfo_0_single__q)
    );
    wire [32:0] _T_1109;
    BITS #(.width(65), .high(32), .low(0)) bits_4855 (
        .y(_T_1109),
        .in(wdata0)
    );
    wire [64:0] _T_1111;
    wire [64:0] _WTEMP_681;
    PAD_UNSIGNED #(.width(33), .n(65)) u_pad_4856 (
        .y(_WTEMP_681),
        .in(_T_1109)
    );
    BITWISEOR #(.width(65)) bitwiseor_4857 (
        .y(_T_1111),
        .a(_WTEMP_681),
        .b(65'hE004000000000000)
    );
    wire [64:0] wdata;
    MUX_UNSIGNED #(.width(65)) u_mux_4858 (
        .y(wdata),
        .sel(wsingle),
        .a(_T_1111),
        .b(wdata0)
    );
    wire [1:0] _T_1113;
    wire [1:0] _WTEMP_682;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_4859 (
        .y(_WTEMP_682),
        .in(1'h1)
    );
    BITWISEAND #(.width(2)) bitwiseand_4860 (
        .y(_T_1113),
        .a(_wbInfo_0_pipeid__q),
        .b(_WTEMP_682)
    );
    wire _T_1115;
    GEQ_UNSIGNED #(.width(2)) u_geq_4861 (
        .y(_T_1115),
        .a(_wbInfo_0_pipeid__q),
        .b(2'h2)
    );
    wire [1:0] _T_1117;
    assign _T_1117 = 2'h0;
    wire _T_1119;
    wire [1:0] _WTEMP_683;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_4862 (
        .y(_WTEMP_683),
        .in(1'h1)
    );
    GEQ_UNSIGNED #(.width(2)) u_geq_4863 (
        .y(_T_1119),
        .a(_T_1113),
        .b(_WTEMP_683)
    );
    wire [4:0] _T_1120;
    MUX_UNSIGNED #(.width(5)) u_mux_4864 (
        .y(_T_1120),
        .sel(_T_1119),
        .a(_FPUFMAPipe__io_out_bits_exc),
        .b(_sfma__io_out_bits_exc)
    );
    wire [1:0] _T_1122;
    assign _T_1122 = 2'h0;
    wire _T_1124;
    wire [1:0] _WTEMP_684;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_4865 (
        .y(_WTEMP_684),
        .in(1'h1)
    );
    GEQ_UNSIGNED #(.width(2)) u_geq_4866 (
        .y(_T_1124),
        .a(_T_1113),
        .b(_WTEMP_684)
    );
    wire [4:0] _T_1125;
    MUX_UNSIGNED #(.width(5)) u_mux_4867 (
        .y(_T_1125),
        .sel(_T_1124),
        .a(_ifpu__io_out_bits_exc),
        .b(_fpmu__io_out_bits_exc)
    );
    wire [4:0] wexc;
    MUX_UNSIGNED #(.width(5)) u_mux_4868 (
        .y(wexc),
        .sel(_T_1115),
        .a(_T_1120),
        .b(_T_1125)
    );
    wire _T_1127;
    EQ_UNSIGNED #(.width(1)) u_eq_4869 (
        .y(_T_1127),
        .a(_wbInfo_0_cp__q),
        .b(1'h0)
    );
    wire _T_1128;
    BITS #(.width(3), .high(0), .low(0)) bits_4870 (
        .y(_T_1128),
        .in(_wen__q)
    );
    wire _T_1129;
    BITWISEAND #(.width(1)) bitwiseand_4871 (
        .y(_T_1129),
        .a(_T_1127),
        .b(_T_1128)
    );
    wire _T_1130;
    BITWISEOR #(.width(1)) bitwiseor_4872 (
        .y(_T_1130),
        .a(_T_1129),
        .b(_divSqrt_wen__q)
    );
    assign regfile__T_1131_addr = waddr;
    assign regfile__T_1131_en = _T_1130;
    assign regfile__T_1131_clk = clock;
    assign regfile__T_1131_mask = 1'h1;
    wire _T_1132;
    BITS #(.width(3), .high(0), .low(0)) bits_4873 (
        .y(_T_1132),
        .in(_wen__q)
    );
    wire _T_1133;
    BITWISEAND #(.width(1)) bitwiseand_4874 (
        .y(_T_1133),
        .a(_wbInfo_0_cp__q),
        .b(_T_1132)
    );
    wire [63:0] _node_69;
    wire [63:0] _WTEMP_685;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_4875 (
        .y(_WTEMP_685),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_4876 (
        .y(_node_69),
        .sel(_T_870),
        .a(_fpiu__io_out_bits_toint),
        .b(_WTEMP_685)
    );
    wire _node_70;
    MUX_UNSIGNED #(.width(1)) u_mux_4877 (
        .y(_node_70),
        .sel(_T_870),
        .a(1'h1),
        .b(1'h0)
    );
    wire _T_1136;
    EQ_UNSIGNED #(.width(1)) u_eq_4878 (
        .y(_T_1136),
        .a(_ex_reg_valid__q),
        .b(1'h0)
    );
    wire wb_toint_valid;
    BITWISEAND #(.width(1)) bitwiseand_4879 (
        .y(wb_toint_valid),
        .a(_wb_reg_valid__q),
        .b(_wb_ctrl_toint__q)
    );
    wire [4:0] _wb_toint_exc__q;
    wire [4:0] _wb_toint_exc__d;
    DFF_POSCLK #(.width(5)) wb_toint_exc (
        .q(_wb_toint_exc__q),
        .d(_wb_toint_exc__d),
        .clk(clock)
    );
    wire _T_1138;
    BITWISEOR #(.width(1)) bitwiseor_4880 (
        .y(_T_1138),
        .a(wb_toint_valid),
        .b(_divSqrt_wen__q)
    );
    wire _T_1139;
    BITS #(.width(3), .high(0), .low(0)) bits_4881 (
        .y(_T_1139),
        .in(_wen__q)
    );
    wire _T_1140;
    BITWISEOR #(.width(1)) bitwiseor_4882 (
        .y(_T_1140),
        .a(_T_1138),
        .b(_T_1139)
    );
    wire [4:0] _T_1142;
    wire [4:0] _WTEMP_686;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_4883 (
        .y(_WTEMP_686),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(5)) u_mux_4884 (
        .y(_T_1142),
        .sel(wb_toint_valid),
        .a(_wb_toint_exc__q),
        .b(_WTEMP_686)
    );
    wire [4:0] _T_1144;
    wire [4:0] _WTEMP_687;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_4885 (
        .y(_WTEMP_687),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(5)) u_mux_4886 (
        .y(_T_1144),
        .sel(_divSqrt_wen__q),
        .a(divSqrt_flags),
        .b(_WTEMP_687)
    );
    wire [4:0] _T_1145;
    BITWISEOR #(.width(5)) bitwiseor_4887 (
        .y(_T_1145),
        .a(_T_1142),
        .b(_T_1144)
    );
    wire _T_1146;
    BITS #(.width(3), .high(0), .low(0)) bits_4888 (
        .y(_T_1146),
        .in(_wen__q)
    );
    wire [4:0] _T_1148;
    wire [4:0] _WTEMP_688;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_4889 (
        .y(_WTEMP_688),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(5)) u_mux_4890 (
        .y(_T_1148),
        .sel(_T_1146),
        .a(wexc),
        .b(_WTEMP_688)
    );
    wire [4:0] _T_1149;
    BITWISEOR #(.width(5)) bitwiseor_4891 (
        .y(_T_1149),
        .a(_T_1145),
        .b(_T_1148)
    );
    wire _T_1150;
    BITWISEOR #(.width(1)) bitwiseor_4892 (
        .y(_T_1150),
        .a(_mem_ctrl_div__q),
        .b(_mem_ctrl_sqrt__q)
    );
    wire _T_1151;
    BITWISEAND #(.width(1)) bitwiseand_4893 (
        .y(_T_1151),
        .a(_mem_reg_valid__q),
        .b(_T_1150)
    );
    wire _T_1153;
    EQ_UNSIGNED #(.width(1)) u_eq_4894 (
        .y(_T_1153),
        .a(divSqrt_inReady),
        .b(1'h0)
    );
    wire _T_1155;
    wire [2:0] _WTEMP_689;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_4895 (
        .y(_WTEMP_689),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(3)) u_neq_4896 (
        .y(_T_1155),
        .a(_wen__q),
        .b(_WTEMP_689)
    );
    wire _T_1156;
    BITWISEOR #(.width(1)) bitwiseor_4897 (
        .y(_T_1156),
        .a(_T_1153),
        .b(_T_1155)
    );
    wire units_busy;
    BITWISEAND #(.width(1)) bitwiseand_4898 (
        .y(units_busy),
        .a(_T_1151),
        .b(_T_1156)
    );
    wire _T_1157;
    BITWISEAND #(.width(1)) bitwiseand_4899 (
        .y(_T_1157),
        .a(_ex_reg_valid__q),
        .b(ex_ctrl_wflags)
    );
    wire _T_1158;
    BITWISEAND #(.width(1)) bitwiseand_4900 (
        .y(_T_1158),
        .a(_mem_reg_valid__q),
        .b(_mem_ctrl_wflags__q)
    );
    wire _T_1159;
    BITWISEOR #(.width(1)) bitwiseor_4901 (
        .y(_T_1159),
        .a(_T_1157),
        .b(_T_1158)
    );
    wire _T_1160;
    BITWISEAND #(.width(1)) bitwiseand_4902 (
        .y(_T_1160),
        .a(_wb_reg_valid__q),
        .b(_wb_ctrl_toint__q)
    );
    wire _T_1161;
    BITWISEOR #(.width(1)) bitwiseor_4903 (
        .y(_T_1161),
        .a(_T_1159),
        .b(_T_1160)
    );
    wire _T_1163;
    wire [2:0] _WTEMP_690;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_4904 (
        .y(_WTEMP_690),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(3)) u_neq_4905 (
        .y(_T_1163),
        .a(_wen__q),
        .b(_WTEMP_690)
    );
    wire _T_1164;
    BITWISEOR #(.width(1)) bitwiseor_4906 (
        .y(_T_1164),
        .a(_T_1161),
        .b(_T_1163)
    );
    wire _T_1165;
    BITWISEOR #(.width(1)) bitwiseor_4907 (
        .y(_T_1165),
        .a(_T_1164),
        .b(_divSqrt_in_flight__q)
    );
    wire _T_1167;
    EQ_UNSIGNED #(.width(1)) u_eq_4908 (
        .y(_T_1167),
        .a(_T_1165),
        .b(1'h0)
    );
    wire _T_1168;
    BITWISEOR #(.width(1)) bitwiseor_4909 (
        .y(_T_1168),
        .a(units_busy),
        .b(_write_port_busy__q)
    );
    wire _T_1169;
    BITWISEOR #(.width(1)) bitwiseor_4910 (
        .y(_T_1169),
        .a(_T_1168),
        .b(_divSqrt_in_flight__q)
    );
    wire _T_1171;
    EQ_UNSIGNED #(.width(1)) u_eq_4911 (
        .y(_T_1171),
        .a(_wb_cp_valid__q),
        .b(1'h0)
    );
    wire _T_1172;
    BITWISEAND #(.width(1)) bitwiseand_4912 (
        .y(_T_1172),
        .a(_wb_reg_valid__q),
        .b(_T_1171)
    );
    wire _T_1174;
    EQ_UNSIGNED #(.width(1)) u_eq_4913 (
        .y(_T_1174),
        .a(_mem_ctrl_single__q),
        .b(1'h0)
    );
    wire _T_1175;
    BITWISEAND #(.width(1)) bitwiseand_4914 (
        .y(_T_1175),
        .a(_mem_ctrl_fma__q),
        .b(_T_1174)
    );
    wire _T_1177;
    BITWISEOR #(.width(1)) bitwiseor_4915 (
        .y(_T_1177),
        .a(1'h0),
        .b(_T_1175)
    );
    wire _T_1178;
    BITWISEOR #(.width(1)) bitwiseor_4916 (
        .y(_T_1178),
        .a(_T_1177),
        .b(_mem_ctrl_div__q)
    );
    wire _T_1179;
    BITWISEOR #(.width(1)) bitwiseor_4917 (
        .y(_T_1179),
        .a(_T_1178),
        .b(_mem_ctrl_sqrt__q)
    );
    wire __T_1180__q;
    wire __T_1180__d;
    DFF_POSCLK #(.width(1)) _T_1180 (
        .q(__T_1180__q),
        .d(__T_1180__d),
        .clk(clock)
    );
    wire _T_1181;
    BITWISEAND #(.width(1)) bitwiseand_4918 (
        .y(_T_1181),
        .a(_T_1172),
        .b(__T_1180__q)
    );
    wire _T_1183;
    EQ_UNSIGNED #(.width(1)) u_eq_4919 (
        .y(_T_1183),
        .a(_wb_cp_valid__q),
        .b(1'h0)
    );
    wire _T_1184;
    BITS #(.width(3), .high(0), .low(0)) bits_4920 (
        .y(_T_1184),
        .in(_wen__q)
    );
    wire _T_1186;
    EQ_UNSIGNED #(.width(2)) u_eq_4921 (
        .y(_T_1186),
        .a(_wbInfo_0_pipeid__q),
        .b(2'h3)
    );
    wire _T_1188;
    BITWISEOR #(.width(1)) bitwiseor_4922 (
        .y(_T_1188),
        .a(1'h0),
        .b(_T_1186)
    );
    wire _T_1189;
    BITWISEAND #(.width(1)) bitwiseand_4923 (
        .y(_T_1189),
        .a(_T_1184),
        .b(_T_1188)
    );
    wire _T_1190;
    BITWISEOR #(.width(1)) bitwiseor_4924 (
        .y(_T_1190),
        .a(_divSqrt_wen__q),
        .b(_T_1189)
    );
    wire _T_1191;
    BITWISEAND #(.width(1)) bitwiseand_4925 (
        .y(_T_1191),
        .a(_T_1183),
        .b(_T_1190)
    );
    wire _T_1192;
    BITS #(.width(32), .high(14), .low(14)) bits_4926 (
        .y(_T_1192),
        .in(io_inst)
    );
    wire [1:0] _T_1193;
    BITS #(.width(32), .high(13), .low(12)) bits_4927 (
        .y(_T_1193),
        .in(io_inst)
    );
    wire _T_1195;
    LT_UNSIGNED #(.width(2)) u_lt_4928 (
        .y(_T_1195),
        .a(_T_1193),
        .b(2'h3)
    );
    wire _T_1197;
    GEQ_UNSIGNED #(.width(3)) u_geq_4929 (
        .y(_T_1197),
        .a(io_fcsr_rm),
        .b(3'h4)
    );
    wire _T_1198;
    BITWISEOR #(.width(1)) bitwiseor_4930 (
        .y(_T_1198),
        .a(_T_1195),
        .b(_T_1197)
    );
    wire _T_1199;
    BITWISEAND #(.width(1)) bitwiseand_4931 (
        .y(_T_1199),
        .a(_T_1192),
        .b(_T_1198)
    );
    wire [1:0] __T_1203__q;
    wire [1:0] __T_1203__d;
    DFF_POSCLK #(.width(2)) _T_1203 (
        .q(__T_1203__q),
        .d(__T_1203__d),
        .clk(clock)
    );
    wire [4:0] __T_1205__q;
    wire [4:0] __T_1205__d;
    DFF_POSCLK #(.width(5)) _T_1205 (
        .q(__T_1205__q),
        .d(__T_1205__d),
        .clk(clock)
    );
    wire [64:0] __T_1207__q;
    wire [64:0] __T_1207__d;
    DFF_POSCLK #(.width(65)) _T_1207 (
        .q(__T_1207__q),
        .d(__T_1207__d),
        .clk(clock)
    );
    wire _DivSqrtRecF64__clock;
    wire _DivSqrtRecF64__reset;
    wire _DivSqrtRecF64__io_inReady_div;
    wire _DivSqrtRecF64__io_inReady_sqrt;
    wire _DivSqrtRecF64__io_inValid;
    wire _DivSqrtRecF64__io_sqrtOp;
    wire [64:0] _DivSqrtRecF64__io_a;
    wire [64:0] _DivSqrtRecF64__io_b;
    wire [1:0] _DivSqrtRecF64__io_roundingMode;
    wire _DivSqrtRecF64__io_outValid_div;
    wire _DivSqrtRecF64__io_outValid_sqrt;
    wire [64:0] _DivSqrtRecF64__io_out;
    wire [4:0] _DivSqrtRecF64__io_exceptionFlags;
    DivSqrtRecF64 DivSqrtRecF64 (
        .clock(_DivSqrtRecF64__clock),
        .reset(_DivSqrtRecF64__reset),
        .io_inReady_div(_DivSqrtRecF64__io_inReady_div),
        .io_inReady_sqrt(_DivSqrtRecF64__io_inReady_sqrt),
        .io_inValid(_DivSqrtRecF64__io_inValid),
        .io_sqrtOp(_DivSqrtRecF64__io_sqrtOp),
        .io_a(_DivSqrtRecF64__io_a),
        .io_b(_DivSqrtRecF64__io_b),
        .io_roundingMode(_DivSqrtRecF64__io_roundingMode),
        .io_outValid_div(_DivSqrtRecF64__io_outValid_div),
        .io_outValid_sqrt(_DivSqrtRecF64__io_outValid_sqrt),
        .io_out(_DivSqrtRecF64__io_out),
        .io_exceptionFlags(_DivSqrtRecF64__io_exceptionFlags)
    );
    wire _T_1208;
    MUX_UNSIGNED #(.width(1)) u_mux_6280 (
        .y(_T_1208),
        .sel(_DivSqrtRecF64__io_sqrtOp),
        .a(_DivSqrtRecF64__io_inReady_sqrt),
        .b(_DivSqrtRecF64__io_inReady_div)
    );
    wire _T_1209;
    BITWISEOR #(.width(1)) bitwiseor_6281 (
        .y(_T_1209),
        .a(_DivSqrtRecF64__io_outValid_div),
        .b(_DivSqrtRecF64__io_outValid_sqrt)
    );
    wire _T_1210;
    BITWISEOR #(.width(1)) bitwiseor_6282 (
        .y(_T_1210),
        .a(_mem_ctrl_div__q),
        .b(_mem_ctrl_sqrt__q)
    );
    wire _T_1211;
    BITWISEAND #(.width(1)) bitwiseand_6283 (
        .y(_T_1211),
        .a(_mem_reg_valid__q),
        .b(_T_1210)
    );
    wire _T_1213;
    EQ_UNSIGNED #(.width(1)) u_eq_6284 (
        .y(_T_1213),
        .a(_divSqrt_in_flight__q),
        .b(1'h0)
    );
    wire _T_1214;
    BITWISEAND #(.width(1)) bitwiseand_6285 (
        .y(_T_1214),
        .a(_T_1211),
        .b(_T_1213)
    );
    wire _T_1215;
    BITWISEAND #(.width(1)) bitwiseand_6286 (
        .y(_T_1215),
        .a(_DivSqrtRecF64__io_inValid),
        .b(divSqrt_inReady)
    );
    wire [4:0] _T_1217;
    BITS #(.width(32), .high(11), .low(7)) bits_6287 (
        .y(_T_1217),
        .in(_mem_reg_inst__q)
    );
    wire _T_1219;
    EQ_UNSIGNED #(.width(1)) u_eq_6288 (
        .y(_T_1219),
        .a(_divSqrt_killed__q),
        .b(1'h0)
    );
    wire _node_73;
    MUX_UNSIGNED #(.width(1)) u_mux_6289 (
        .y(_node_73),
        .sel(_T_1215),
        .a(1'h1),
        .b(_divSqrt_in_flight__q)
    );
    wire _RecFNToRecFN__clock;
    wire _RecFNToRecFN__reset;
    wire [64:0] _RecFNToRecFN__io_in;
    wire [1:0] _RecFNToRecFN__io_roundingMode;
    wire [32:0] _RecFNToRecFN__io_out;
    wire [4:0] _RecFNToRecFN__io_exceptionFlags;
    RecFNToRecFN_2 RecFNToRecFN (
        .clock(_RecFNToRecFN__clock),
        .reset(_RecFNToRecFN__reset),
        .io_in(_RecFNToRecFN__io_in),
        .io_roundingMode(_RecFNToRecFN__io_roundingMode),
        .io_out(_RecFNToRecFN__io_out),
        .io_exceptionFlags(_RecFNToRecFN__io_exceptionFlags)
    );
    wire [64:0] _T_1221;
    wire [64:0] _WTEMP_921;
    PAD_UNSIGNED #(.width(33), .n(65)) u_pad_6530 (
        .y(_WTEMP_921),
        .in(_RecFNToRecFN__io_out)
    );
    MUX_UNSIGNED #(.width(65)) u_mux_6531 (
        .y(_T_1221),
        .sel(_divSqrt_single__q),
        .a(_WTEMP_921),
        .b(__T_1207__q)
    );
    wire [4:0] _T_1223;
    wire [4:0] _WTEMP_922;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_6532 (
        .y(_WTEMP_922),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(5)) u_mux_6533 (
        .y(_T_1223),
        .sel(_divSqrt_single__q),
        .a(_RecFNToRecFN__io_exceptionFlags),
        .b(_WTEMP_922)
    );
    wire [4:0] _T_1224;
    BITWISEOR #(.width(5)) bitwiseor_6534 (
        .y(_T_1224),
        .a(__T_1205__q),
        .b(_T_1223)
    );
    assign _DivSqrtRecF64__clock = clock;
    assign _DivSqrtRecF64__io_a = _fpiu__io_as_double_in1;
    assign _DivSqrtRecF64__io_b = _fpiu__io_as_double_in2;
    assign _DivSqrtRecF64__io_inValid = _T_1214;
    BITS #(.width(3), .high(1), .low(0)) bits_6535 (
        .y(_DivSqrtRecF64__io_roundingMode),
        .in(_fpiu__io_as_double_rm)
    );
    assign _DivSqrtRecF64__io_sqrtOp = _mem_ctrl_sqrt__q;
    assign _DivSqrtRecF64__reset = reset;
    assign _FPUFMAPipe__clock = clock;
    assign _FPUFMAPipe__io_in_bits_cmd = req_cmd;
    assign _FPUFMAPipe__io_in_bits_div = req_div;
    assign _FPUFMAPipe__io_in_bits_fastpipe = req_fastpipe;
    assign _FPUFMAPipe__io_in_bits_fma = req_fma;
    assign _FPUFMAPipe__io_in_bits_fromint = req_fromint;
    assign _FPUFMAPipe__io_in_bits_in1 = req_in1;
    assign _FPUFMAPipe__io_in_bits_in2 = req_in2;
    assign _FPUFMAPipe__io_in_bits_in3 = req_in3;
    assign _FPUFMAPipe__io_in_bits_ldst = req_ldst;
    assign _FPUFMAPipe__io_in_bits_ren1 = req_ren1;
    assign _FPUFMAPipe__io_in_bits_ren2 = req_ren2;
    assign _FPUFMAPipe__io_in_bits_ren3 = req_ren3;
    assign _FPUFMAPipe__io_in_bits_rm = req_rm;
    assign _FPUFMAPipe__io_in_bits_single = req_single;
    assign _FPUFMAPipe__io_in_bits_sqrt = req_sqrt;
    assign _FPUFMAPipe__io_in_bits_swap12 = req_swap12;
    assign _FPUFMAPipe__io_in_bits_swap23 = req_swap23;
    assign _FPUFMAPipe__io_in_bits_toint = req_toint;
    assign _FPUFMAPipe__io_in_bits_typ = req_typ;
    assign _FPUFMAPipe__io_in_bits_wen = req_wen;
    assign _FPUFMAPipe__io_in_bits_wflags = req_wflags;
    assign _FPUFMAPipe__io_in_valid = _T_886;
    assign _FPUFMAPipe__reset = reset;
    assign _RecFNToRecFN__clock = clock;
    assign _RecFNToRecFN__io_in = __T_1207__q;
    assign _RecFNToRecFN__io_roundingMode = __T_1203__q;
    assign _RecFNToRecFN__reset = reset;
    assign __T_1180__d = _T_1179;
    MUX_UNSIGNED #(.width(2)) u_mux_6536 (
        .y(__T_1203__d),
        .sel(_T_1215),
        .a(_DivSqrtRecF64__io_roundingMode),
        .b(__T_1203__q)
    );
    MUX_UNSIGNED #(.width(5)) u_mux_6537 (
        .y(__T_1205__d),
        .sel(_T_1209),
        .a(_DivSqrtRecF64__io_exceptionFlags),
        .b(__T_1205__q)
    );
    MUX_UNSIGNED #(.width(65)) u_mux_6538 (
        .y(__T_1207__d),
        .sel(_T_1209),
        .a(_DivSqrtRecF64__io_out),
        .b(__T_1207__q)
    );
    MUX_UNSIGNED #(.width(5)) u_mux_6539 (
        .y(__T_282_cmd__d),
        .sel(io_valid),
        .a(_fp_decoder__io_sigs_cmd),
        .b(__T_282_cmd__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6540 (
        .y(__T_282_div__d),
        .sel(io_valid),
        .a(_fp_decoder__io_sigs_div),
        .b(__T_282_div__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6541 (
        .y(__T_282_fastpipe__d),
        .sel(io_valid),
        .a(_fp_decoder__io_sigs_fastpipe),
        .b(__T_282_fastpipe__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6542 (
        .y(__T_282_fma__d),
        .sel(io_valid),
        .a(_fp_decoder__io_sigs_fma),
        .b(__T_282_fma__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6543 (
        .y(__T_282_fromint__d),
        .sel(io_valid),
        .a(_fp_decoder__io_sigs_fromint),
        .b(__T_282_fromint__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6544 (
        .y(__T_282_ldst__d),
        .sel(io_valid),
        .a(_fp_decoder__io_sigs_ldst),
        .b(__T_282_ldst__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6545 (
        .y(__T_282_ren1__d),
        .sel(io_valid),
        .a(_fp_decoder__io_sigs_ren1),
        .b(__T_282_ren1__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6546 (
        .y(__T_282_ren2__d),
        .sel(io_valid),
        .a(_fp_decoder__io_sigs_ren2),
        .b(__T_282_ren2__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6547 (
        .y(__T_282_ren3__d),
        .sel(io_valid),
        .a(_fp_decoder__io_sigs_ren3),
        .b(__T_282_ren3__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6548 (
        .y(__T_282_single__d),
        .sel(io_valid),
        .a(_fp_decoder__io_sigs_single),
        .b(__T_282_single__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6549 (
        .y(__T_282_sqrt__d),
        .sel(io_valid),
        .a(_fp_decoder__io_sigs_sqrt),
        .b(__T_282_sqrt__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6550 (
        .y(__T_282_swap12__d),
        .sel(io_valid),
        .a(_fp_decoder__io_sigs_swap12),
        .b(__T_282_swap12__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6551 (
        .y(__T_282_swap23__d),
        .sel(io_valid),
        .a(_fp_decoder__io_sigs_swap23),
        .b(__T_282_swap23__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6552 (
        .y(__T_282_toint__d),
        .sel(io_valid),
        .a(_fp_decoder__io_sigs_toint),
        .b(__T_282_toint__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6553 (
        .y(__T_282_wen__d),
        .sel(io_valid),
        .a(_fp_decoder__io_sigs_wen),
        .b(__T_282_wen__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6554 (
        .y(__T_282_wflags__d),
        .sel(io_valid),
        .a(_fp_decoder__io_sigs_wflags),
        .b(__T_282_wflags__q)
    );
    assign cp_ctrl_cmd = io_cp_req_bits_cmd;
    assign cp_ctrl_div = io_cp_req_bits_div;
    assign cp_ctrl_fastpipe = io_cp_req_bits_fastpipe;
    assign cp_ctrl_fma = io_cp_req_bits_fma;
    assign cp_ctrl_fromint = io_cp_req_bits_fromint;
    assign cp_ctrl_ldst = io_cp_req_bits_ldst;
    assign cp_ctrl_ren1 = io_cp_req_bits_ren1;
    assign cp_ctrl_ren2 = io_cp_req_bits_ren2;
    assign cp_ctrl_ren3 = io_cp_req_bits_ren3;
    assign cp_ctrl_single = io_cp_req_bits_single;
    assign cp_ctrl_sqrt = io_cp_req_bits_sqrt;
    assign cp_ctrl_swap12 = io_cp_req_bits_swap12;
    assign cp_ctrl_swap23 = io_cp_req_bits_swap23;
    assign cp_ctrl_toint = io_cp_req_bits_toint;
    assign cp_ctrl_wen = io_cp_req_bits_wen;
    assign cp_ctrl_wflags = io_cp_req_bits_wflags;
    assign divSqrt_flags = _T_1224;
    assign divSqrt_inReady = _T_1208;
    MUX_UNSIGNED #(.width(1)) u_mux_6555 (
        .y(_WTEMP_477),
        .sel(_T_1209),
        .a(1'h0),
        .b(_node_73)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6556 (
        .y(_divSqrt_killed__d),
        .sel(_T_1215),
        .a(killm),
        .b(_divSqrt_killed__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6557 (
        .y(_divSqrt_single__d),
        .sel(_T_1215),
        .a(_mem_ctrl_single__q),
        .b(_divSqrt_single__q)
    );
    MUX_UNSIGNED #(.width(5)) u_mux_6558 (
        .y(_divSqrt_waddr__d),
        .sel(_T_1215),
        .a(_T_1217),
        .b(_divSqrt_waddr__q)
    );
    assign divSqrt_wdata = _T_1221;
    MUX_UNSIGNED #(.width(1)) u_mux_6559 (
        .y(_divSqrt_wen__d),
        .sel(_T_1209),
        .a(_T_1219),
        .b(1'h0)
    );
    MUX_UNSIGNED #(.width(5)) u_mux_6560 (
        .y(_ex_ra1__d),
        .sel(io_valid),
        .a(_node_10),
        .b(_ex_ra1__q)
    );
    MUX_UNSIGNED #(.width(5)) u_mux_6561 (
        .y(_ex_ra2__d),
        .sel(io_valid),
        .a(_node_11),
        .b(_ex_ra2__q)
    );
    MUX_UNSIGNED #(.width(5)) u_mux_6562 (
        .y(_ex_ra3__d),
        .sel(io_valid),
        .a(_node_12),
        .b(_ex_ra3__q)
    );
    MUX_UNSIGNED #(.width(32)) u_mux_6563 (
        .y(_ex_reg_inst__d),
        .sel(io_valid),
        .a(io_inst),
        .b(_ex_reg_inst__q)
    );
    assign _WTEMP_0 = io_valid;
    assign _fp_decoder__clock = clock;
    assign _fp_decoder__io_inst = io_inst;
    assign _fp_decoder__reset = reset;
    assign _fpiu__clock = clock;
    assign _fpiu__io_in_bits_cmd = req_cmd;
    assign _fpiu__io_in_bits_div = req_div;
    assign _fpiu__io_in_bits_fastpipe = req_fastpipe;
    assign _fpiu__io_in_bits_fma = req_fma;
    assign _fpiu__io_in_bits_fromint = req_fromint;
    assign _fpiu__io_in_bits_in1 = req_in1;
    assign _fpiu__io_in_bits_in2 = req_in2;
    assign _fpiu__io_in_bits_in3 = req_in3;
    assign _fpiu__io_in_bits_ldst = req_ldst;
    assign _fpiu__io_in_bits_ren1 = req_ren1;
    assign _fpiu__io_in_bits_ren2 = req_ren2;
    assign _fpiu__io_in_bits_ren3 = req_ren3;
    assign _fpiu__io_in_bits_rm = req_rm;
    assign _fpiu__io_in_bits_single = req_single;
    assign _fpiu__io_in_bits_sqrt = req_sqrt;
    assign _fpiu__io_in_bits_swap12 = req_swap12;
    assign _fpiu__io_in_bits_swap23 = req_swap23;
    assign _fpiu__io_in_bits_toint = req_toint;
    assign _fpiu__io_in_bits_typ = req_typ;
    assign _fpiu__io_in_bits_wen = req_wen;
    assign _fpiu__io_in_bits_wflags = req_wflags;
    assign _fpiu__io_in_valid = _T_868;
    assign _fpiu__reset = reset;
    assign _fpmu__clock = clock;
    assign _fpmu__io_in_bits_cmd = req_cmd;
    assign _fpmu__io_in_bits_div = req_div;
    assign _fpmu__io_in_bits_fastpipe = req_fastpipe;
    assign _fpmu__io_in_bits_fma = req_fma;
    assign _fpmu__io_in_bits_fromint = req_fromint;
    assign _fpmu__io_in_bits_in1 = req_in1;
    assign _fpmu__io_in_bits_in2 = req_in2;
    assign _fpmu__io_in_bits_in3 = req_in3;
    assign _fpmu__io_in_bits_ldst = req_ldst;
    assign _fpmu__io_in_bits_ren1 = req_ren1;
    assign _fpmu__io_in_bits_ren2 = req_ren2;
    assign _fpmu__io_in_bits_ren3 = req_ren3;
    assign _fpmu__io_in_bits_rm = req_rm;
    assign _fpmu__io_in_bits_single = req_single;
    assign _fpmu__io_in_bits_sqrt = req_sqrt;
    assign _fpmu__io_in_bits_swap12 = req_swap12;
    assign _fpmu__io_in_bits_swap23 = req_swap23;
    assign _fpmu__io_in_bits_toint = req_toint;
    assign _fpmu__io_in_bits_typ = req_typ;
    assign _fpmu__io_in_bits_wen = req_wen;
    assign _fpmu__io_in_bits_wflags = req_wflags;
    assign _fpmu__io_in_valid = _T_874;
    assign _fpmu__io_lt = _fpiu__io_out_bits_lt;
    assign _fpmu__reset = reset;
    assign _ifpu__clock = clock;
    assign _ifpu__io_in_bits_cmd = req_cmd;
    assign _ifpu__io_in_bits_div = req_div;
    assign _ifpu__io_in_bits_fastpipe = req_fastpipe;
    assign _ifpu__io_in_bits_fma = req_fma;
    assign _ifpu__io_in_bits_fromint = req_fromint;
    assign _ifpu__io_in_bits_in1 = _T_873;
    assign _ifpu__io_in_bits_in2 = req_in2;
    assign _ifpu__io_in_bits_in3 = req_in3;
    assign _ifpu__io_in_bits_ldst = req_ldst;
    assign _ifpu__io_in_bits_ren1 = req_ren1;
    assign _ifpu__io_in_bits_ren2 = req_ren2;
    assign _ifpu__io_in_bits_ren3 = req_ren3;
    assign _ifpu__io_in_bits_rm = req_rm;
    assign _ifpu__io_in_bits_single = req_single;
    assign _ifpu__io_in_bits_sqrt = req_sqrt;
    assign _ifpu__io_in_bits_swap12 = req_swap12;
    assign _ifpu__io_in_bits_swap23 = req_swap23;
    assign _ifpu__io_in_bits_toint = req_toint;
    assign _ifpu__io_in_bits_typ = req_typ;
    assign _ifpu__io_in_bits_wen = req_wen;
    assign _ifpu__io_in_bits_wflags = req_wflags;
    assign _ifpu__io_in_valid = _T_872;
    assign _ifpu__reset = reset;
    assign io_cp_req_ready = _T_1136;
    wire [64:0] _WTEMP_923;
    PAD_UNSIGNED #(.width(64), .n(65)) u_pad_6564 (
        .y(_WTEMP_923),
        .in(_node_69)
    );
    MUX_UNSIGNED #(.width(65)) u_mux_6565 (
        .y(io_cp_resp_bits_data),
        .sel(_T_1133),
        .a(wdata),
        .b(_WTEMP_923)
    );
    assign io_cp_resp_bits_exc = 5'h0;
    MUX_UNSIGNED #(.width(1)) u_mux_6566 (
        .y(io_cp_resp_valid),
        .sel(_T_1133),
        .a(1'h1),
        .b(_node_70)
    );
    assign io_dec_cmd = _fp_decoder__io_sigs_cmd;
    assign io_dec_div = _fp_decoder__io_sigs_div;
    assign io_dec_fastpipe = _fp_decoder__io_sigs_fastpipe;
    assign io_dec_fma = _fp_decoder__io_sigs_fma;
    assign io_dec_fromint = _fp_decoder__io_sigs_fromint;
    assign io_dec_ldst = _fp_decoder__io_sigs_ldst;
    assign io_dec_ren1 = _fp_decoder__io_sigs_ren1;
    assign io_dec_ren2 = _fp_decoder__io_sigs_ren2;
    assign io_dec_ren3 = _fp_decoder__io_sigs_ren3;
    assign io_dec_single = _fp_decoder__io_sigs_single;
    assign io_dec_sqrt = _fp_decoder__io_sigs_sqrt;
    assign io_dec_swap12 = _fp_decoder__io_sigs_swap12;
    assign io_dec_swap23 = _fp_decoder__io_sigs_swap23;
    assign io_dec_toint = _fp_decoder__io_sigs_toint;
    assign io_dec_wen = _fp_decoder__io_sigs_wen;
    assign io_dec_wflags = _fp_decoder__io_sigs_wflags;
    assign io_fcsr_flags_bits = _T_1149;
    assign io_fcsr_flags_valid = _T_1140;
    assign io_fcsr_rdy = _T_1167;
    assign io_illegal_rm = _T_1199;
    assign io_nack_mem = _T_1169;
    assign io_sboard_clr = _T_1191;
    assign io_sboard_clra = waddr;
    assign io_sboard_set = _T_1181;
    assign io_store_data = _fpiu__io_out_bits_store;
    assign io_toint_data = _fpiu__io_out_bits_toint;
    assign _load_wb__d = io_dmem_resp_val;
    MUX_UNSIGNED #(.width(64)) u_mux_6567 (
        .y(_load_wb_data__d),
        .sel(io_dmem_resp_val),
        .a(io_dmem_resp_data),
        .b(_load_wb_data__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6568 (
        .y(_load_wb_single__d),
        .sel(io_dmem_resp_val),
        .a(_T_383),
        .b(_load_wb_single__q)
    );
    MUX_UNSIGNED #(.width(5)) u_mux_6569 (
        .y(_load_wb_tag__d),
        .sel(io_dmem_resp_val),
        .a(io_dmem_resp_tag),
        .b(_load_wb_tag__q)
    );
    assign _WTEMP_2 = ex_cp_valid;
    MUX_UNSIGNED #(.width(5)) u_mux_6570 (
        .y(_mem_ctrl_cmd__d),
        .sel(req_valid),
        .a(ex_ctrl_cmd),
        .b(_mem_ctrl_cmd__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6571 (
        .y(_mem_ctrl_div__d),
        .sel(req_valid),
        .a(ex_ctrl_div),
        .b(_mem_ctrl_div__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6572 (
        .y(_mem_ctrl_fastpipe__d),
        .sel(req_valid),
        .a(ex_ctrl_fastpipe),
        .b(_mem_ctrl_fastpipe__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6573 (
        .y(_mem_ctrl_fma__d),
        .sel(req_valid),
        .a(ex_ctrl_fma),
        .b(_mem_ctrl_fma__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6574 (
        .y(_mem_ctrl_fromint__d),
        .sel(req_valid),
        .a(ex_ctrl_fromint),
        .b(_mem_ctrl_fromint__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6575 (
        .y(_mem_ctrl_ldst__d),
        .sel(req_valid),
        .a(ex_ctrl_ldst),
        .b(_mem_ctrl_ldst__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6576 (
        .y(_mem_ctrl_ren1__d),
        .sel(req_valid),
        .a(ex_ctrl_ren1),
        .b(_mem_ctrl_ren1__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6577 (
        .y(_mem_ctrl_ren2__d),
        .sel(req_valid),
        .a(ex_ctrl_ren2),
        .b(_mem_ctrl_ren2__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6578 (
        .y(_mem_ctrl_ren3__d),
        .sel(req_valid),
        .a(ex_ctrl_ren3),
        .b(_mem_ctrl_ren3__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6579 (
        .y(_mem_ctrl_single__d),
        .sel(req_valid),
        .a(ex_ctrl_single),
        .b(_mem_ctrl_single__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6580 (
        .y(_mem_ctrl_sqrt__d),
        .sel(req_valid),
        .a(ex_ctrl_sqrt),
        .b(_mem_ctrl_sqrt__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6581 (
        .y(_mem_ctrl_swap12__d),
        .sel(req_valid),
        .a(ex_ctrl_swap12),
        .b(_mem_ctrl_swap12__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6582 (
        .y(_mem_ctrl_swap23__d),
        .sel(req_valid),
        .a(ex_ctrl_swap23),
        .b(_mem_ctrl_swap23__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6583 (
        .y(_mem_ctrl_toint__d),
        .sel(req_valid),
        .a(ex_ctrl_toint),
        .b(_mem_ctrl_toint__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6584 (
        .y(_mem_ctrl_wen__d),
        .sel(req_valid),
        .a(ex_ctrl_wen),
        .b(_mem_ctrl_wen__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6585 (
        .y(_mem_ctrl_wflags__d),
        .sel(req_valid),
        .a(ex_ctrl_wflags),
        .b(_mem_ctrl_wflags__q)
    );
    MUX_UNSIGNED #(.width(32)) u_mux_6586 (
        .y(_mem_reg_inst__d),
        .sel(_ex_reg_valid__q),
        .a(_ex_reg_inst__q),
        .b(_mem_reg_inst__q)
    );
    assign _WTEMP_1 = _T_217;
    assign regfile__T_1131_data = wdata;
    assign regfile__T_782_data = load_wb_data_recoded;
    MUX_UNSIGNED #(.width(5)) u_mux_6587 (
        .y(req_cmd),
        .sel(ex_cp_valid),
        .a(io_cp_req_bits_cmd),
        .b(ex_ctrl_cmd)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6588 (
        .y(req_div),
        .sel(ex_cp_valid),
        .a(io_cp_req_bits_div),
        .b(ex_ctrl_div)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6589 (
        .y(req_fastpipe),
        .sel(ex_cp_valid),
        .a(io_cp_req_bits_fastpipe),
        .b(ex_ctrl_fastpipe)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6590 (
        .y(req_fma),
        .sel(ex_cp_valid),
        .a(io_cp_req_bits_fma),
        .b(ex_ctrl_fma)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6591 (
        .y(req_fromint),
        .sel(ex_cp_valid),
        .a(io_cp_req_bits_fromint),
        .b(ex_ctrl_fromint)
    );
    MUX_UNSIGNED #(.width(65)) u_mux_6592 (
        .y(req_in1),
        .sel(ex_cp_valid),
        .a(io_cp_req_bits_in1),
        .b(regfile__T_849_data)
    );
    MUX_UNSIGNED #(.width(65)) u_mux_6593 (
        .y(req_in2),
        .sel(ex_cp_valid),
        .a(_node_13),
        .b(regfile__T_853_data)
    );
    MUX_UNSIGNED #(.width(65)) u_mux_6594 (
        .y(req_in3),
        .sel(ex_cp_valid),
        .a(_node_14),
        .b(regfile__T_857_data)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6595 (
        .y(req_ldst),
        .sel(ex_cp_valid),
        .a(io_cp_req_bits_ldst),
        .b(ex_ctrl_ldst)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6596 (
        .y(req_ren1),
        .sel(ex_cp_valid),
        .a(io_cp_req_bits_ren1),
        .b(ex_ctrl_ren1)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6597 (
        .y(req_ren2),
        .sel(ex_cp_valid),
        .a(io_cp_req_bits_ren2),
        .b(ex_ctrl_ren2)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6598 (
        .y(req_ren3),
        .sel(ex_cp_valid),
        .a(io_cp_req_bits_ren3),
        .b(ex_ctrl_ren3)
    );
    MUX_UNSIGNED #(.width(3)) u_mux_6599 (
        .y(req_rm),
        .sel(ex_cp_valid),
        .a(io_cp_req_bits_rm),
        .b(ex_rm)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6600 (
        .y(req_single),
        .sel(ex_cp_valid),
        .a(io_cp_req_bits_single),
        .b(ex_ctrl_single)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6601 (
        .y(req_sqrt),
        .sel(ex_cp_valid),
        .a(io_cp_req_bits_sqrt),
        .b(ex_ctrl_sqrt)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6602 (
        .y(req_swap12),
        .sel(ex_cp_valid),
        .a(io_cp_req_bits_swap12),
        .b(ex_ctrl_swap12)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6603 (
        .y(req_swap23),
        .sel(ex_cp_valid),
        .a(io_cp_req_bits_swap23),
        .b(ex_ctrl_swap23)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6604 (
        .y(req_toint),
        .sel(ex_cp_valid),
        .a(io_cp_req_bits_toint),
        .b(ex_ctrl_toint)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_6605 (
        .y(req_typ),
        .sel(ex_cp_valid),
        .a(io_cp_req_bits_typ),
        .b(_T_858)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6606 (
        .y(req_wen),
        .sel(ex_cp_valid),
        .a(io_cp_req_bits_wen),
        .b(ex_ctrl_wen)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6607 (
        .y(req_wflags),
        .sel(ex_cp_valid),
        .a(io_cp_req_bits_wflags),
        .b(ex_ctrl_wflags)
    );
    assign _sfma__clock = clock;
    assign _sfma__io_in_bits_cmd = req_cmd;
    assign _sfma__io_in_bits_div = req_div;
    assign _sfma__io_in_bits_fastpipe = req_fastpipe;
    assign _sfma__io_in_bits_fma = req_fma;
    assign _sfma__io_in_bits_fromint = req_fromint;
    assign _sfma__io_in_bits_in1 = req_in1;
    assign _sfma__io_in_bits_in2 = req_in2;
    assign _sfma__io_in_bits_in3 = req_in3;
    assign _sfma__io_in_bits_ldst = req_ldst;
    assign _sfma__io_in_bits_ren1 = req_ren1;
    assign _sfma__io_in_bits_ren2 = req_ren2;
    assign _sfma__io_in_bits_ren3 = req_ren3;
    assign _sfma__io_in_bits_rm = req_rm;
    assign _sfma__io_in_bits_single = req_single;
    assign _sfma__io_in_bits_sqrt = req_sqrt;
    assign _sfma__io_in_bits_swap12 = req_swap12;
    assign _sfma__io_in_bits_swap23 = req_swap23;
    assign _sfma__io_in_bits_toint = req_toint;
    assign _sfma__io_in_bits_typ = req_typ;
    assign _sfma__io_in_bits_wen = req_wen;
    assign _sfma__io_in_bits_wflags = req_wflags;
    assign _sfma__io_in_valid = _T_860;
    assign _sfma__reset = reset;
    MUX_UNSIGNED #(.width(1)) u_mux_6608 (
        .y(_wbInfo_0_cp__d),
        .sel(mem_wen),
        .a(_node_48),
        .b(_node_49)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_6609 (
        .y(_wbInfo_0_pipeid__d),
        .sel(mem_wen),
        .a(_node_50),
        .b(_node_51)
    );
    MUX_UNSIGNED #(.width(5)) u_mux_6610 (
        .y(_wbInfo_0_rd__d),
        .sel(mem_wen),
        .a(_node_52),
        .b(_node_53)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6611 (
        .y(_wbInfo_0_single__d),
        .sel(mem_wen),
        .a(_node_54),
        .b(_node_55)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6612 (
        .y(_wbInfo_1_cp__d),
        .sel(mem_wen),
        .a(_node_56),
        .b(_node_57)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_6613 (
        .y(_wbInfo_1_pipeid__d),
        .sel(mem_wen),
        .a(_node_58),
        .b(_node_59)
    );
    MUX_UNSIGNED #(.width(5)) u_mux_6614 (
        .y(_wbInfo_1_rd__d),
        .sel(mem_wen),
        .a(_node_60),
        .b(_node_61)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6615 (
        .y(_wbInfo_1_single__d),
        .sel(mem_wen),
        .a(_node_62),
        .b(_node_63)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6616 (
        .y(_wbInfo_2_cp__d),
        .sel(mem_wen),
        .a(_node_64),
        .b(_wbInfo_2_cp__q)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_6617 (
        .y(_wbInfo_2_pipeid__d),
        .sel(mem_wen),
        .a(_node_65),
        .b(_wbInfo_2_pipeid__q)
    );
    MUX_UNSIGNED #(.width(5)) u_mux_6618 (
        .y(_wbInfo_2_rd__d),
        .sel(mem_wen),
        .a(_node_66),
        .b(_wbInfo_2_rd__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6619 (
        .y(_wbInfo_2_single__d),
        .sel(mem_wen),
        .a(_node_67),
        .b(_wbInfo_2_single__q)
    );
    assign _WTEMP_4 = _mem_cp_valid__q;
    MUX_UNSIGNED #(.width(5)) u_mux_6620 (
        .y(_wb_ctrl_cmd__d),
        .sel(_mem_reg_valid__q),
        .a(_mem_ctrl_cmd__q),
        .b(_wb_ctrl_cmd__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6621 (
        .y(_wb_ctrl_div__d),
        .sel(_mem_reg_valid__q),
        .a(_mem_ctrl_div__q),
        .b(_wb_ctrl_div__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6622 (
        .y(_wb_ctrl_fastpipe__d),
        .sel(_mem_reg_valid__q),
        .a(_mem_ctrl_fastpipe__q),
        .b(_wb_ctrl_fastpipe__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6623 (
        .y(_wb_ctrl_fma__d),
        .sel(_mem_reg_valid__q),
        .a(_mem_ctrl_fma__q),
        .b(_wb_ctrl_fma__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6624 (
        .y(_wb_ctrl_fromint__d),
        .sel(_mem_reg_valid__q),
        .a(_mem_ctrl_fromint__q),
        .b(_wb_ctrl_fromint__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6625 (
        .y(_wb_ctrl_ldst__d),
        .sel(_mem_reg_valid__q),
        .a(_mem_ctrl_ldst__q),
        .b(_wb_ctrl_ldst__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6626 (
        .y(_wb_ctrl_ren1__d),
        .sel(_mem_reg_valid__q),
        .a(_mem_ctrl_ren1__q),
        .b(_wb_ctrl_ren1__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6627 (
        .y(_wb_ctrl_ren2__d),
        .sel(_mem_reg_valid__q),
        .a(_mem_ctrl_ren2__q),
        .b(_wb_ctrl_ren2__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6628 (
        .y(_wb_ctrl_ren3__d),
        .sel(_mem_reg_valid__q),
        .a(_mem_ctrl_ren3__q),
        .b(_wb_ctrl_ren3__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6629 (
        .y(_wb_ctrl_single__d),
        .sel(_mem_reg_valid__q),
        .a(_mem_ctrl_single__q),
        .b(_wb_ctrl_single__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6630 (
        .y(_wb_ctrl_sqrt__d),
        .sel(_mem_reg_valid__q),
        .a(_mem_ctrl_sqrt__q),
        .b(_wb_ctrl_sqrt__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6631 (
        .y(_wb_ctrl_swap12__d),
        .sel(_mem_reg_valid__q),
        .a(_mem_ctrl_swap12__q),
        .b(_wb_ctrl_swap12__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6632 (
        .y(_wb_ctrl_swap23__d),
        .sel(_mem_reg_valid__q),
        .a(_mem_ctrl_swap23__q),
        .b(_wb_ctrl_swap23__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6633 (
        .y(_wb_ctrl_toint__d),
        .sel(_mem_reg_valid__q),
        .a(_mem_ctrl_toint__q),
        .b(_wb_ctrl_toint__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6634 (
        .y(_wb_ctrl_wen__d),
        .sel(_mem_reg_valid__q),
        .a(_mem_ctrl_wen__q),
        .b(_wb_ctrl_wen__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6635 (
        .y(_wb_ctrl_wflags__d),
        .sel(_mem_reg_valid__q),
        .a(_mem_ctrl_wflags__q),
        .b(_wb_ctrl_wflags__q)
    );
    assign _WTEMP_3 = _T_227;
    MUX_UNSIGNED #(.width(5)) u_mux_6636 (
        .y(_wb_toint_exc__d),
        .sel(_mem_ctrl_toint__q),
        .a(_fpiu__io_out_bits_exc),
        .b(_wb_toint_exc__q)
    );
    wire [2:0] _WTEMP_924;
    PAD_UNSIGNED #(.width(2), .n(3)) u_pad_6637 (
        .y(_WTEMP_924),
        .in(_T_1017)
    );
    MUX_UNSIGNED #(.width(3)) u_mux_6638 (
        .y(_WTEMP_650),
        .sel(mem_wen),
        .a(_node_68),
        .b(_WTEMP_924)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6639 (
        .y(_write_port_busy__d),
        .sel(req_valid),
        .a(_T_1013),
        .b(_write_port_busy__q)
    );
endmodule //FPU
module DFF_POSCLK(q, d, clk);
    parameter width = 4;
    output reg [width-1:0] q;
    input [width-1:0] d;
    input clk;
    always @(posedge clk) begin
        q <= d;
    end
endmodule // DFF_POSCLK
module MUX_UNSIGNED(y, sel, a, b);
    parameter width = 4;
    output [width-1:0] y;
    input sel;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = sel ? a : b;
endmodule // MUX_UNSIGNED
module BITWISEOR(y, a, b);
    parameter width = 4;
    output [width-1:0] y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a | b;
endmodule // BITWISEOR
module BITWISEAND(y, a, b);
    parameter width = 4;
    output [width-1:0] y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a & b;
endmodule // BITWISEAND
module EQ_UNSIGNED(y, a, b);
    parameter width = 4;
    output y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a == b;
endmodule // EQ_UNSIGNED
module FPUDecoder(
    input clock,
    input reset,
    input [31:0] io_inst,
    output [4:0] io_sigs_cmd,
    output io_sigs_ldst,
    output io_sigs_wen,
    output io_sigs_ren1,
    output io_sigs_ren2,
    output io_sigs_ren3,
    output io_sigs_swap12,
    output io_sigs_swap23,
    output io_sigs_single,
    output io_sigs_fromint,
    output io_sigs_toint,
    output io_sigs_fastpipe,
    output io_sigs_fma,
    output io_sigs_div,
    output io_sigs_sqrt,
    output io_sigs_wflags
);
    wire [31:0] _T_22;
    BITWISEAND #(.width(32)) bitwiseand_17 (
        .y(_T_22),
        .a(io_inst),
        .b(32'h4)
    );
    wire _T_24;
    EQ_UNSIGNED #(.width(32)) u_eq_18 (
        .y(_T_24),
        .a(_T_22),
        .b(32'h4)
    );
    wire [31:0] _T_26;
    BITWISEAND #(.width(32)) bitwiseand_19 (
        .y(_T_26),
        .a(io_inst),
        .b(32'h8000010)
    );
    wire _T_28;
    EQ_UNSIGNED #(.width(32)) u_eq_20 (
        .y(_T_28),
        .a(_T_26),
        .b(32'h8000010)
    );
    wire _T_30;
    BITWISEOR #(.width(1)) bitwiseor_21 (
        .y(_T_30),
        .a(1'h0),
        .b(_T_24)
    );
    wire _T_31;
    BITWISEOR #(.width(1)) bitwiseor_22 (
        .y(_T_31),
        .a(_T_30),
        .b(_T_28)
    );
    wire [31:0] _T_33;
    BITWISEAND #(.width(32)) bitwiseand_23 (
        .y(_T_33),
        .a(io_inst),
        .b(32'h8)
    );
    wire _T_35;
    EQ_UNSIGNED #(.width(32)) u_eq_24 (
        .y(_T_35),
        .a(_T_33),
        .b(32'h8)
    );
    wire [31:0] _T_37;
    BITWISEAND #(.width(32)) bitwiseand_25 (
        .y(_T_37),
        .a(io_inst),
        .b(32'h10000010)
    );
    wire _T_39;
    EQ_UNSIGNED #(.width(32)) u_eq_26 (
        .y(_T_39),
        .a(_T_37),
        .b(32'h10000010)
    );
    wire _T_41;
    BITWISEOR #(.width(1)) bitwiseor_27 (
        .y(_T_41),
        .a(1'h0),
        .b(_T_35)
    );
    wire _T_42;
    BITWISEOR #(.width(1)) bitwiseor_28 (
        .y(_T_42),
        .a(_T_41),
        .b(_T_39)
    );
    wire [31:0] _T_44;
    BITWISEAND #(.width(32)) bitwiseand_29 (
        .y(_T_44),
        .a(io_inst),
        .b(32'h40)
    );
    wire _T_46;
    EQ_UNSIGNED #(.width(32)) u_eq_30 (
        .y(_T_46),
        .a(_T_44),
        .b(32'h0)
    );
    wire [31:0] _T_48;
    BITWISEAND #(.width(32)) bitwiseand_31 (
        .y(_T_48),
        .a(io_inst),
        .b(32'h20000000)
    );
    wire _T_50;
    EQ_UNSIGNED #(.width(32)) u_eq_32 (
        .y(_T_50),
        .a(_T_48),
        .b(32'h20000000)
    );
    wire _T_52;
    BITWISEOR #(.width(1)) bitwiseor_33 (
        .y(_T_52),
        .a(1'h0),
        .b(_T_46)
    );
    wire _T_53;
    BITWISEOR #(.width(1)) bitwiseor_34 (
        .y(_T_53),
        .a(_T_52),
        .b(_T_50)
    );
    wire [31:0] _T_55;
    BITWISEAND #(.width(32)) bitwiseand_35 (
        .y(_T_55),
        .a(io_inst),
        .b(32'h40000000)
    );
    wire _T_57;
    EQ_UNSIGNED #(.width(32)) u_eq_36 (
        .y(_T_57),
        .a(_T_55),
        .b(32'h40000000)
    );
    wire _T_59;
    BITWISEOR #(.width(1)) bitwiseor_37 (
        .y(_T_59),
        .a(1'h0),
        .b(_T_46)
    );
    wire _T_60;
    BITWISEOR #(.width(1)) bitwiseor_38 (
        .y(_T_60),
        .a(_T_59),
        .b(_T_57)
    );
    wire [31:0] _T_62;
    BITWISEAND #(.width(32)) bitwiseand_39 (
        .y(_T_62),
        .a(io_inst),
        .b(32'h10)
    );
    wire _T_64;
    EQ_UNSIGNED #(.width(32)) u_eq_40 (
        .y(_T_64),
        .a(_T_62),
        .b(32'h0)
    );
    wire _T_66;
    BITWISEOR #(.width(1)) bitwiseor_41 (
        .y(_T_66),
        .a(1'h0),
        .b(_T_64)
    );
    wire [1:0] _T_67;
    CAT #(.width_a(1), .width_b(1)) cat_42 (
        .y(_T_67),
        .a(_T_42),
        .b(_T_31)
    );
    wire [1:0] _T_68;
    CAT #(.width_a(1), .width_b(1)) cat_43 (
        .y(_T_68),
        .a(_T_66),
        .b(_T_60)
    );
    wire [2:0] _T_69;
    CAT #(.width_a(2), .width_b(1)) cat_44 (
        .y(_T_69),
        .a(_T_68),
        .b(_T_53)
    );
    wire [4:0] decoder_0;
    CAT #(.width_a(3), .width_b(2)) cat_45 (
        .y(decoder_0),
        .a(_T_69),
        .b(_T_67)
    );
    wire decoder_1;
    BITWISEOR #(.width(1)) bitwiseor_46 (
        .y(decoder_1),
        .a(1'h0),
        .b(_T_46)
    );
    wire [31:0] _T_72;
    BITWISEAND #(.width(32)) bitwiseand_47 (
        .y(_T_72),
        .a(io_inst),
        .b(32'h80000020)
    );
    wire _T_74;
    EQ_UNSIGNED #(.width(32)) u_eq_48 (
        .y(_T_74),
        .a(_T_72),
        .b(32'h0)
    );
    wire [31:0] _T_76;
    BITWISEAND #(.width(32)) bitwiseand_49 (
        .y(_T_76),
        .a(io_inst),
        .b(32'h30)
    );
    wire _T_78;
    EQ_UNSIGNED #(.width(32)) u_eq_50 (
        .y(_T_78),
        .a(_T_76),
        .b(32'h0)
    );
    wire [31:0] _T_80;
    BITWISEAND #(.width(32)) bitwiseand_51 (
        .y(_T_80),
        .a(io_inst),
        .b(32'h10000020)
    );
    wire _T_82;
    EQ_UNSIGNED #(.width(32)) u_eq_52 (
        .y(_T_82),
        .a(_T_80),
        .b(32'h10000000)
    );
    wire _T_84;
    BITWISEOR #(.width(1)) bitwiseor_53 (
        .y(_T_84),
        .a(1'h0),
        .b(_T_74)
    );
    wire _T_85;
    BITWISEOR #(.width(1)) bitwiseor_54 (
        .y(_T_85),
        .a(_T_84),
        .b(_T_78)
    );
    wire decoder_2;
    BITWISEOR #(.width(1)) bitwiseor_55 (
        .y(decoder_2),
        .a(_T_85),
        .b(_T_82)
    );
    wire [31:0] _T_87;
    BITWISEAND #(.width(32)) bitwiseand_56 (
        .y(_T_87),
        .a(io_inst),
        .b(32'h80000004)
    );
    wire _T_89;
    EQ_UNSIGNED #(.width(32)) u_eq_57 (
        .y(_T_89),
        .a(_T_87),
        .b(32'h0)
    );
    wire [31:0] _T_91;
    BITWISEAND #(.width(32)) bitwiseand_58 (
        .y(_T_91),
        .a(io_inst),
        .b(32'h10000004)
    );
    wire _T_93;
    EQ_UNSIGNED #(.width(32)) u_eq_59 (
        .y(_T_93),
        .a(_T_91),
        .b(32'h0)
    );
    wire [31:0] _T_95;
    BITWISEAND #(.width(32)) bitwiseand_60 (
        .y(_T_95),
        .a(io_inst),
        .b(32'h50)
    );
    wire _T_97;
    EQ_UNSIGNED #(.width(32)) u_eq_61 (
        .y(_T_97),
        .a(_T_95),
        .b(32'h40)
    );
    wire _T_99;
    BITWISEOR #(.width(1)) bitwiseor_62 (
        .y(_T_99),
        .a(1'h0),
        .b(_T_89)
    );
    wire _T_100;
    BITWISEOR #(.width(1)) bitwiseor_63 (
        .y(_T_100),
        .a(_T_99),
        .b(_T_93)
    );
    wire decoder_3;
    BITWISEOR #(.width(1)) bitwiseor_64 (
        .y(decoder_3),
        .a(_T_100),
        .b(_T_97)
    );
    wire [31:0] _T_102;
    BITWISEAND #(.width(32)) bitwiseand_65 (
        .y(_T_102),
        .a(io_inst),
        .b(32'h40000004)
    );
    wire _T_104;
    EQ_UNSIGNED #(.width(32)) u_eq_66 (
        .y(_T_104),
        .a(_T_102),
        .b(32'h0)
    );
    wire [31:0] _T_106;
    BITWISEAND #(.width(32)) bitwiseand_67 (
        .y(_T_106),
        .a(io_inst),
        .b(32'h20)
    );
    wire _T_108;
    EQ_UNSIGNED #(.width(32)) u_eq_68 (
        .y(_T_108),
        .a(_T_106),
        .b(32'h20)
    );
    wire _T_110;
    BITWISEOR #(.width(1)) bitwiseor_69 (
        .y(_T_110),
        .a(1'h0),
        .b(_T_104)
    );
    wire _T_111;
    BITWISEOR #(.width(1)) bitwiseor_70 (
        .y(_T_111),
        .a(_T_110),
        .b(_T_108)
    );
    wire decoder_4;
    BITWISEOR #(.width(1)) bitwiseor_71 (
        .y(decoder_4),
        .a(_T_111),
        .b(_T_97)
    );
    wire decoder_5;
    BITWISEOR #(.width(1)) bitwiseor_72 (
        .y(decoder_5),
        .a(1'h0),
        .b(_T_97)
    );
    wire [31:0] _T_114;
    BITWISEAND #(.width(32)) bitwiseand_73 (
        .y(_T_114),
        .a(io_inst),
        .b(32'h50000010)
    );
    wire _T_116;
    EQ_UNSIGNED #(.width(32)) u_eq_74 (
        .y(_T_116),
        .a(_T_114),
        .b(32'h50000010)
    );
    wire _T_118;
    BITWISEOR #(.width(1)) bitwiseor_75 (
        .y(_T_118),
        .a(1'h0),
        .b(_T_46)
    );
    wire decoder_6;
    BITWISEOR #(.width(1)) bitwiseor_76 (
        .y(decoder_6),
        .a(_T_118),
        .b(_T_116)
    );
    wire [31:0] _T_120;
    BITWISEAND #(.width(32)) bitwiseand_77 (
        .y(_T_120),
        .a(io_inst),
        .b(32'h30000010)
    );
    wire _T_122;
    EQ_UNSIGNED #(.width(32)) u_eq_78 (
        .y(_T_122),
        .a(_T_120),
        .b(32'h10)
    );
    wire decoder_7;
    BITWISEOR #(.width(1)) bitwiseor_79 (
        .y(decoder_7),
        .a(1'h0),
        .b(_T_122)
    );
    wire [31:0] _T_125;
    BITWISEAND #(.width(32)) bitwiseand_80 (
        .y(_T_125),
        .a(io_inst),
        .b(32'h1040)
    );
    wire _T_127;
    EQ_UNSIGNED #(.width(32)) u_eq_81 (
        .y(_T_127),
        .a(_T_125),
        .b(32'h0)
    );
    wire [31:0] _T_129;
    BITWISEAND #(.width(32)) bitwiseand_82 (
        .y(_T_129),
        .a(io_inst),
        .b(32'h2000040)
    );
    wire _T_131;
    EQ_UNSIGNED #(.width(32)) u_eq_83 (
        .y(_T_131),
        .a(_T_129),
        .b(32'h40)
    );
    wire _T_133;
    BITWISEOR #(.width(1)) bitwiseor_84 (
        .y(_T_133),
        .a(1'h0),
        .b(_T_127)
    );
    wire decoder_8;
    BITWISEOR #(.width(1)) bitwiseor_85 (
        .y(decoder_8),
        .a(_T_133),
        .b(_T_131)
    );
    wire [31:0] _T_135;
    BITWISEAND #(.width(32)) bitwiseand_86 (
        .y(_T_135),
        .a(io_inst),
        .b(32'h90000010)
    );
    wire _T_137;
    EQ_UNSIGNED #(.width(32)) u_eq_87 (
        .y(_T_137),
        .a(_T_135),
        .b(32'h90000010)
    );
    wire decoder_9;
    BITWISEOR #(.width(1)) bitwiseor_88 (
        .y(decoder_9),
        .a(1'h0),
        .b(_T_137)
    );
    wire [31:0] _T_140;
    BITWISEAND #(.width(32)) bitwiseand_89 (
        .y(_T_140),
        .a(io_inst),
        .b(32'h90000010)
    );
    wire _T_142;
    EQ_UNSIGNED #(.width(32)) u_eq_90 (
        .y(_T_142),
        .a(_T_140),
        .b(32'h80000010)
    );
    wire _T_144;
    BITWISEOR #(.width(1)) bitwiseor_91 (
        .y(_T_144),
        .a(1'h0),
        .b(_T_108)
    );
    wire decoder_10;
    BITWISEOR #(.width(1)) bitwiseor_92 (
        .y(decoder_10),
        .a(_T_144),
        .b(_T_142)
    );
    wire [31:0] _T_146;
    BITWISEAND #(.width(32)) bitwiseand_93 (
        .y(_T_146),
        .a(io_inst),
        .b(32'hA0000010)
    );
    wire _T_148;
    EQ_UNSIGNED #(.width(32)) u_eq_94 (
        .y(_T_148),
        .a(_T_146),
        .b(32'h20000010)
    );
    wire [31:0] _T_150;
    BITWISEAND #(.width(32)) bitwiseand_95 (
        .y(_T_150),
        .a(io_inst),
        .b(32'hD0000010)
    );
    wire _T_152;
    EQ_UNSIGNED #(.width(32)) u_eq_96 (
        .y(_T_152),
        .a(_T_150),
        .b(32'h40000010)
    );
    wire _T_154;
    BITWISEOR #(.width(1)) bitwiseor_97 (
        .y(_T_154),
        .a(1'h0),
        .b(_T_148)
    );
    wire decoder_11;
    BITWISEOR #(.width(1)) bitwiseor_98 (
        .y(decoder_11),
        .a(_T_154),
        .b(_T_152)
    );
    wire [31:0] _T_156;
    BITWISEAND #(.width(32)) bitwiseand_99 (
        .y(_T_156),
        .a(io_inst),
        .b(32'h70000004)
    );
    wire _T_158;
    EQ_UNSIGNED #(.width(32)) u_eq_100 (
        .y(_T_158),
        .a(_T_156),
        .b(32'h0)
    );
    wire [31:0] _T_160;
    BITWISEAND #(.width(32)) bitwiseand_101 (
        .y(_T_160),
        .a(io_inst),
        .b(32'h68000004)
    );
    wire _T_162;
    EQ_UNSIGNED #(.width(32)) u_eq_102 (
        .y(_T_162),
        .a(_T_160),
        .b(32'h0)
    );
    wire _T_164;
    BITWISEOR #(.width(1)) bitwiseor_103 (
        .y(_T_164),
        .a(1'h0),
        .b(_T_158)
    );
    wire _T_165;
    BITWISEOR #(.width(1)) bitwiseor_104 (
        .y(_T_165),
        .a(_T_164),
        .b(_T_162)
    );
    wire decoder_12;
    BITWISEOR #(.width(1)) bitwiseor_105 (
        .y(decoder_12),
        .a(_T_165),
        .b(_T_97)
    );
    wire [31:0] _T_167;
    BITWISEAND #(.width(32)) bitwiseand_106 (
        .y(_T_167),
        .a(io_inst),
        .b(32'h58000010)
    );
    wire _T_169;
    EQ_UNSIGNED #(.width(32)) u_eq_107 (
        .y(_T_169),
        .a(_T_167),
        .b(32'h18000010)
    );
    wire decoder_13;
    BITWISEOR #(.width(1)) bitwiseor_108 (
        .y(decoder_13),
        .a(1'h0),
        .b(_T_169)
    );
    wire [31:0] _T_172;
    BITWISEAND #(.width(32)) bitwiseand_109 (
        .y(_T_172),
        .a(io_inst),
        .b(32'hD0000010)
    );
    wire _T_174;
    EQ_UNSIGNED #(.width(32)) u_eq_110 (
        .y(_T_174),
        .a(_T_172),
        .b(32'h50000010)
    );
    wire decoder_14;
    BITWISEOR #(.width(1)) bitwiseor_111 (
        .y(decoder_14),
        .a(1'h0),
        .b(_T_174)
    );
    wire [31:0] _T_177;
    BITWISEAND #(.width(32)) bitwiseand_112 (
        .y(_T_177),
        .a(io_inst),
        .b(32'h20000004)
    );
    wire _T_179;
    EQ_UNSIGNED #(.width(32)) u_eq_113 (
        .y(_T_179),
        .a(_T_177),
        .b(32'h0)
    );
    wire [31:0] _T_181;
    BITWISEAND #(.width(32)) bitwiseand_114 (
        .y(_T_181),
        .a(io_inst),
        .b(32'h8002000)
    );
    wire _T_183;
    EQ_UNSIGNED #(.width(32)) u_eq_115 (
        .y(_T_183),
        .a(_T_181),
        .b(32'h8000000)
    );
    wire [31:0] _T_185;
    BITWISEAND #(.width(32)) bitwiseand_116 (
        .y(_T_185),
        .a(io_inst),
        .b(32'hC0000004)
    );
    wire _T_187;
    EQ_UNSIGNED #(.width(32)) u_eq_117 (
        .y(_T_187),
        .a(_T_185),
        .b(32'h80000000)
    );
    wire _T_189;
    BITWISEOR #(.width(1)) bitwiseor_118 (
        .y(_T_189),
        .a(1'h0),
        .b(_T_179)
    );
    wire _T_190;
    BITWISEOR #(.width(1)) bitwiseor_119 (
        .y(_T_190),
        .a(_T_189),
        .b(_T_97)
    );
    wire _T_191;
    BITWISEOR #(.width(1)) bitwiseor_120 (
        .y(_T_191),
        .a(_T_190),
        .b(_T_183)
    );
    wire decoder_15;
    BITWISEOR #(.width(1)) bitwiseor_121 (
        .y(decoder_15),
        .a(_T_191),
        .b(_T_187)
    );
    assign io_sigs_cmd = decoder_0;
    assign io_sigs_div = decoder_13;
    assign io_sigs_fastpipe = decoder_11;
    assign io_sigs_fma = decoder_12;
    assign io_sigs_fromint = decoder_9;
    assign io_sigs_ldst = decoder_1;
    assign io_sigs_ren1 = decoder_3;
    assign io_sigs_ren2 = decoder_4;
    assign io_sigs_ren3 = decoder_5;
    assign io_sigs_single = decoder_8;
    assign io_sigs_sqrt = decoder_14;
    assign io_sigs_swap12 = decoder_6;
    assign io_sigs_swap23 = decoder_7;
    assign io_sigs_toint = decoder_10;
    assign io_sigs_wen = decoder_2;
    assign io_sigs_wflags = decoder_15;
endmodule //FPUDecoder
module CAT(y, a, b);
    parameter width_a = 4;
    parameter width_b = 4;
    output [width_a+width_b-1:0] y;
    input [width_a-1:0] a;
    input [width_b-1:0] b;
    assign y = {a, b};
endmodule // CAT
module BITS(y, in);
    parameter width = 4;
    parameter high = 2;
    parameter low = 0;
    output [high-low:0] y;
    input [width-1:0] in;
    assign y = in[high:low];
endmodule // BITS
module PAD_UNSIGNED(y, in);
    parameter width = 4;
    parameter n = 4;
    output [(n > width ? n : width)-1:0] y;
    input [width-1:0] in;
    assign y = (n > width) ? {{(n - width){1'b0}}, in} : in;
endmodule // PAD_UNSIGNED
module SHL_UNSIGNED(y, in);
    parameter width = 4;
    parameter n = 4;
    output [width+n-1:0] y;
    input [width-1:0] in;
    wire [width+n-1:0] temp;
    assign temp = {{n{1'b0}}, in};
    assign y = temp << n;
endmodule // SHL_UNSIGNED
module NEQ_UNSIGNED(y, a, b);
    parameter width = 4;
    output y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a != b;
endmodule // NEQ_UNSIGNED
module BITWISENOT(y, in);
    parameter width = 4;
    output [width-1:0] y;
    input [width-1:0] in;
    assign y = ~in;
endmodule // BITWISENOT
module DSHL_UNSIGNED(y, in, n);
    parameter width_in = 4;
    parameter width_n = 2;
    output [(width_in+2**width_n-1)-1:0] y;
    input [width_in-1:0] in;
    input [width_n-1:0] n;
    wire [(width_in+2**width_n-1)-1:0] temp;
    assign temp = {{(2**width_n-1){1'b0}}, in};
    assign y = temp << n;
endmodule // DSHL_UNSIGNED
module BITWISEXOR(y, a, b);
    parameter width = 4;
    output [width-1:0] y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a ^ b;
endmodule // BITWISEXOR
module ADD_UNSIGNED(y, a, b);
    parameter width = 4;
    output [width:0] y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a + b;
endmodule // ADD_UNSIGNED
module TAIL(y, in);
    parameter width = 4;
    parameter n = 2;
    output [width-n-1:0] y;
    input [width-1:0] in;
    assign y = in[width-n-1:0];
endmodule // TAIL
module MRMWMEM(read_datas, read_clks, read_ens, read_addrs, write_clks, write_ens, write_masks, write_addrs, write_datas);
    parameter depth = 16;
    parameter addrbits = 4;
    parameter width = 32;
    parameter readernum = 2;
    parameter writernum = 2;
    parameter isSyncRead = 0;
    output [(width*readernum-1):0] read_datas;
    input [(1*readernum-1):0] read_clks;
    input [(1*readernum-1):0] read_ens;
    input [(addrbits*readernum-1):0] read_addrs;
    input [1*writernum-1:0] write_clks;
    input [1*writernum-1:0] write_ens;
    input [1*writernum-1:0] write_masks;
    input [(addrbits*writernum-1):0] write_addrs;
    input [(width*writernum-1):0] write_datas;
    reg [width-1:0] memcore [0:depth-1];
    wire [(addrbits*readernum-1):0] final_read_addrs;
    genvar gv_n;
    generate
        for (gv_n = 0; gv_n < readernum; gv_n = gv_n + 1) begin: get_final_raddrs
            if (isSyncRead) begin: raddr_processor
                reg [addrbits-1:0] read_addr_pipe_0;
                always @(posedge read_clks[gv_n]) begin
                    if (read_ens[gv_n]) begin
                        read_addr_pipe_0 <= read_addrs[gv_n*addrbits +: addrbits];
                    end
                end
                assign final_read_addrs[gv_n*addrbits +: addrbits] = read_addr_pipe_0;
            end else begin: raddr_processor
                assign final_read_addrs[gv_n*addrbits +: addrbits] = read_addrs[gv_n*addrbits +: addrbits];
            end
        end
    endgenerate
    genvar gv_k;
    generate
        for (gv_k = 0; gv_k < readernum; gv_k = gv_k + 1) begin: form_read_datas
            assign read_datas[gv_k*width +: width] = memcore[final_read_addrs[gv_k*addrbits +: addrbits]];
        end
    endgenerate
    integer i;
    always @(posedge write_clks[0]) begin
        for (i = 0; i < writernum; i = i + 1) begin
            if (write_ens[i] & write_masks[i]) begin
                memcore[write_addrs[i*addrbits +: addrbits]] <= write_datas[i*width +: width];
            end
        end
    end
endmodule // MRMWMEM
module FPUFMAPipe(
    input clock,
    input reset,
    input io_in_valid,
    input [4:0] io_in_bits_cmd,
    input io_in_bits_ldst,
    input io_in_bits_wen,
    input io_in_bits_ren1,
    input io_in_bits_ren2,
    input io_in_bits_ren3,
    input io_in_bits_swap12,
    input io_in_bits_swap23,
    input io_in_bits_single,
    input io_in_bits_fromint,
    input io_in_bits_toint,
    input io_in_bits_fastpipe,
    input io_in_bits_fma,
    input io_in_bits_div,
    input io_in_bits_sqrt,
    input io_in_bits_wflags,
    input [2:0] io_in_bits_rm,
    input [1:0] io_in_bits_typ,
    input [64:0] io_in_bits_in1,
    input [64:0] io_in_bits_in2,
    input [64:0] io_in_bits_in3,
    output io_out_valid,
    output [64:0] io_out_bits_data,
    output [4:0] io_out_bits_exc
);
    wire [31:0] one;
    assign one = 32'h80000000;
    wire _T_131;
    BITS #(.width(65), .high(32), .low(32)) bits_547 (
        .y(_T_131),
        .in(io_in_bits_in1)
    );
    wire _T_132;
    BITS #(.width(65), .high(32), .low(32)) bits_548 (
        .y(_T_132),
        .in(io_in_bits_in2)
    );
    wire _T_133;
    BITWISEXOR #(.width(1)) bitwisexor_549 (
        .y(_T_133),
        .a(_T_131),
        .b(_T_132)
    );
    wire [32:0] zero;
    SHL_UNSIGNED #(.width(1), .n(32)) u_shl_550 (
        .y(zero),
        .in(_T_133)
    );
    wire _valid__q;
    wire _valid__d;
    DFF_POSCLK #(.width(1)) valid (
        .q(_valid__q),
        .d(_valid__d),
        .clk(clock)
    );
    wire [4:0] _in_cmd__q;
    wire [4:0] _in_cmd__d;
    DFF_POSCLK #(.width(5)) in_cmd (
        .q(_in_cmd__q),
        .d(_in_cmd__d),
        .clk(clock)
    );
    wire _in_ldst__q;
    wire _in_ldst__d;
    DFF_POSCLK #(.width(1)) in_ldst (
        .q(_in_ldst__q),
        .d(_in_ldst__d),
        .clk(clock)
    );
    wire _in_wen__q;
    wire _in_wen__d;
    DFF_POSCLK #(.width(1)) in_wen (
        .q(_in_wen__q),
        .d(_in_wen__d),
        .clk(clock)
    );
    wire _in_ren1__q;
    wire _in_ren1__d;
    DFF_POSCLK #(.width(1)) in_ren1 (
        .q(_in_ren1__q),
        .d(_in_ren1__d),
        .clk(clock)
    );
    wire _in_ren2__q;
    wire _in_ren2__d;
    DFF_POSCLK #(.width(1)) in_ren2 (
        .q(_in_ren2__q),
        .d(_in_ren2__d),
        .clk(clock)
    );
    wire _in_ren3__q;
    wire _in_ren3__d;
    DFF_POSCLK #(.width(1)) in_ren3 (
        .q(_in_ren3__q),
        .d(_in_ren3__d),
        .clk(clock)
    );
    wire _in_swap12__q;
    wire _in_swap12__d;
    DFF_POSCLK #(.width(1)) in_swap12 (
        .q(_in_swap12__q),
        .d(_in_swap12__d),
        .clk(clock)
    );
    wire _in_swap23__q;
    wire _in_swap23__d;
    DFF_POSCLK #(.width(1)) in_swap23 (
        .q(_in_swap23__q),
        .d(_in_swap23__d),
        .clk(clock)
    );
    wire _in_single__q;
    wire _in_single__d;
    DFF_POSCLK #(.width(1)) in_single (
        .q(_in_single__q),
        .d(_in_single__d),
        .clk(clock)
    );
    wire _in_fromint__q;
    wire _in_fromint__d;
    DFF_POSCLK #(.width(1)) in_fromint (
        .q(_in_fromint__q),
        .d(_in_fromint__d),
        .clk(clock)
    );
    wire _in_toint__q;
    wire _in_toint__d;
    DFF_POSCLK #(.width(1)) in_toint (
        .q(_in_toint__q),
        .d(_in_toint__d),
        .clk(clock)
    );
    wire _in_fastpipe__q;
    wire _in_fastpipe__d;
    DFF_POSCLK #(.width(1)) in_fastpipe (
        .q(_in_fastpipe__q),
        .d(_in_fastpipe__d),
        .clk(clock)
    );
    wire _in_fma__q;
    wire _in_fma__d;
    DFF_POSCLK #(.width(1)) in_fma (
        .q(_in_fma__q),
        .d(_in_fma__d),
        .clk(clock)
    );
    wire _in_div__q;
    wire _in_div__d;
    DFF_POSCLK #(.width(1)) in_div (
        .q(_in_div__q),
        .d(_in_div__d),
        .clk(clock)
    );
    wire _in_sqrt__q;
    wire _in_sqrt__d;
    DFF_POSCLK #(.width(1)) in_sqrt (
        .q(_in_sqrt__q),
        .d(_in_sqrt__d),
        .clk(clock)
    );
    wire _in_wflags__q;
    wire _in_wflags__d;
    DFF_POSCLK #(.width(1)) in_wflags (
        .q(_in_wflags__q),
        .d(_in_wflags__d),
        .clk(clock)
    );
    wire [2:0] _in_rm__q;
    wire [2:0] _in_rm__d;
    DFF_POSCLK #(.width(3)) in_rm (
        .q(_in_rm__q),
        .d(_in_rm__d),
        .clk(clock)
    );
    wire [1:0] _in_typ__q;
    wire [1:0] _in_typ__d;
    DFF_POSCLK #(.width(2)) in_typ (
        .q(_in_typ__q),
        .d(_in_typ__d),
        .clk(clock)
    );
    wire [64:0] _in_in1__q;
    wire [64:0] _in_in1__d;
    DFF_POSCLK #(.width(65)) in_in1 (
        .q(_in_in1__q),
        .d(_in_in1__d),
        .clk(clock)
    );
    wire [64:0] _in_in2__q;
    wire [64:0] _in_in2__d;
    DFF_POSCLK #(.width(65)) in_in2 (
        .q(_in_in2__q),
        .d(_in_in2__d),
        .clk(clock)
    );
    wire [64:0] _in_in3__q;
    wire [64:0] _in_in3__d;
    DFF_POSCLK #(.width(65)) in_in3 (
        .q(_in_in3__q),
        .d(_in_in3__d),
        .clk(clock)
    );
    wire _T_177;
    BITS #(.width(5), .high(1), .low(1)) bits_551 (
        .y(_T_177),
        .in(io_in_bits_cmd)
    );
    wire _T_178;
    BITWISEOR #(.width(1)) bitwiseor_552 (
        .y(_T_178),
        .a(io_in_bits_ren3),
        .b(io_in_bits_swap23)
    );
    wire _T_179;
    BITWISEAND #(.width(1)) bitwiseand_553 (
        .y(_T_179),
        .a(_T_177),
        .b(_T_178)
    );
    wire _T_180;
    BITS #(.width(5), .high(0), .low(0)) bits_554 (
        .y(_T_180),
        .in(io_in_bits_cmd)
    );
    wire [1:0] _T_181;
    CAT #(.width_a(1), .width_b(1)) cat_555 (
        .y(_T_181),
        .a(_T_179),
        .b(_T_180)
    );
    wire _T_182;
    BITWISEOR #(.width(1)) bitwiseor_556 (
        .y(_T_182),
        .a(io_in_bits_ren3),
        .b(io_in_bits_swap23)
    );
    wire _T_184;
    EQ_UNSIGNED #(.width(1)) u_eq_557 (
        .y(_T_184),
        .a(_T_182),
        .b(1'h0)
    );
    wire [64:0] _node_15;
    wire [64:0] _WTEMP_71;
    PAD_UNSIGNED #(.width(32), .n(65)) u_pad_558 (
        .y(_WTEMP_71),
        .in(32'h80000000)
    );
    MUX_UNSIGNED #(.width(65)) u_mux_559 (
        .y(_node_15),
        .sel(io_in_bits_swap23),
        .a(_WTEMP_71),
        .b(io_in_bits_in2)
    );
    wire [64:0] _node_16;
    wire [64:0] _WTEMP_72;
    PAD_UNSIGNED #(.width(33), .n(65)) u_pad_560 (
        .y(_WTEMP_72),
        .in(zero)
    );
    MUX_UNSIGNED #(.width(65)) u_mux_561 (
        .y(_node_16),
        .sel(_T_184),
        .a(_WTEMP_72),
        .b(io_in_bits_in3)
    );
    wire _fma__clock;
    wire _fma__reset;
    wire [1:0] _fma__io_op;
    wire [32:0] _fma__io_a;
    wire [32:0] _fma__io_b;
    wire [32:0] _fma__io_c;
    wire [1:0] _fma__io_roundingMode;
    wire [32:0] _fma__io_out;
    wire [4:0] _fma__io_exceptionFlags;
    MulAddRecFN fma (
        .clock(_fma__clock),
        .reset(_fma__reset),
        .io_op(_fma__io_op),
        .io_a(_fma__io_a),
        .io_b(_fma__io_b),
        .io_c(_fma__io_c),
        .io_roundingMode(_fma__io_roundingMode),
        .io_out(_fma__io_out),
        .io_exceptionFlags(_fma__io_exceptionFlags)
    );
    wire [64:0] res_data;
    wire [4:0] res_exc;
    wire __T_192__q;
    wire __T_192__d;
    DFF_POSCLK #(.width(1)) _T_192 (
        .q(__T_192__q),
        .d(__T_192__d),
        .clk(clock)
    );
    wire _WTEMP_184;
    MUX_UNSIGNED #(.width(1)) u_mux_1421 (
        .y(__T_192__d),
        .sel(reset),
        .a(1'h0),
        .b(_WTEMP_184)
    );
    wire [64:0] __T_196_data__q;
    wire [64:0] __T_196_data__d;
    DFF_POSCLK #(.width(65)) _T_196_data (
        .q(__T_196_data__q),
        .d(__T_196_data__d),
        .clk(clock)
    );
    wire [4:0] __T_196_exc__q;
    wire [4:0] __T_196_exc__d;
    DFF_POSCLK #(.width(5)) _T_196_exc (
        .q(__T_196_exc__q),
        .d(__T_196_exc__d),
        .clk(clock)
    );
    wire __T_201__q;
    wire __T_201__d;
    DFF_POSCLK #(.width(1)) _T_201 (
        .q(__T_201__q),
        .d(__T_201__d),
        .clk(clock)
    );
    wire _WTEMP_185;
    MUX_UNSIGNED #(.width(1)) u_mux_1422 (
        .y(__T_201__d),
        .sel(reset),
        .a(1'h0),
        .b(_WTEMP_185)
    );
    wire [64:0] __T_205_data__q;
    wire [64:0] __T_205_data__d;
    DFF_POSCLK #(.width(65)) _T_205_data (
        .q(__T_205_data__q),
        .d(__T_205_data__d),
        .clk(clock)
    );
    wire [4:0] __T_205_exc__q;
    wire [4:0] __T_205_exc__d;
    DFF_POSCLK #(.width(5)) _T_205_exc (
        .q(__T_205_exc__q),
        .d(__T_205_exc__d),
        .clk(clock)
    );
    wire _T_217_valid;
    wire [64:0] _T_217_bits_data;
    wire [4:0] _T_217_bits_exc;
    assign _WTEMP_184 = _valid__q;
    MUX_UNSIGNED #(.width(65)) u_mux_1423 (
        .y(__T_196_data__d),
        .sel(_valid__q),
        .a(res_data),
        .b(__T_196_data__q)
    );
    MUX_UNSIGNED #(.width(5)) u_mux_1424 (
        .y(__T_196_exc__d),
        .sel(_valid__q),
        .a(res_exc),
        .b(__T_196_exc__q)
    );
    assign _WTEMP_185 = __T_192__q;
    MUX_UNSIGNED #(.width(65)) u_mux_1425 (
        .y(__T_205_data__d),
        .sel(__T_192__q),
        .a(__T_196_data__q),
        .b(__T_205_data__q)
    );
    MUX_UNSIGNED #(.width(5)) u_mux_1426 (
        .y(__T_205_exc__d),
        .sel(__T_192__q),
        .a(__T_196_exc__q),
        .b(__T_205_exc__q)
    );
    assign _T_217_bits_data = __T_205_data__q;
    assign _T_217_bits_exc = __T_205_exc__q;
    assign _T_217_valid = __T_201__q;
    assign _fma__clock = clock;
    BITS #(.width(65), .high(32), .low(0)) bits_1427 (
        .y(_fma__io_a),
        .in(_in_in1__q)
    );
    BITS #(.width(65), .high(32), .low(0)) bits_1428 (
        .y(_fma__io_b),
        .in(_in_in2__q)
    );
    BITS #(.width(65), .high(32), .low(0)) bits_1429 (
        .y(_fma__io_c),
        .in(_in_in3__q)
    );
    BITS #(.width(5), .high(1), .low(0)) bits_1430 (
        .y(_fma__io_op),
        .in(_in_cmd__q)
    );
    BITS #(.width(3), .high(1), .low(0)) bits_1431 (
        .y(_fma__io_roundingMode),
        .in(_in_rm__q)
    );
    assign _fma__reset = reset;
    wire [4:0] _WTEMP_186;
    PAD_UNSIGNED #(.width(2), .n(5)) u_pad_1432 (
        .y(_WTEMP_186),
        .in(_T_181)
    );
    MUX_UNSIGNED #(.width(5)) u_mux_1433 (
        .y(_in_cmd__d),
        .sel(io_in_valid),
        .a(_WTEMP_186),
        .b(_in_cmd__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_1434 (
        .y(_in_div__d),
        .sel(io_in_valid),
        .a(io_in_bits_div),
        .b(_in_div__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_1435 (
        .y(_in_fastpipe__d),
        .sel(io_in_valid),
        .a(io_in_bits_fastpipe),
        .b(_in_fastpipe__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_1436 (
        .y(_in_fma__d),
        .sel(io_in_valid),
        .a(io_in_bits_fma),
        .b(_in_fma__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_1437 (
        .y(_in_fromint__d),
        .sel(io_in_valid),
        .a(io_in_bits_fromint),
        .b(_in_fromint__q)
    );
    MUX_UNSIGNED #(.width(65)) u_mux_1438 (
        .y(_in_in1__d),
        .sel(io_in_valid),
        .a(io_in_bits_in1),
        .b(_in_in1__q)
    );
    MUX_UNSIGNED #(.width(65)) u_mux_1439 (
        .y(_in_in2__d),
        .sel(io_in_valid),
        .a(_node_15),
        .b(_in_in2__q)
    );
    MUX_UNSIGNED #(.width(65)) u_mux_1440 (
        .y(_in_in3__d),
        .sel(io_in_valid),
        .a(_node_16),
        .b(_in_in3__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_1441 (
        .y(_in_ldst__d),
        .sel(io_in_valid),
        .a(io_in_bits_ldst),
        .b(_in_ldst__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_1442 (
        .y(_in_ren1__d),
        .sel(io_in_valid),
        .a(io_in_bits_ren1),
        .b(_in_ren1__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_1443 (
        .y(_in_ren2__d),
        .sel(io_in_valid),
        .a(io_in_bits_ren2),
        .b(_in_ren2__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_1444 (
        .y(_in_ren3__d),
        .sel(io_in_valid),
        .a(io_in_bits_ren3),
        .b(_in_ren3__q)
    );
    MUX_UNSIGNED #(.width(3)) u_mux_1445 (
        .y(_in_rm__d),
        .sel(io_in_valid),
        .a(io_in_bits_rm),
        .b(_in_rm__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_1446 (
        .y(_in_single__d),
        .sel(io_in_valid),
        .a(io_in_bits_single),
        .b(_in_single__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_1447 (
        .y(_in_sqrt__d),
        .sel(io_in_valid),
        .a(io_in_bits_sqrt),
        .b(_in_sqrt__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_1448 (
        .y(_in_swap12__d),
        .sel(io_in_valid),
        .a(io_in_bits_swap12),
        .b(_in_swap12__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_1449 (
        .y(_in_swap23__d),
        .sel(io_in_valid),
        .a(io_in_bits_swap23),
        .b(_in_swap23__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_1450 (
        .y(_in_toint__d),
        .sel(io_in_valid),
        .a(io_in_bits_toint),
        .b(_in_toint__q)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_1451 (
        .y(_in_typ__d),
        .sel(io_in_valid),
        .a(io_in_bits_typ),
        .b(_in_typ__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_1452 (
        .y(_in_wen__d),
        .sel(io_in_valid),
        .a(io_in_bits_wen),
        .b(_in_wen__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_1453 (
        .y(_in_wflags__d),
        .sel(io_in_valid),
        .a(io_in_bits_wflags),
        .b(_in_wflags__q)
    );
    assign io_out_bits_data = _T_217_bits_data;
    assign io_out_bits_exc = _T_217_bits_exc;
    assign io_out_valid = _T_217_valid;
    PAD_UNSIGNED #(.width(33), .n(65)) u_pad_1454 (
        .y(res_data),
        .in(_fma__io_out)
    );
    assign res_exc = _fma__io_exceptionFlags;
    assign _valid__d = io_in_valid;
endmodule //FPUFMAPipe
module MulAddRecFN(
    input clock,
    input reset,
    input [1:0] io_op,
    input [32:0] io_a,
    input [32:0] io_b,
    input [32:0] io_c,
    input [1:0] io_roundingMode,
    output [32:0] io_out,
    output [4:0] io_exceptionFlags
);
    wire _mulAddRecFN_preMul__clock;
    wire _mulAddRecFN_preMul__reset;
    wire [1:0] _mulAddRecFN_preMul__io_op;
    wire [32:0] _mulAddRecFN_preMul__io_a;
    wire [32:0] _mulAddRecFN_preMul__io_b;
    wire [32:0] _mulAddRecFN_preMul__io_c;
    wire [1:0] _mulAddRecFN_preMul__io_roundingMode;
    wire [23:0] _mulAddRecFN_preMul__io_mulAddA;
    wire [23:0] _mulAddRecFN_preMul__io_mulAddB;
    wire [47:0] _mulAddRecFN_preMul__io_mulAddC;
    wire [2:0] _mulAddRecFN_preMul__io_toPostMul_highExpA;
    wire _mulAddRecFN_preMul__io_toPostMul_isNaN_isQuietNaNA;
    wire [2:0] _mulAddRecFN_preMul__io_toPostMul_highExpB;
    wire _mulAddRecFN_preMul__io_toPostMul_isNaN_isQuietNaNB;
    wire _mulAddRecFN_preMul__io_toPostMul_signProd;
    wire _mulAddRecFN_preMul__io_toPostMul_isZeroProd;
    wire _mulAddRecFN_preMul__io_toPostMul_opSignC;
    wire [2:0] _mulAddRecFN_preMul__io_toPostMul_highExpC;
    wire _mulAddRecFN_preMul__io_toPostMul_isNaN_isQuietNaNC;
    wire _mulAddRecFN_preMul__io_toPostMul_isCDominant;
    wire _mulAddRecFN_preMul__io_toPostMul_CAlignDist_0;
    wire [6:0] _mulAddRecFN_preMul__io_toPostMul_CAlignDist;
    wire _mulAddRecFN_preMul__io_toPostMul_bit0AlignedNegSigC;
    wire [25:0] _mulAddRecFN_preMul__io_toPostMul_highAlignedNegSigC;
    wire [10:0] _mulAddRecFN_preMul__io_toPostMul_sExpSum;
    wire [1:0] _mulAddRecFN_preMul__io_toPostMul_roundingMode;
    MulAddRecFN_preMul mulAddRecFN_preMul (
        .clock(_mulAddRecFN_preMul__clock),
        .reset(_mulAddRecFN_preMul__reset),
        .io_op(_mulAddRecFN_preMul__io_op),
        .io_a(_mulAddRecFN_preMul__io_a),
        .io_b(_mulAddRecFN_preMul__io_b),
        .io_c(_mulAddRecFN_preMul__io_c),
        .io_roundingMode(_mulAddRecFN_preMul__io_roundingMode),
        .io_mulAddA(_mulAddRecFN_preMul__io_mulAddA),
        .io_mulAddB(_mulAddRecFN_preMul__io_mulAddB),
        .io_mulAddC(_mulAddRecFN_preMul__io_mulAddC),
        .io_toPostMul_highExpA(_mulAddRecFN_preMul__io_toPostMul_highExpA),
        .io_toPostMul_isNaN_isQuietNaNA(_mulAddRecFN_preMul__io_toPostMul_isNaN_isQuietNaNA),
        .io_toPostMul_highExpB(_mulAddRecFN_preMul__io_toPostMul_highExpB),
        .io_toPostMul_isNaN_isQuietNaNB(_mulAddRecFN_preMul__io_toPostMul_isNaN_isQuietNaNB),
        .io_toPostMul_signProd(_mulAddRecFN_preMul__io_toPostMul_signProd),
        .io_toPostMul_isZeroProd(_mulAddRecFN_preMul__io_toPostMul_isZeroProd),
        .io_toPostMul_opSignC(_mulAddRecFN_preMul__io_toPostMul_opSignC),
        .io_toPostMul_highExpC(_mulAddRecFN_preMul__io_toPostMul_highExpC),
        .io_toPostMul_isNaN_isQuietNaNC(_mulAddRecFN_preMul__io_toPostMul_isNaN_isQuietNaNC),
        .io_toPostMul_isCDominant(_mulAddRecFN_preMul__io_toPostMul_isCDominant),
        .io_toPostMul_CAlignDist_0(_mulAddRecFN_preMul__io_toPostMul_CAlignDist_0),
        .io_toPostMul_CAlignDist(_mulAddRecFN_preMul__io_toPostMul_CAlignDist),
        .io_toPostMul_bit0AlignedNegSigC(_mulAddRecFN_preMul__io_toPostMul_bit0AlignedNegSigC),
        .io_toPostMul_highAlignedNegSigC(_mulAddRecFN_preMul__io_toPostMul_highAlignedNegSigC),
        .io_toPostMul_sExpSum(_mulAddRecFN_preMul__io_toPostMul_sExpSum),
        .io_toPostMul_roundingMode(_mulAddRecFN_preMul__io_toPostMul_roundingMode)
    );
    wire _mulAddRecFN_postMul__clock;
    wire _mulAddRecFN_postMul__reset;
    wire [2:0] _mulAddRecFN_postMul__io_fromPreMul_highExpA;
    wire _mulAddRecFN_postMul__io_fromPreMul_isNaN_isQuietNaNA;
    wire [2:0] _mulAddRecFN_postMul__io_fromPreMul_highExpB;
    wire _mulAddRecFN_postMul__io_fromPreMul_isNaN_isQuietNaNB;
    wire _mulAddRecFN_postMul__io_fromPreMul_signProd;
    wire _mulAddRecFN_postMul__io_fromPreMul_isZeroProd;
    wire _mulAddRecFN_postMul__io_fromPreMul_opSignC;
    wire [2:0] _mulAddRecFN_postMul__io_fromPreMul_highExpC;
    wire _mulAddRecFN_postMul__io_fromPreMul_isNaN_isQuietNaNC;
    wire _mulAddRecFN_postMul__io_fromPreMul_isCDominant;
    wire _mulAddRecFN_postMul__io_fromPreMul_CAlignDist_0;
    wire [6:0] _mulAddRecFN_postMul__io_fromPreMul_CAlignDist;
    wire _mulAddRecFN_postMul__io_fromPreMul_bit0AlignedNegSigC;
    wire [25:0] _mulAddRecFN_postMul__io_fromPreMul_highAlignedNegSigC;
    wire [10:0] _mulAddRecFN_postMul__io_fromPreMul_sExpSum;
    wire [1:0] _mulAddRecFN_postMul__io_fromPreMul_roundingMode;
    wire [48:0] _mulAddRecFN_postMul__io_mulAddResult;
    wire [32:0] _mulAddRecFN_postMul__io_out;
    wire [4:0] _mulAddRecFN_postMul__io_exceptionFlags;
    MulAddRecFN_postMul mulAddRecFN_postMul (
        .clock(_mulAddRecFN_postMul__clock),
        .reset(_mulAddRecFN_postMul__reset),
        .io_fromPreMul_highExpA(_mulAddRecFN_postMul__io_fromPreMul_highExpA),
        .io_fromPreMul_isNaN_isQuietNaNA(_mulAddRecFN_postMul__io_fromPreMul_isNaN_isQuietNaNA),
        .io_fromPreMul_highExpB(_mulAddRecFN_postMul__io_fromPreMul_highExpB),
        .io_fromPreMul_isNaN_isQuietNaNB(_mulAddRecFN_postMul__io_fromPreMul_isNaN_isQuietNaNB),
        .io_fromPreMul_signProd(_mulAddRecFN_postMul__io_fromPreMul_signProd),
        .io_fromPreMul_isZeroProd(_mulAddRecFN_postMul__io_fromPreMul_isZeroProd),
        .io_fromPreMul_opSignC(_mulAddRecFN_postMul__io_fromPreMul_opSignC),
        .io_fromPreMul_highExpC(_mulAddRecFN_postMul__io_fromPreMul_highExpC),
        .io_fromPreMul_isNaN_isQuietNaNC(_mulAddRecFN_postMul__io_fromPreMul_isNaN_isQuietNaNC),
        .io_fromPreMul_isCDominant(_mulAddRecFN_postMul__io_fromPreMul_isCDominant),
        .io_fromPreMul_CAlignDist_0(_mulAddRecFN_postMul__io_fromPreMul_CAlignDist_0),
        .io_fromPreMul_CAlignDist(_mulAddRecFN_postMul__io_fromPreMul_CAlignDist),
        .io_fromPreMul_bit0AlignedNegSigC(_mulAddRecFN_postMul__io_fromPreMul_bit0AlignedNegSigC),
        .io_fromPreMul_highAlignedNegSigC(_mulAddRecFN_postMul__io_fromPreMul_highAlignedNegSigC),
        .io_fromPreMul_sExpSum(_mulAddRecFN_postMul__io_fromPreMul_sExpSum),
        .io_fromPreMul_roundingMode(_mulAddRecFN_postMul__io_fromPreMul_roundingMode),
        .io_mulAddResult(_mulAddRecFN_postMul__io_mulAddResult),
        .io_out(_mulAddRecFN_postMul__io_out),
        .io_exceptionFlags(_mulAddRecFN_postMul__io_exceptionFlags)
    );
    wire [47:0] _T_16;
    MUL2_UNSIGNED #(.width_a(24), .width_b(24)) u_mul2_1416 (
        .y(_T_16),
        .a(_mulAddRecFN_preMul__io_mulAddA),
        .b(_mulAddRecFN_preMul__io_mulAddB)
    );
    wire [48:0] _T_18;
    CAT #(.width_a(1), .width_b(48)) cat_1417 (
        .y(_T_18),
        .a(1'h0),
        .b(_mulAddRecFN_preMul__io_mulAddC)
    );
    wire [49:0] _T_19;
    wire [48:0] _WTEMP_183;
    PAD_UNSIGNED #(.width(48), .n(49)) u_pad_1418 (
        .y(_WTEMP_183),
        .in(_T_16)
    );
    ADD_UNSIGNED #(.width(49)) u_add_1419 (
        .y(_T_19),
        .a(_WTEMP_183),
        .b(_T_18)
    );
    wire [48:0] _T_20;
    TAIL #(.width(50), .n(1)) tail_1420 (
        .y(_T_20),
        .in(_T_19)
    );
    assign io_exceptionFlags = _mulAddRecFN_postMul__io_exceptionFlags;
    assign io_out = _mulAddRecFN_postMul__io_out;
    assign _mulAddRecFN_postMul__clock = clock;
    assign _mulAddRecFN_postMul__io_fromPreMul_CAlignDist = _mulAddRecFN_preMul__io_toPostMul_CAlignDist;
    assign _mulAddRecFN_postMul__io_fromPreMul_CAlignDist_0 = _mulAddRecFN_preMul__io_toPostMul_CAlignDist_0;
    assign _mulAddRecFN_postMul__io_fromPreMul_bit0AlignedNegSigC = _mulAddRecFN_preMul__io_toPostMul_bit0AlignedNegSigC;
    assign _mulAddRecFN_postMul__io_fromPreMul_highAlignedNegSigC = _mulAddRecFN_preMul__io_toPostMul_highAlignedNegSigC;
    assign _mulAddRecFN_postMul__io_fromPreMul_highExpA = _mulAddRecFN_preMul__io_toPostMul_highExpA;
    assign _mulAddRecFN_postMul__io_fromPreMul_highExpB = _mulAddRecFN_preMul__io_toPostMul_highExpB;
    assign _mulAddRecFN_postMul__io_fromPreMul_highExpC = _mulAddRecFN_preMul__io_toPostMul_highExpC;
    assign _mulAddRecFN_postMul__io_fromPreMul_isCDominant = _mulAddRecFN_preMul__io_toPostMul_isCDominant;
    assign _mulAddRecFN_postMul__io_fromPreMul_isNaN_isQuietNaNA = _mulAddRecFN_preMul__io_toPostMul_isNaN_isQuietNaNA;
    assign _mulAddRecFN_postMul__io_fromPreMul_isNaN_isQuietNaNB = _mulAddRecFN_preMul__io_toPostMul_isNaN_isQuietNaNB;
    assign _mulAddRecFN_postMul__io_fromPreMul_isNaN_isQuietNaNC = _mulAddRecFN_preMul__io_toPostMul_isNaN_isQuietNaNC;
    assign _mulAddRecFN_postMul__io_fromPreMul_isZeroProd = _mulAddRecFN_preMul__io_toPostMul_isZeroProd;
    assign _mulAddRecFN_postMul__io_fromPreMul_opSignC = _mulAddRecFN_preMul__io_toPostMul_opSignC;
    assign _mulAddRecFN_postMul__io_fromPreMul_roundingMode = _mulAddRecFN_preMul__io_toPostMul_roundingMode;
    assign _mulAddRecFN_postMul__io_fromPreMul_sExpSum = _mulAddRecFN_preMul__io_toPostMul_sExpSum;
    assign _mulAddRecFN_postMul__io_fromPreMul_signProd = _mulAddRecFN_preMul__io_toPostMul_signProd;
    assign _mulAddRecFN_postMul__io_mulAddResult = _T_20;
    assign _mulAddRecFN_postMul__reset = reset;
    assign _mulAddRecFN_preMul__clock = clock;
    assign _mulAddRecFN_preMul__io_a = io_a;
    assign _mulAddRecFN_preMul__io_b = io_b;
    assign _mulAddRecFN_preMul__io_c = io_c;
    assign _mulAddRecFN_preMul__io_op = io_op;
    assign _mulAddRecFN_preMul__io_roundingMode = io_roundingMode;
    assign _mulAddRecFN_preMul__reset = reset;
endmodule //MulAddRecFN
module MulAddRecFN_preMul(
    input clock,
    input reset,
    input [1:0] io_op,
    input [32:0] io_a,
    input [32:0] io_b,
    input [32:0] io_c,
    input [1:0] io_roundingMode,
    output [23:0] io_mulAddA,
    output [23:0] io_mulAddB,
    output [47:0] io_mulAddC,
    output [2:0] io_toPostMul_highExpA,
    output io_toPostMul_isNaN_isQuietNaNA,
    output [2:0] io_toPostMul_highExpB,
    output io_toPostMul_isNaN_isQuietNaNB,
    output io_toPostMul_signProd,
    output io_toPostMul_isZeroProd,
    output io_toPostMul_opSignC,
    output [2:0] io_toPostMul_highExpC,
    output io_toPostMul_isNaN_isQuietNaNC,
    output io_toPostMul_isCDominant,
    output io_toPostMul_CAlignDist_0,
    output [6:0] io_toPostMul_CAlignDist,
    output io_toPostMul_bit0AlignedNegSigC,
    output [25:0] io_toPostMul_highAlignedNegSigC,
    output [10:0] io_toPostMul_sExpSum,
    output [1:0] io_toPostMul_roundingMode
);
    wire signA;
    BITS #(.width(33), .high(32), .low(32)) bits_562 (
        .y(signA),
        .in(io_a)
    );
    wire [8:0] expA;
    BITS #(.width(33), .high(31), .low(23)) bits_563 (
        .y(expA),
        .in(io_a)
    );
    wire [22:0] fractA;
    BITS #(.width(33), .high(22), .low(0)) bits_564 (
        .y(fractA),
        .in(io_a)
    );
    wire [2:0] _T_52;
    BITS #(.width(9), .high(8), .low(6)) bits_565 (
        .y(_T_52),
        .in(expA)
    );
    wire isZeroA;
    wire [2:0] _WTEMP_73;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_566 (
        .y(_WTEMP_73),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(3)) u_eq_567 (
        .y(isZeroA),
        .a(_T_52),
        .b(_WTEMP_73)
    );
    wire _T_55;
    EQ_UNSIGNED #(.width(1)) u_eq_568 (
        .y(_T_55),
        .a(isZeroA),
        .b(1'h0)
    );
    wire [23:0] sigA;
    CAT #(.width_a(1), .width_b(23)) cat_569 (
        .y(sigA),
        .a(_T_55),
        .b(fractA)
    );
    wire signB;
    BITS #(.width(33), .high(32), .low(32)) bits_570 (
        .y(signB),
        .in(io_b)
    );
    wire [8:0] expB;
    BITS #(.width(33), .high(31), .low(23)) bits_571 (
        .y(expB),
        .in(io_b)
    );
    wire [22:0] fractB;
    BITS #(.width(33), .high(22), .low(0)) bits_572 (
        .y(fractB),
        .in(io_b)
    );
    wire [2:0] _T_56;
    BITS #(.width(9), .high(8), .low(6)) bits_573 (
        .y(_T_56),
        .in(expB)
    );
    wire isZeroB;
    wire [2:0] _WTEMP_74;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_574 (
        .y(_WTEMP_74),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(3)) u_eq_575 (
        .y(isZeroB),
        .a(_T_56),
        .b(_WTEMP_74)
    );
    wire _T_59;
    EQ_UNSIGNED #(.width(1)) u_eq_576 (
        .y(_T_59),
        .a(isZeroB),
        .b(1'h0)
    );
    wire [23:0] sigB;
    CAT #(.width_a(1), .width_b(23)) cat_577 (
        .y(sigB),
        .a(_T_59),
        .b(fractB)
    );
    wire _T_60;
    BITS #(.width(33), .high(32), .low(32)) bits_578 (
        .y(_T_60),
        .in(io_c)
    );
    wire _T_61;
    BITS #(.width(2), .high(0), .low(0)) bits_579 (
        .y(_T_61),
        .in(io_op)
    );
    wire opSignC;
    BITWISEXOR #(.width(1)) bitwisexor_580 (
        .y(opSignC),
        .a(_T_60),
        .b(_T_61)
    );
    wire [8:0] expC;
    BITS #(.width(33), .high(31), .low(23)) bits_581 (
        .y(expC),
        .in(io_c)
    );
    wire [22:0] fractC;
    BITS #(.width(33), .high(22), .low(0)) bits_582 (
        .y(fractC),
        .in(io_c)
    );
    wire [2:0] _T_62;
    BITS #(.width(9), .high(8), .low(6)) bits_583 (
        .y(_T_62),
        .in(expC)
    );
    wire isZeroC;
    wire [2:0] _WTEMP_75;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_584 (
        .y(_WTEMP_75),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(3)) u_eq_585 (
        .y(isZeroC),
        .a(_T_62),
        .b(_WTEMP_75)
    );
    wire _T_65;
    EQ_UNSIGNED #(.width(1)) u_eq_586 (
        .y(_T_65),
        .a(isZeroC),
        .b(1'h0)
    );
    wire [23:0] sigC;
    CAT #(.width_a(1), .width_b(23)) cat_587 (
        .y(sigC),
        .a(_T_65),
        .b(fractC)
    );
    wire _T_66;
    BITWISEXOR #(.width(1)) bitwisexor_588 (
        .y(_T_66),
        .a(signA),
        .b(signB)
    );
    wire _T_67;
    BITS #(.width(2), .high(1), .low(1)) bits_589 (
        .y(_T_67),
        .in(io_op)
    );
    wire signProd;
    BITWISEXOR #(.width(1)) bitwisexor_590 (
        .y(signProd),
        .a(_T_66),
        .b(_T_67)
    );
    wire isZeroProd;
    BITWISEOR #(.width(1)) bitwiseor_591 (
        .y(isZeroProd),
        .a(isZeroA),
        .b(isZeroB)
    );
    wire _T_68;
    BITS #(.width(9), .high(8), .low(8)) bits_592 (
        .y(_T_68),
        .in(expB)
    );
    wire _T_70;
    EQ_UNSIGNED #(.width(1)) u_eq_593 (
        .y(_T_70),
        .a(_T_68),
        .b(1'h0)
    );
    wire _T_71;
    BITS #(.width(1), .high(0), .low(0)) bits_594 (
        .y(_T_71),
        .in(_T_70)
    );
    wire [2:0] _T_74;
    MUX_UNSIGNED #(.width(3)) u_mux_595 (
        .y(_T_74),
        .sel(_T_71),
        .a(3'h7),
        .b(3'h0)
    );
    wire [7:0] _T_75;
    BITS #(.width(9), .high(7), .low(0)) bits_596 (
        .y(_T_75),
        .in(expB)
    );
    wire [10:0] _T_76;
    CAT #(.width_a(3), .width_b(8)) cat_597 (
        .y(_T_76),
        .a(_T_74),
        .b(_T_75)
    );
    wire [11:0] _T_77;
    wire [10:0] _WTEMP_76;
    PAD_UNSIGNED #(.width(9), .n(11)) u_pad_598 (
        .y(_WTEMP_76),
        .in(expA)
    );
    ADD_UNSIGNED #(.width(11)) u_add_599 (
        .y(_T_77),
        .a(_WTEMP_76),
        .b(_T_76)
    );
    wire [10:0] _T_78;
    TAIL #(.width(12), .n(1)) tail_600 (
        .y(_T_78),
        .in(_T_77)
    );
    wire [11:0] _T_80;
    wire [10:0] _WTEMP_77;
    PAD_UNSIGNED #(.width(5), .n(11)) u_pad_601 (
        .y(_WTEMP_77),
        .in(5'h1B)
    );
    ADD_UNSIGNED #(.width(11)) u_add_602 (
        .y(_T_80),
        .a(_T_78),
        .b(_WTEMP_77)
    );
    wire [10:0] sExpAlignedProd;
    TAIL #(.width(12), .n(1)) tail_603 (
        .y(sExpAlignedProd),
        .in(_T_80)
    );
    wire doSubMags;
    BITWISEXOR #(.width(1)) bitwisexor_604 (
        .y(doSubMags),
        .a(signProd),
        .b(opSignC)
    );
    wire [11:0] _T_81;
    wire [10:0] _WTEMP_78;
    PAD_UNSIGNED #(.width(9), .n(11)) u_pad_605 (
        .y(_WTEMP_78),
        .in(expC)
    );
    SUB_UNSIGNED #(.width(11)) u_sub_606 (
        .y(_T_81),
        .a(sExpAlignedProd),
        .b(_WTEMP_78)
    );
    wire [11:0] _T_82;
    ASUINT #(.width(12)) asuint_607 (
        .y(_T_82),
        .in(_T_81)
    );
    wire [10:0] sNatCAlignDist;
    TAIL #(.width(12), .n(1)) tail_608 (
        .y(sNatCAlignDist),
        .in(_T_82)
    );
    wire _T_83;
    BITS #(.width(11), .high(10), .low(10)) bits_609 (
        .y(_T_83),
        .in(sNatCAlignDist)
    );
    wire CAlignDist_floor;
    BITWISEOR #(.width(1)) bitwiseor_610 (
        .y(CAlignDist_floor),
        .a(isZeroProd),
        .b(_T_83)
    );
    wire [9:0] _T_84;
    BITS #(.width(11), .high(9), .low(0)) bits_611 (
        .y(_T_84),
        .in(sNatCAlignDist)
    );
    wire _T_86;
    wire [9:0] _WTEMP_79;
    PAD_UNSIGNED #(.width(1), .n(10)) u_pad_612 (
        .y(_WTEMP_79),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(10)) u_eq_613 (
        .y(_T_86),
        .a(_T_84),
        .b(_WTEMP_79)
    );
    wire CAlignDist_0;
    BITWISEOR #(.width(1)) bitwiseor_614 (
        .y(CAlignDist_0),
        .a(CAlignDist_floor),
        .b(_T_86)
    );
    wire _T_88;
    EQ_UNSIGNED #(.width(1)) u_eq_615 (
        .y(_T_88),
        .a(isZeroC),
        .b(1'h0)
    );
    wire [9:0] _T_89;
    BITS #(.width(11), .high(9), .low(0)) bits_616 (
        .y(_T_89),
        .in(sNatCAlignDist)
    );
    wire _T_91;
    wire [9:0] _WTEMP_80;
    PAD_UNSIGNED #(.width(5), .n(10)) u_pad_617 (
        .y(_WTEMP_80),
        .in(5'h19)
    );
    LT_UNSIGNED #(.width(10)) u_lt_618 (
        .y(_T_91),
        .a(_T_89),
        .b(_WTEMP_80)
    );
    wire _T_92;
    BITWISEOR #(.width(1)) bitwiseor_619 (
        .y(_T_92),
        .a(CAlignDist_floor),
        .b(_T_91)
    );
    wire isCDominant;
    BITWISEAND #(.width(1)) bitwiseand_620 (
        .y(isCDominant),
        .a(_T_88),
        .b(_T_92)
    );
    wire [9:0] _T_94;
    BITS #(.width(11), .high(9), .low(0)) bits_621 (
        .y(_T_94),
        .in(sNatCAlignDist)
    );
    wire _T_96;
    wire [9:0] _WTEMP_81;
    PAD_UNSIGNED #(.width(7), .n(10)) u_pad_622 (
        .y(_WTEMP_81),
        .in(7'h4A)
    );
    LT_UNSIGNED #(.width(10)) u_lt_623 (
        .y(_T_96),
        .a(_T_94),
        .b(_WTEMP_81)
    );
    wire [6:0] _T_97;
    BITS #(.width(11), .high(6), .low(0)) bits_624 (
        .y(_T_97),
        .in(sNatCAlignDist)
    );
    wire [6:0] _T_99;
    MUX_UNSIGNED #(.width(7)) u_mux_625 (
        .y(_T_99),
        .sel(_T_96),
        .a(_T_97),
        .b(7'h4A)
    );
    wire [6:0] CAlignDist;
    wire [6:0] _WTEMP_82;
    PAD_UNSIGNED #(.width(1), .n(7)) u_pad_626 (
        .y(_WTEMP_82),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(7)) u_mux_627 (
        .y(CAlignDist),
        .sel(CAlignDist_floor),
        .a(_WTEMP_82),
        .b(_T_99)
    );
    wire [10:0] sExpSum;
    wire [10:0] _WTEMP_83;
    PAD_UNSIGNED #(.width(9), .n(11)) u_pad_628 (
        .y(_WTEMP_83),
        .in(expC)
    );
    MUX_UNSIGNED #(.width(11)) u_mux_629 (
        .y(sExpSum),
        .sel(CAlignDist_floor),
        .a(_WTEMP_83),
        .b(sExpAlignedProd)
    );
    wire _T_100;
    BITS #(.width(7), .high(6), .low(6)) bits_630 (
        .y(_T_100),
        .in(CAlignDist)
    );
    wire [5:0] _T_101;
    BITS #(.width(7), .high(5), .low(0)) bits_631 (
        .y(_T_101),
        .in(CAlignDist)
    );
    wire [64:0] _T_103;
    DSHR_SIGNED #(.width_in(65), .width_n(6)) s_dshr_632 (
        .y(_T_103),
        .in(-65'sh10000000000000000),
        .n(_T_101)
    );
    wire [9:0] _T_104;
    BITS #(.width(65), .high(63), .low(54)) bits_633 (
        .y(_T_104),
        .in(_T_103)
    );
    wire [7:0] _T_105;
    BITS #(.width(10), .high(7), .low(0)) bits_634 (
        .y(_T_105),
        .in(_T_104)
    );
    wire [7:0] _T_108;
    assign _T_108 = 8'hF0;
    wire [7:0] _T_109;
    assign _T_109 = 8'hF;
    wire [3:0] _T_110;
    SHR_UNSIGNED #(.width(8), .n(4)) u_shr_635 (
        .y(_T_110),
        .in(_T_105)
    );
    wire [7:0] _T_111;
    wire [7:0] _WTEMP_84;
    PAD_UNSIGNED #(.width(4), .n(8)) u_pad_636 (
        .y(_WTEMP_84),
        .in(_T_110)
    );
    BITWISEAND #(.width(8)) bitwiseand_637 (
        .y(_T_111),
        .a(_WTEMP_84),
        .b(_T_109)
    );
    wire [3:0] _T_112;
    BITS #(.width(8), .high(3), .low(0)) bits_638 (
        .y(_T_112),
        .in(_T_105)
    );
    wire [7:0] _T_113;
    SHL_UNSIGNED #(.width(4), .n(4)) u_shl_639 (
        .y(_T_113),
        .in(_T_112)
    );
    wire [7:0] _T_114;
    assign _T_114 = 8'hF0;
    wire [7:0] _T_115;
    BITWISEAND #(.width(8)) bitwiseand_640 (
        .y(_T_115),
        .a(_T_113),
        .b(_T_114)
    );
    wire [7:0] _T_116;
    BITWISEOR #(.width(8)) bitwiseor_641 (
        .y(_T_116),
        .a(_T_111),
        .b(_T_115)
    );
    wire [5:0] _T_117;
    assign _T_117 = 6'hF;
    wire [7:0] _T_118;
    assign _T_118 = 8'h3C;
    wire [7:0] _T_119;
    assign _T_119 = 8'h33;
    wire [5:0] _T_120;
    SHR_UNSIGNED #(.width(8), .n(2)) u_shr_642 (
        .y(_T_120),
        .in(_T_116)
    );
    wire [7:0] _T_121;
    wire [7:0] _WTEMP_85;
    PAD_UNSIGNED #(.width(6), .n(8)) u_pad_643 (
        .y(_WTEMP_85),
        .in(_T_120)
    );
    BITWISEAND #(.width(8)) bitwiseand_644 (
        .y(_T_121),
        .a(_WTEMP_85),
        .b(_T_119)
    );
    wire [5:0] _T_122;
    BITS #(.width(8), .high(5), .low(0)) bits_645 (
        .y(_T_122),
        .in(_T_116)
    );
    wire [7:0] _T_123;
    SHL_UNSIGNED #(.width(6), .n(2)) u_shl_646 (
        .y(_T_123),
        .in(_T_122)
    );
    wire [7:0] _T_124;
    assign _T_124 = 8'hCC;
    wire [7:0] _T_125;
    BITWISEAND #(.width(8)) bitwiseand_647 (
        .y(_T_125),
        .a(_T_123),
        .b(_T_124)
    );
    wire [7:0] _T_126;
    BITWISEOR #(.width(8)) bitwiseor_648 (
        .y(_T_126),
        .a(_T_121),
        .b(_T_125)
    );
    wire [6:0] _T_127;
    assign _T_127 = 7'h33;
    wire [7:0] _T_128;
    assign _T_128 = 8'h66;
    wire [7:0] _T_129;
    assign _T_129 = 8'h55;
    wire [6:0] _T_130;
    SHR_UNSIGNED #(.width(8), .n(1)) u_shr_649 (
        .y(_T_130),
        .in(_T_126)
    );
    wire [7:0] _T_131;
    wire [7:0] _WTEMP_86;
    PAD_UNSIGNED #(.width(7), .n(8)) u_pad_650 (
        .y(_WTEMP_86),
        .in(_T_130)
    );
    BITWISEAND #(.width(8)) bitwiseand_651 (
        .y(_T_131),
        .a(_WTEMP_86),
        .b(_T_129)
    );
    wire [6:0] _T_132;
    BITS #(.width(8), .high(6), .low(0)) bits_652 (
        .y(_T_132),
        .in(_T_126)
    );
    wire [7:0] _T_133;
    SHL_UNSIGNED #(.width(7), .n(1)) u_shl_653 (
        .y(_T_133),
        .in(_T_132)
    );
    wire [7:0] _T_134;
    assign _T_134 = 8'hAA;
    wire [7:0] _T_135;
    BITWISEAND #(.width(8)) bitwiseand_654 (
        .y(_T_135),
        .a(_T_133),
        .b(_T_134)
    );
    wire [7:0] _T_136;
    BITWISEOR #(.width(8)) bitwiseor_655 (
        .y(_T_136),
        .a(_T_131),
        .b(_T_135)
    );
    wire [1:0] _T_137;
    BITS #(.width(10), .high(9), .low(8)) bits_656 (
        .y(_T_137),
        .in(_T_104)
    );
    wire _T_138;
    BITS #(.width(2), .high(0), .low(0)) bits_657 (
        .y(_T_138),
        .in(_T_137)
    );
    wire _T_139;
    BITS #(.width(2), .high(1), .low(1)) bits_658 (
        .y(_T_139),
        .in(_T_137)
    );
    wire [1:0] _T_140;
    CAT #(.width_a(1), .width_b(1)) cat_659 (
        .y(_T_140),
        .a(_T_138),
        .b(_T_139)
    );
    wire [9:0] _T_141;
    CAT #(.width_a(8), .width_b(2)) cat_660 (
        .y(_T_141),
        .a(_T_136),
        .b(_T_140)
    );
    wire [23:0] _T_143;
    CAT #(.width_a(10), .width_b(14)) cat_661 (
        .y(_T_143),
        .a(_T_141),
        .b(14'h3FFF)
    );
    wire [64:0] _T_145;
    DSHR_SIGNED #(.width_in(65), .width_n(6)) s_dshr_662 (
        .y(_T_145),
        .in(-65'sh10000000000000000),
        .n(_T_101)
    );
    wire [13:0] _T_146;
    BITS #(.width(65), .high(13), .low(0)) bits_663 (
        .y(_T_146),
        .in(_T_145)
    );
    wire [7:0] _T_147;
    BITS #(.width(14), .high(7), .low(0)) bits_664 (
        .y(_T_147),
        .in(_T_146)
    );
    wire [7:0] _T_150;
    assign _T_150 = 8'hF0;
    wire [7:0] _T_151;
    assign _T_151 = 8'hF;
    wire [3:0] _T_152;
    SHR_UNSIGNED #(.width(8), .n(4)) u_shr_665 (
        .y(_T_152),
        .in(_T_147)
    );
    wire [7:0] _T_153;
    wire [7:0] _WTEMP_87;
    PAD_UNSIGNED #(.width(4), .n(8)) u_pad_666 (
        .y(_WTEMP_87),
        .in(_T_152)
    );
    BITWISEAND #(.width(8)) bitwiseand_667 (
        .y(_T_153),
        .a(_WTEMP_87),
        .b(_T_151)
    );
    wire [3:0] _T_154;
    BITS #(.width(8), .high(3), .low(0)) bits_668 (
        .y(_T_154),
        .in(_T_147)
    );
    wire [7:0] _T_155;
    SHL_UNSIGNED #(.width(4), .n(4)) u_shl_669 (
        .y(_T_155),
        .in(_T_154)
    );
    wire [7:0] _T_156;
    assign _T_156 = 8'hF0;
    wire [7:0] _T_157;
    BITWISEAND #(.width(8)) bitwiseand_670 (
        .y(_T_157),
        .a(_T_155),
        .b(_T_156)
    );
    wire [7:0] _T_158;
    BITWISEOR #(.width(8)) bitwiseor_671 (
        .y(_T_158),
        .a(_T_153),
        .b(_T_157)
    );
    wire [5:0] _T_159;
    assign _T_159 = 6'hF;
    wire [7:0] _T_160;
    assign _T_160 = 8'h3C;
    wire [7:0] _T_161;
    assign _T_161 = 8'h33;
    wire [5:0] _T_162;
    SHR_UNSIGNED #(.width(8), .n(2)) u_shr_672 (
        .y(_T_162),
        .in(_T_158)
    );
    wire [7:0] _T_163;
    wire [7:0] _WTEMP_88;
    PAD_UNSIGNED #(.width(6), .n(8)) u_pad_673 (
        .y(_WTEMP_88),
        .in(_T_162)
    );
    BITWISEAND #(.width(8)) bitwiseand_674 (
        .y(_T_163),
        .a(_WTEMP_88),
        .b(_T_161)
    );
    wire [5:0] _T_164;
    BITS #(.width(8), .high(5), .low(0)) bits_675 (
        .y(_T_164),
        .in(_T_158)
    );
    wire [7:0] _T_165;
    SHL_UNSIGNED #(.width(6), .n(2)) u_shl_676 (
        .y(_T_165),
        .in(_T_164)
    );
    wire [7:0] _T_166;
    assign _T_166 = 8'hCC;
    wire [7:0] _T_167;
    BITWISEAND #(.width(8)) bitwiseand_677 (
        .y(_T_167),
        .a(_T_165),
        .b(_T_166)
    );
    wire [7:0] _T_168;
    BITWISEOR #(.width(8)) bitwiseor_678 (
        .y(_T_168),
        .a(_T_163),
        .b(_T_167)
    );
    wire [6:0] _T_169;
    assign _T_169 = 7'h33;
    wire [7:0] _T_170;
    assign _T_170 = 8'h66;
    wire [7:0] _T_171;
    assign _T_171 = 8'h55;
    wire [6:0] _T_172;
    SHR_UNSIGNED #(.width(8), .n(1)) u_shr_679 (
        .y(_T_172),
        .in(_T_168)
    );
    wire [7:0] _T_173;
    wire [7:0] _WTEMP_89;
    PAD_UNSIGNED #(.width(7), .n(8)) u_pad_680 (
        .y(_WTEMP_89),
        .in(_T_172)
    );
    BITWISEAND #(.width(8)) bitwiseand_681 (
        .y(_T_173),
        .a(_WTEMP_89),
        .b(_T_171)
    );
    wire [6:0] _T_174;
    BITS #(.width(8), .high(6), .low(0)) bits_682 (
        .y(_T_174),
        .in(_T_168)
    );
    wire [7:0] _T_175;
    SHL_UNSIGNED #(.width(7), .n(1)) u_shl_683 (
        .y(_T_175),
        .in(_T_174)
    );
    wire [7:0] _T_176;
    assign _T_176 = 8'hAA;
    wire [7:0] _T_177;
    BITWISEAND #(.width(8)) bitwiseand_684 (
        .y(_T_177),
        .a(_T_175),
        .b(_T_176)
    );
    wire [7:0] _T_178;
    BITWISEOR #(.width(8)) bitwiseor_685 (
        .y(_T_178),
        .a(_T_173),
        .b(_T_177)
    );
    wire [5:0] _T_179;
    BITS #(.width(14), .high(13), .low(8)) bits_686 (
        .y(_T_179),
        .in(_T_146)
    );
    wire [3:0] _T_180;
    BITS #(.width(6), .high(3), .low(0)) bits_687 (
        .y(_T_180),
        .in(_T_179)
    );
    wire [1:0] _T_181;
    BITS #(.width(4), .high(1), .low(0)) bits_688 (
        .y(_T_181),
        .in(_T_180)
    );
    wire _T_182;
    BITS #(.width(2), .high(0), .low(0)) bits_689 (
        .y(_T_182),
        .in(_T_181)
    );
    wire _T_183;
    BITS #(.width(2), .high(1), .low(1)) bits_690 (
        .y(_T_183),
        .in(_T_181)
    );
    wire [1:0] _T_184;
    CAT #(.width_a(1), .width_b(1)) cat_691 (
        .y(_T_184),
        .a(_T_182),
        .b(_T_183)
    );
    wire [1:0] _T_185;
    BITS #(.width(4), .high(3), .low(2)) bits_692 (
        .y(_T_185),
        .in(_T_180)
    );
    wire _T_186;
    BITS #(.width(2), .high(0), .low(0)) bits_693 (
        .y(_T_186),
        .in(_T_185)
    );
    wire _T_187;
    BITS #(.width(2), .high(1), .low(1)) bits_694 (
        .y(_T_187),
        .in(_T_185)
    );
    wire [1:0] _T_188;
    CAT #(.width_a(1), .width_b(1)) cat_695 (
        .y(_T_188),
        .a(_T_186),
        .b(_T_187)
    );
    wire [3:0] _T_189;
    CAT #(.width_a(2), .width_b(2)) cat_696 (
        .y(_T_189),
        .a(_T_184),
        .b(_T_188)
    );
    wire [1:0] _T_190;
    BITS #(.width(6), .high(5), .low(4)) bits_697 (
        .y(_T_190),
        .in(_T_179)
    );
    wire _T_191;
    BITS #(.width(2), .high(0), .low(0)) bits_698 (
        .y(_T_191),
        .in(_T_190)
    );
    wire _T_192;
    BITS #(.width(2), .high(1), .low(1)) bits_699 (
        .y(_T_192),
        .in(_T_190)
    );
    wire [1:0] _T_193;
    CAT #(.width_a(1), .width_b(1)) cat_700 (
        .y(_T_193),
        .a(_T_191),
        .b(_T_192)
    );
    wire [5:0] _T_194;
    CAT #(.width_a(4), .width_b(2)) cat_701 (
        .y(_T_194),
        .a(_T_189),
        .b(_T_193)
    );
    wire [13:0] _T_195;
    CAT #(.width_a(8), .width_b(6)) cat_702 (
        .y(_T_195),
        .a(_T_178),
        .b(_T_194)
    );
    wire [23:0] CExtraMask;
    wire [23:0] _WTEMP_90;
    PAD_UNSIGNED #(.width(14), .n(24)) u_pad_703 (
        .y(_WTEMP_90),
        .in(_T_195)
    );
    MUX_UNSIGNED #(.width(24)) u_mux_704 (
        .y(CExtraMask),
        .sel(_T_100),
        .a(_T_143),
        .b(_WTEMP_90)
    );
    wire [23:0] _T_196;
    BITWISENOT #(.width(24)) bitwisenot_705 (
        .y(_T_196),
        .in(sigC)
    );
    wire [23:0] negSigC;
    MUX_UNSIGNED #(.width(24)) u_mux_706 (
        .y(negSigC),
        .sel(doSubMags),
        .a(_T_196),
        .b(sigC)
    );
    wire _T_197;
    BITS #(.width(1), .high(0), .low(0)) bits_707 (
        .y(_T_197),
        .in(doSubMags)
    );
    wire [49:0] _T_200;
    MUX_UNSIGNED #(.width(50)) u_mux_708 (
        .y(_T_200),
        .sel(_T_197),
        .a(50'h3FFFFFFFFFFFF),
        .b(50'h0)
    );
    wire [24:0] _T_201;
    CAT #(.width_a(1), .width_b(24)) cat_709 (
        .y(_T_201),
        .a(doSubMags),
        .b(negSigC)
    );
    wire [74:0] _T_202;
    CAT #(.width_a(25), .width_b(50)) cat_710 (
        .y(_T_202),
        .a(_T_201),
        .b(_T_200)
    );
    wire [74:0] _T_203;
    ASSINT #(.width(75)) assint_711 (
        .y(_T_203),
        .in(_T_202)
    );
    wire [74:0] _T_204;
    DSHR_SIGNED #(.width_in(75), .width_n(7)) s_dshr_712 (
        .y(_T_204),
        .in(_T_203),
        .n(CAlignDist)
    );
    wire [23:0] _T_205;
    BITWISEAND #(.width(24)) bitwiseand_713 (
        .y(_T_205),
        .a(sigC),
        .b(CExtraMask)
    );
    wire _T_207;
    wire [23:0] _WTEMP_91;
    PAD_UNSIGNED #(.width(1), .n(24)) u_pad_714 (
        .y(_WTEMP_91),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(24)) u_neq_715 (
        .y(_T_207),
        .a(_T_205),
        .b(_WTEMP_91)
    );
    wire _T_208;
    BITWISEXOR #(.width(1)) bitwisexor_716 (
        .y(_T_208),
        .a(_T_207),
        .b(doSubMags)
    );
    wire [74:0] _T_209;
    ASUINT #(.width(75)) asuint_717 (
        .y(_T_209),
        .in(_T_204)
    );
    wire [75:0] _T_210;
    CAT #(.width_a(75), .width_b(1)) cat_718 (
        .y(_T_210),
        .a(_T_209),
        .b(_T_208)
    );
    wire [74:0] alignedNegSigC;
    BITS #(.width(76), .high(74), .low(0)) bits_719 (
        .y(alignedNegSigC),
        .in(_T_210)
    );
    wire [47:0] _T_211;
    BITS #(.width(75), .high(48), .low(1)) bits_720 (
        .y(_T_211),
        .in(alignedNegSigC)
    );
    wire [2:0] _T_212;
    BITS #(.width(9), .high(8), .low(6)) bits_721 (
        .y(_T_212),
        .in(expA)
    );
    wire _T_213;
    BITS #(.width(23), .high(22), .low(22)) bits_722 (
        .y(_T_213),
        .in(fractA)
    );
    wire [2:0] _T_214;
    BITS #(.width(9), .high(8), .low(6)) bits_723 (
        .y(_T_214),
        .in(expB)
    );
    wire _T_215;
    BITS #(.width(23), .high(22), .low(22)) bits_724 (
        .y(_T_215),
        .in(fractB)
    );
    wire [2:0] _T_216;
    BITS #(.width(9), .high(8), .low(6)) bits_725 (
        .y(_T_216),
        .in(expC)
    );
    wire _T_217;
    BITS #(.width(23), .high(22), .low(22)) bits_726 (
        .y(_T_217),
        .in(fractC)
    );
    wire _T_218;
    BITS #(.width(75), .high(0), .low(0)) bits_727 (
        .y(_T_218),
        .in(alignedNegSigC)
    );
    wire [25:0] _T_219;
    BITS #(.width(75), .high(74), .low(49)) bits_728 (
        .y(_T_219),
        .in(alignedNegSigC)
    );
    assign io_mulAddA = sigA;
    assign io_mulAddB = sigB;
    assign io_mulAddC = _T_211;
    assign io_toPostMul_CAlignDist = CAlignDist;
    assign io_toPostMul_CAlignDist_0 = CAlignDist_0;
    assign io_toPostMul_bit0AlignedNegSigC = _T_218;
    assign io_toPostMul_highAlignedNegSigC = _T_219;
    assign io_toPostMul_highExpA = _T_212;
    assign io_toPostMul_highExpB = _T_214;
    assign io_toPostMul_highExpC = _T_216;
    assign io_toPostMul_isCDominant = isCDominant;
    assign io_toPostMul_isNaN_isQuietNaNA = _T_213;
    assign io_toPostMul_isNaN_isQuietNaNB = _T_215;
    assign io_toPostMul_isNaN_isQuietNaNC = _T_217;
    assign io_toPostMul_isZeroProd = isZeroProd;
    assign io_toPostMul_opSignC = opSignC;
    assign io_toPostMul_roundingMode = io_roundingMode;
    assign io_toPostMul_sExpSum = sExpSum;
    assign io_toPostMul_signProd = signProd;
endmodule //MulAddRecFN_preMul
module SUB_UNSIGNED(y, a, b);
    parameter width = 4;
    output [width:0] y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a - b;
endmodule // SUB_UNSIGNED
module ASUINT(y, in);
    parameter width = 4;
    output [width-1:0] y;
    input [width-1:0] in;
    assign y = $unsigned(in);
endmodule // ASUINT
module LT_UNSIGNED(y, a, b);
    parameter width = 4;
    output y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a < b;
endmodule // LT_UNSIGNED
module DSHR_SIGNED(y, in, n);
    parameter width_in = 4;
    parameter width_n = 2;
    output [width_in-1:0] y;
    input [width_in-1:0] in;
    input [width_n-1:0] n;
    assign y = $signed(in) >>> n;
endmodule // DSHR_SIGNED
module SHR_UNSIGNED(y, in);
    parameter width = 4;
    parameter n = 2;
    output [(n < width ? (width-n-1) : 0):0] y;
    input [width-1:0] in;
    assign y = n < width ? in[width-1:n] : 1'b0;
endmodule // SHR_UNSIGNED
module ASSINT(y, in);
    parameter width = 4;
    output [width-1:0] y;
    input [width-1:0] in;
    assign y = $signed(in);
endmodule // ASSINT
module MulAddRecFN_postMul(
    input clock,
    input reset,
    input [2:0] io_fromPreMul_highExpA,
    input io_fromPreMul_isNaN_isQuietNaNA,
    input [2:0] io_fromPreMul_highExpB,
    input io_fromPreMul_isNaN_isQuietNaNB,
    input io_fromPreMul_signProd,
    input io_fromPreMul_isZeroProd,
    input io_fromPreMul_opSignC,
    input [2:0] io_fromPreMul_highExpC,
    input io_fromPreMul_isNaN_isQuietNaNC,
    input io_fromPreMul_isCDominant,
    input io_fromPreMul_CAlignDist_0,
    input [6:0] io_fromPreMul_CAlignDist,
    input io_fromPreMul_bit0AlignedNegSigC,
    input [25:0] io_fromPreMul_highAlignedNegSigC,
    input [10:0] io_fromPreMul_sExpSum,
    input [1:0] io_fromPreMul_roundingMode,
    input [48:0] io_mulAddResult,
    output [32:0] io_out,
    output [4:0] io_exceptionFlags
);
    wire isZeroA;
    wire [2:0] _WTEMP_92;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_729 (
        .y(_WTEMP_92),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(3)) u_eq_730 (
        .y(isZeroA),
        .a(io_fromPreMul_highExpA),
        .b(_WTEMP_92)
    );
    wire [1:0] _T_43;
    BITS #(.width(3), .high(2), .low(1)) bits_731 (
        .y(_T_43),
        .in(io_fromPreMul_highExpA)
    );
    wire isSpecialA;
    EQ_UNSIGNED #(.width(2)) u_eq_732 (
        .y(isSpecialA),
        .a(_T_43),
        .b(2'h3)
    );
    wire _T_45;
    BITS #(.width(3), .high(0), .low(0)) bits_733 (
        .y(_T_45),
        .in(io_fromPreMul_highExpA)
    );
    wire _T_47;
    EQ_UNSIGNED #(.width(1)) u_eq_734 (
        .y(_T_47),
        .a(_T_45),
        .b(1'h0)
    );
    wire isInfA;
    BITWISEAND #(.width(1)) bitwiseand_735 (
        .y(isInfA),
        .a(isSpecialA),
        .b(_T_47)
    );
    wire _T_48;
    BITS #(.width(3), .high(0), .low(0)) bits_736 (
        .y(_T_48),
        .in(io_fromPreMul_highExpA)
    );
    wire isNaNA;
    BITWISEAND #(.width(1)) bitwiseand_737 (
        .y(isNaNA),
        .a(isSpecialA),
        .b(_T_48)
    );
    wire _T_50;
    EQ_UNSIGNED #(.width(1)) u_eq_738 (
        .y(_T_50),
        .a(io_fromPreMul_isNaN_isQuietNaNA),
        .b(1'h0)
    );
    wire isSigNaNA;
    BITWISEAND #(.width(1)) bitwiseand_739 (
        .y(isSigNaNA),
        .a(isNaNA),
        .b(_T_50)
    );
    wire isZeroB;
    wire [2:0] _WTEMP_93;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_740 (
        .y(_WTEMP_93),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(3)) u_eq_741 (
        .y(isZeroB),
        .a(io_fromPreMul_highExpB),
        .b(_WTEMP_93)
    );
    wire [1:0] _T_52;
    BITS #(.width(3), .high(2), .low(1)) bits_742 (
        .y(_T_52),
        .in(io_fromPreMul_highExpB)
    );
    wire isSpecialB;
    EQ_UNSIGNED #(.width(2)) u_eq_743 (
        .y(isSpecialB),
        .a(_T_52),
        .b(2'h3)
    );
    wire _T_54;
    BITS #(.width(3), .high(0), .low(0)) bits_744 (
        .y(_T_54),
        .in(io_fromPreMul_highExpB)
    );
    wire _T_56;
    EQ_UNSIGNED #(.width(1)) u_eq_745 (
        .y(_T_56),
        .a(_T_54),
        .b(1'h0)
    );
    wire isInfB;
    BITWISEAND #(.width(1)) bitwiseand_746 (
        .y(isInfB),
        .a(isSpecialB),
        .b(_T_56)
    );
    wire _T_57;
    BITS #(.width(3), .high(0), .low(0)) bits_747 (
        .y(_T_57),
        .in(io_fromPreMul_highExpB)
    );
    wire isNaNB;
    BITWISEAND #(.width(1)) bitwiseand_748 (
        .y(isNaNB),
        .a(isSpecialB),
        .b(_T_57)
    );
    wire _T_59;
    EQ_UNSIGNED #(.width(1)) u_eq_749 (
        .y(_T_59),
        .a(io_fromPreMul_isNaN_isQuietNaNB),
        .b(1'h0)
    );
    wire isSigNaNB;
    BITWISEAND #(.width(1)) bitwiseand_750 (
        .y(isSigNaNB),
        .a(isNaNB),
        .b(_T_59)
    );
    wire isZeroC;
    wire [2:0] _WTEMP_94;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_751 (
        .y(_WTEMP_94),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(3)) u_eq_752 (
        .y(isZeroC),
        .a(io_fromPreMul_highExpC),
        .b(_WTEMP_94)
    );
    wire [1:0] _T_61;
    BITS #(.width(3), .high(2), .low(1)) bits_753 (
        .y(_T_61),
        .in(io_fromPreMul_highExpC)
    );
    wire isSpecialC;
    EQ_UNSIGNED #(.width(2)) u_eq_754 (
        .y(isSpecialC),
        .a(_T_61),
        .b(2'h3)
    );
    wire _T_63;
    BITS #(.width(3), .high(0), .low(0)) bits_755 (
        .y(_T_63),
        .in(io_fromPreMul_highExpC)
    );
    wire _T_65;
    EQ_UNSIGNED #(.width(1)) u_eq_756 (
        .y(_T_65),
        .a(_T_63),
        .b(1'h0)
    );
    wire isInfC;
    BITWISEAND #(.width(1)) bitwiseand_757 (
        .y(isInfC),
        .a(isSpecialC),
        .b(_T_65)
    );
    wire _T_66;
    BITS #(.width(3), .high(0), .low(0)) bits_758 (
        .y(_T_66),
        .in(io_fromPreMul_highExpC)
    );
    wire isNaNC;
    BITWISEAND #(.width(1)) bitwiseand_759 (
        .y(isNaNC),
        .a(isSpecialC),
        .b(_T_66)
    );
    wire _T_68;
    EQ_UNSIGNED #(.width(1)) u_eq_760 (
        .y(_T_68),
        .a(io_fromPreMul_isNaN_isQuietNaNC),
        .b(1'h0)
    );
    wire isSigNaNC;
    BITWISEAND #(.width(1)) bitwiseand_761 (
        .y(isSigNaNC),
        .a(isNaNC),
        .b(_T_68)
    );
    wire roundingMode_nearest_even;
    EQ_UNSIGNED #(.width(2)) u_eq_762 (
        .y(roundingMode_nearest_even),
        .a(io_fromPreMul_roundingMode),
        .b(2'h0)
    );
    wire roundingMode_minMag;
    EQ_UNSIGNED #(.width(2)) u_eq_763 (
        .y(roundingMode_minMag),
        .a(io_fromPreMul_roundingMode),
        .b(2'h1)
    );
    wire roundingMode_min;
    EQ_UNSIGNED #(.width(2)) u_eq_764 (
        .y(roundingMode_min),
        .a(io_fromPreMul_roundingMode),
        .b(2'h2)
    );
    wire roundingMode_max;
    EQ_UNSIGNED #(.width(2)) u_eq_765 (
        .y(roundingMode_max),
        .a(io_fromPreMul_roundingMode),
        .b(2'h3)
    );
    wire signZeroNotEqOpSigns;
    MUX_UNSIGNED #(.width(1)) u_mux_766 (
        .y(signZeroNotEqOpSigns),
        .sel(roundingMode_min),
        .a(1'h1),
        .b(1'h0)
    );
    wire doSubMags;
    BITWISEXOR #(.width(1)) bitwisexor_767 (
        .y(doSubMags),
        .a(io_fromPreMul_signProd),
        .b(io_fromPreMul_opSignC)
    );
    wire _T_71;
    BITS #(.width(49), .high(48), .low(48)) bits_768 (
        .y(_T_71),
        .in(io_mulAddResult)
    );
    wire [26:0] _T_73;
    wire [25:0] _WTEMP_95;
    PAD_UNSIGNED #(.width(1), .n(26)) u_pad_769 (
        .y(_WTEMP_95),
        .in(1'h1)
    );
    ADD_UNSIGNED #(.width(26)) u_add_770 (
        .y(_T_73),
        .a(io_fromPreMul_highAlignedNegSigC),
        .b(_WTEMP_95)
    );
    wire [25:0] _T_74;
    TAIL #(.width(27), .n(1)) tail_771 (
        .y(_T_74),
        .in(_T_73)
    );
    wire [25:0] _T_75;
    MUX_UNSIGNED #(.width(26)) u_mux_772 (
        .y(_T_75),
        .sel(_T_71),
        .a(_T_74),
        .b(io_fromPreMul_highAlignedNegSigC)
    );
    wire [47:0] _T_76;
    BITS #(.width(49), .high(47), .low(0)) bits_773 (
        .y(_T_76),
        .in(io_mulAddResult)
    );
    wire [73:0] _T_77;
    CAT #(.width_a(26), .width_b(48)) cat_774 (
        .y(_T_77),
        .a(_T_75),
        .b(_T_76)
    );
    wire [74:0] sigSum;
    CAT #(.width_a(74), .width_b(1)) cat_775 (
        .y(sigSum),
        .a(_T_77),
        .b(io_fromPreMul_bit0AlignedNegSigC)
    );
    wire [49:0] _T_79;
    BITS #(.width(75), .high(50), .low(1)) bits_776 (
        .y(_T_79),
        .in(sigSum)
    );
    wire [49:0] _T_80;
    BITWISEXOR #(.width(50)) bitwisexor_777 (
        .y(_T_80),
        .a(50'h0),
        .b(_T_79)
    );
    wire [49:0] _T_81;
    BITWISEOR #(.width(50)) bitwiseor_778 (
        .y(_T_81),
        .a(50'h0),
        .b(_T_79)
    );
    wire [50:0] _T_82;
    SHL_UNSIGNED #(.width(50), .n(1)) u_shl_779 (
        .y(_T_82),
        .in(_T_81)
    );
    wire [50:0] _T_83;
    wire [50:0] _WTEMP_96;
    PAD_UNSIGNED #(.width(50), .n(51)) u_pad_780 (
        .y(_WTEMP_96),
        .in(_T_80)
    );
    BITWISEXOR #(.width(51)) bitwisexor_781 (
        .y(_T_83),
        .a(_WTEMP_96),
        .b(_T_82)
    );
    wire [49:0] _T_85;
    BITS #(.width(51), .high(49), .low(0)) bits_782 (
        .y(_T_85),
        .in(_T_83)
    );
    wire [17:0] _T_86;
    BITS #(.width(50), .high(49), .low(32)) bits_783 (
        .y(_T_86),
        .in(_T_85)
    );
    wire [31:0] _T_87;
    BITS #(.width(50), .high(31), .low(0)) bits_784 (
        .y(_T_87),
        .in(_T_85)
    );
    wire _T_89;
    wire [17:0] _WTEMP_97;
    PAD_UNSIGNED #(.width(1), .n(18)) u_pad_785 (
        .y(_WTEMP_97),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(18)) u_neq_786 (
        .y(_T_89),
        .a(_T_86),
        .b(_WTEMP_97)
    );
    wire [1:0] _T_90;
    BITS #(.width(18), .high(17), .low(16)) bits_787 (
        .y(_T_90),
        .in(_T_86)
    );
    wire [15:0] _T_91;
    BITS #(.width(18), .high(15), .low(0)) bits_788 (
        .y(_T_91),
        .in(_T_86)
    );
    wire _T_93;
    wire [1:0] _WTEMP_98;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_789 (
        .y(_WTEMP_98),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(2)) u_neq_790 (
        .y(_T_93),
        .a(_T_90),
        .b(_WTEMP_98)
    );
    wire _T_94;
    BITS #(.width(2), .high(1), .low(1)) bits_791 (
        .y(_T_94),
        .in(_T_90)
    );
    wire [7:0] _T_95;
    BITS #(.width(16), .high(15), .low(8)) bits_792 (
        .y(_T_95),
        .in(_T_91)
    );
    wire [7:0] _T_96;
    BITS #(.width(16), .high(7), .low(0)) bits_793 (
        .y(_T_96),
        .in(_T_91)
    );
    wire _T_98;
    wire [7:0] _WTEMP_99;
    PAD_UNSIGNED #(.width(1), .n(8)) u_pad_794 (
        .y(_WTEMP_99),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(8)) u_neq_795 (
        .y(_T_98),
        .a(_T_95),
        .b(_WTEMP_99)
    );
    wire [3:0] _T_99;
    BITS #(.width(8), .high(7), .low(4)) bits_796 (
        .y(_T_99),
        .in(_T_95)
    );
    wire [3:0] _T_100;
    BITS #(.width(8), .high(3), .low(0)) bits_797 (
        .y(_T_100),
        .in(_T_95)
    );
    wire _T_102;
    wire [3:0] _WTEMP_100;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_798 (
        .y(_WTEMP_100),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_799 (
        .y(_T_102),
        .a(_T_99),
        .b(_WTEMP_100)
    );
    wire _T_103;
    BITS #(.width(4), .high(3), .low(3)) bits_800 (
        .y(_T_103),
        .in(_T_99)
    );
    wire _T_105;
    BITS #(.width(4), .high(2), .low(2)) bits_801 (
        .y(_T_105),
        .in(_T_99)
    );
    wire _T_107;
    BITS #(.width(4), .high(1), .low(1)) bits_802 (
        .y(_T_107),
        .in(_T_99)
    );
    wire [1:0] _T_108;
    wire [1:0] _WTEMP_101;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_803 (
        .y(_WTEMP_101),
        .in(_T_107)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_804 (
        .y(_T_108),
        .sel(_T_105),
        .a(2'h2),
        .b(_WTEMP_101)
    );
    wire [1:0] _T_109;
    MUX_UNSIGNED #(.width(2)) u_mux_805 (
        .y(_T_109),
        .sel(_T_103),
        .a(2'h3),
        .b(_T_108)
    );
    wire _T_110;
    BITS #(.width(4), .high(3), .low(3)) bits_806 (
        .y(_T_110),
        .in(_T_100)
    );
    wire _T_112;
    BITS #(.width(4), .high(2), .low(2)) bits_807 (
        .y(_T_112),
        .in(_T_100)
    );
    wire _T_114;
    BITS #(.width(4), .high(1), .low(1)) bits_808 (
        .y(_T_114),
        .in(_T_100)
    );
    wire [1:0] _T_115;
    wire [1:0] _WTEMP_102;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_809 (
        .y(_WTEMP_102),
        .in(_T_114)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_810 (
        .y(_T_115),
        .sel(_T_112),
        .a(2'h2),
        .b(_WTEMP_102)
    );
    wire [1:0] _T_116;
    MUX_UNSIGNED #(.width(2)) u_mux_811 (
        .y(_T_116),
        .sel(_T_110),
        .a(2'h3),
        .b(_T_115)
    );
    wire [1:0] _T_117;
    MUX_UNSIGNED #(.width(2)) u_mux_812 (
        .y(_T_117),
        .sel(_T_102),
        .a(_T_109),
        .b(_T_116)
    );
    wire [2:0] _T_118;
    CAT #(.width_a(1), .width_b(2)) cat_813 (
        .y(_T_118),
        .a(_T_102),
        .b(_T_117)
    );
    wire [3:0] _T_119;
    BITS #(.width(8), .high(7), .low(4)) bits_814 (
        .y(_T_119),
        .in(_T_96)
    );
    wire [3:0] _T_120;
    BITS #(.width(8), .high(3), .low(0)) bits_815 (
        .y(_T_120),
        .in(_T_96)
    );
    wire _T_122;
    wire [3:0] _WTEMP_103;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_816 (
        .y(_WTEMP_103),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_817 (
        .y(_T_122),
        .a(_T_119),
        .b(_WTEMP_103)
    );
    wire _T_123;
    BITS #(.width(4), .high(3), .low(3)) bits_818 (
        .y(_T_123),
        .in(_T_119)
    );
    wire _T_125;
    BITS #(.width(4), .high(2), .low(2)) bits_819 (
        .y(_T_125),
        .in(_T_119)
    );
    wire _T_127;
    BITS #(.width(4), .high(1), .low(1)) bits_820 (
        .y(_T_127),
        .in(_T_119)
    );
    wire [1:0] _T_128;
    wire [1:0] _WTEMP_104;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_821 (
        .y(_WTEMP_104),
        .in(_T_127)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_822 (
        .y(_T_128),
        .sel(_T_125),
        .a(2'h2),
        .b(_WTEMP_104)
    );
    wire [1:0] _T_129;
    MUX_UNSIGNED #(.width(2)) u_mux_823 (
        .y(_T_129),
        .sel(_T_123),
        .a(2'h3),
        .b(_T_128)
    );
    wire _T_130;
    BITS #(.width(4), .high(3), .low(3)) bits_824 (
        .y(_T_130),
        .in(_T_120)
    );
    wire _T_132;
    BITS #(.width(4), .high(2), .low(2)) bits_825 (
        .y(_T_132),
        .in(_T_120)
    );
    wire _T_134;
    BITS #(.width(4), .high(1), .low(1)) bits_826 (
        .y(_T_134),
        .in(_T_120)
    );
    wire [1:0] _T_135;
    wire [1:0] _WTEMP_105;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_827 (
        .y(_WTEMP_105),
        .in(_T_134)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_828 (
        .y(_T_135),
        .sel(_T_132),
        .a(2'h2),
        .b(_WTEMP_105)
    );
    wire [1:0] _T_136;
    MUX_UNSIGNED #(.width(2)) u_mux_829 (
        .y(_T_136),
        .sel(_T_130),
        .a(2'h3),
        .b(_T_135)
    );
    wire [1:0] _T_137;
    MUX_UNSIGNED #(.width(2)) u_mux_830 (
        .y(_T_137),
        .sel(_T_122),
        .a(_T_129),
        .b(_T_136)
    );
    wire [2:0] _T_138;
    CAT #(.width_a(1), .width_b(2)) cat_831 (
        .y(_T_138),
        .a(_T_122),
        .b(_T_137)
    );
    wire [2:0] _T_139;
    MUX_UNSIGNED #(.width(3)) u_mux_832 (
        .y(_T_139),
        .sel(_T_98),
        .a(_T_118),
        .b(_T_138)
    );
    wire [3:0] _T_140;
    CAT #(.width_a(1), .width_b(3)) cat_833 (
        .y(_T_140),
        .a(_T_98),
        .b(_T_139)
    );
    wire [3:0] _T_141;
    wire [3:0] _WTEMP_106;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_834 (
        .y(_WTEMP_106),
        .in(_T_94)
    );
    MUX_UNSIGNED #(.width(4)) u_mux_835 (
        .y(_T_141),
        .sel(_T_93),
        .a(_WTEMP_106),
        .b(_T_140)
    );
    wire [4:0] _T_142;
    CAT #(.width_a(1), .width_b(4)) cat_836 (
        .y(_T_142),
        .a(_T_93),
        .b(_T_141)
    );
    wire [15:0] _T_143;
    BITS #(.width(32), .high(31), .low(16)) bits_837 (
        .y(_T_143),
        .in(_T_87)
    );
    wire [15:0] _T_144;
    BITS #(.width(32), .high(15), .low(0)) bits_838 (
        .y(_T_144),
        .in(_T_87)
    );
    wire _T_146;
    wire [15:0] _WTEMP_107;
    PAD_UNSIGNED #(.width(1), .n(16)) u_pad_839 (
        .y(_WTEMP_107),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(16)) u_neq_840 (
        .y(_T_146),
        .a(_T_143),
        .b(_WTEMP_107)
    );
    wire [7:0] _T_147;
    BITS #(.width(16), .high(15), .low(8)) bits_841 (
        .y(_T_147),
        .in(_T_143)
    );
    wire [7:0] _T_148;
    BITS #(.width(16), .high(7), .low(0)) bits_842 (
        .y(_T_148),
        .in(_T_143)
    );
    wire _T_150;
    wire [7:0] _WTEMP_108;
    PAD_UNSIGNED #(.width(1), .n(8)) u_pad_843 (
        .y(_WTEMP_108),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(8)) u_neq_844 (
        .y(_T_150),
        .a(_T_147),
        .b(_WTEMP_108)
    );
    wire [3:0] _T_151;
    BITS #(.width(8), .high(7), .low(4)) bits_845 (
        .y(_T_151),
        .in(_T_147)
    );
    wire [3:0] _T_152;
    BITS #(.width(8), .high(3), .low(0)) bits_846 (
        .y(_T_152),
        .in(_T_147)
    );
    wire _T_154;
    wire [3:0] _WTEMP_109;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_847 (
        .y(_WTEMP_109),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_848 (
        .y(_T_154),
        .a(_T_151),
        .b(_WTEMP_109)
    );
    wire _T_155;
    BITS #(.width(4), .high(3), .low(3)) bits_849 (
        .y(_T_155),
        .in(_T_151)
    );
    wire _T_157;
    BITS #(.width(4), .high(2), .low(2)) bits_850 (
        .y(_T_157),
        .in(_T_151)
    );
    wire _T_159;
    BITS #(.width(4), .high(1), .low(1)) bits_851 (
        .y(_T_159),
        .in(_T_151)
    );
    wire [1:0] _T_160;
    wire [1:0] _WTEMP_110;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_852 (
        .y(_WTEMP_110),
        .in(_T_159)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_853 (
        .y(_T_160),
        .sel(_T_157),
        .a(2'h2),
        .b(_WTEMP_110)
    );
    wire [1:0] _T_161;
    MUX_UNSIGNED #(.width(2)) u_mux_854 (
        .y(_T_161),
        .sel(_T_155),
        .a(2'h3),
        .b(_T_160)
    );
    wire _T_162;
    BITS #(.width(4), .high(3), .low(3)) bits_855 (
        .y(_T_162),
        .in(_T_152)
    );
    wire _T_164;
    BITS #(.width(4), .high(2), .low(2)) bits_856 (
        .y(_T_164),
        .in(_T_152)
    );
    wire _T_166;
    BITS #(.width(4), .high(1), .low(1)) bits_857 (
        .y(_T_166),
        .in(_T_152)
    );
    wire [1:0] _T_167;
    wire [1:0] _WTEMP_111;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_858 (
        .y(_WTEMP_111),
        .in(_T_166)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_859 (
        .y(_T_167),
        .sel(_T_164),
        .a(2'h2),
        .b(_WTEMP_111)
    );
    wire [1:0] _T_168;
    MUX_UNSIGNED #(.width(2)) u_mux_860 (
        .y(_T_168),
        .sel(_T_162),
        .a(2'h3),
        .b(_T_167)
    );
    wire [1:0] _T_169;
    MUX_UNSIGNED #(.width(2)) u_mux_861 (
        .y(_T_169),
        .sel(_T_154),
        .a(_T_161),
        .b(_T_168)
    );
    wire [2:0] _T_170;
    CAT #(.width_a(1), .width_b(2)) cat_862 (
        .y(_T_170),
        .a(_T_154),
        .b(_T_169)
    );
    wire [3:0] _T_171;
    BITS #(.width(8), .high(7), .low(4)) bits_863 (
        .y(_T_171),
        .in(_T_148)
    );
    wire [3:0] _T_172;
    BITS #(.width(8), .high(3), .low(0)) bits_864 (
        .y(_T_172),
        .in(_T_148)
    );
    wire _T_174;
    wire [3:0] _WTEMP_112;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_865 (
        .y(_WTEMP_112),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_866 (
        .y(_T_174),
        .a(_T_171),
        .b(_WTEMP_112)
    );
    wire _T_175;
    BITS #(.width(4), .high(3), .low(3)) bits_867 (
        .y(_T_175),
        .in(_T_171)
    );
    wire _T_177;
    BITS #(.width(4), .high(2), .low(2)) bits_868 (
        .y(_T_177),
        .in(_T_171)
    );
    wire _T_179;
    BITS #(.width(4), .high(1), .low(1)) bits_869 (
        .y(_T_179),
        .in(_T_171)
    );
    wire [1:0] _T_180;
    wire [1:0] _WTEMP_113;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_870 (
        .y(_WTEMP_113),
        .in(_T_179)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_871 (
        .y(_T_180),
        .sel(_T_177),
        .a(2'h2),
        .b(_WTEMP_113)
    );
    wire [1:0] _T_181;
    MUX_UNSIGNED #(.width(2)) u_mux_872 (
        .y(_T_181),
        .sel(_T_175),
        .a(2'h3),
        .b(_T_180)
    );
    wire _T_182;
    BITS #(.width(4), .high(3), .low(3)) bits_873 (
        .y(_T_182),
        .in(_T_172)
    );
    wire _T_184;
    BITS #(.width(4), .high(2), .low(2)) bits_874 (
        .y(_T_184),
        .in(_T_172)
    );
    wire _T_186;
    BITS #(.width(4), .high(1), .low(1)) bits_875 (
        .y(_T_186),
        .in(_T_172)
    );
    wire [1:0] _T_187;
    wire [1:0] _WTEMP_114;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_876 (
        .y(_WTEMP_114),
        .in(_T_186)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_877 (
        .y(_T_187),
        .sel(_T_184),
        .a(2'h2),
        .b(_WTEMP_114)
    );
    wire [1:0] _T_188;
    MUX_UNSIGNED #(.width(2)) u_mux_878 (
        .y(_T_188),
        .sel(_T_182),
        .a(2'h3),
        .b(_T_187)
    );
    wire [1:0] _T_189;
    MUX_UNSIGNED #(.width(2)) u_mux_879 (
        .y(_T_189),
        .sel(_T_174),
        .a(_T_181),
        .b(_T_188)
    );
    wire [2:0] _T_190;
    CAT #(.width_a(1), .width_b(2)) cat_880 (
        .y(_T_190),
        .a(_T_174),
        .b(_T_189)
    );
    wire [2:0] _T_191;
    MUX_UNSIGNED #(.width(3)) u_mux_881 (
        .y(_T_191),
        .sel(_T_150),
        .a(_T_170),
        .b(_T_190)
    );
    wire [3:0] _T_192;
    CAT #(.width_a(1), .width_b(3)) cat_882 (
        .y(_T_192),
        .a(_T_150),
        .b(_T_191)
    );
    wire [7:0] _T_193;
    BITS #(.width(16), .high(15), .low(8)) bits_883 (
        .y(_T_193),
        .in(_T_144)
    );
    wire [7:0] _T_194;
    BITS #(.width(16), .high(7), .low(0)) bits_884 (
        .y(_T_194),
        .in(_T_144)
    );
    wire _T_196;
    wire [7:0] _WTEMP_115;
    PAD_UNSIGNED #(.width(1), .n(8)) u_pad_885 (
        .y(_WTEMP_115),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(8)) u_neq_886 (
        .y(_T_196),
        .a(_T_193),
        .b(_WTEMP_115)
    );
    wire [3:0] _T_197;
    BITS #(.width(8), .high(7), .low(4)) bits_887 (
        .y(_T_197),
        .in(_T_193)
    );
    wire [3:0] _T_198;
    BITS #(.width(8), .high(3), .low(0)) bits_888 (
        .y(_T_198),
        .in(_T_193)
    );
    wire _T_200;
    wire [3:0] _WTEMP_116;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_889 (
        .y(_WTEMP_116),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_890 (
        .y(_T_200),
        .a(_T_197),
        .b(_WTEMP_116)
    );
    wire _T_201;
    BITS #(.width(4), .high(3), .low(3)) bits_891 (
        .y(_T_201),
        .in(_T_197)
    );
    wire _T_203;
    BITS #(.width(4), .high(2), .low(2)) bits_892 (
        .y(_T_203),
        .in(_T_197)
    );
    wire _T_205;
    BITS #(.width(4), .high(1), .low(1)) bits_893 (
        .y(_T_205),
        .in(_T_197)
    );
    wire [1:0] _T_206;
    wire [1:0] _WTEMP_117;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_894 (
        .y(_WTEMP_117),
        .in(_T_205)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_895 (
        .y(_T_206),
        .sel(_T_203),
        .a(2'h2),
        .b(_WTEMP_117)
    );
    wire [1:0] _T_207;
    MUX_UNSIGNED #(.width(2)) u_mux_896 (
        .y(_T_207),
        .sel(_T_201),
        .a(2'h3),
        .b(_T_206)
    );
    wire _T_208;
    BITS #(.width(4), .high(3), .low(3)) bits_897 (
        .y(_T_208),
        .in(_T_198)
    );
    wire _T_210;
    BITS #(.width(4), .high(2), .low(2)) bits_898 (
        .y(_T_210),
        .in(_T_198)
    );
    wire _T_212;
    BITS #(.width(4), .high(1), .low(1)) bits_899 (
        .y(_T_212),
        .in(_T_198)
    );
    wire [1:0] _T_213;
    wire [1:0] _WTEMP_118;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_900 (
        .y(_WTEMP_118),
        .in(_T_212)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_901 (
        .y(_T_213),
        .sel(_T_210),
        .a(2'h2),
        .b(_WTEMP_118)
    );
    wire [1:0] _T_214;
    MUX_UNSIGNED #(.width(2)) u_mux_902 (
        .y(_T_214),
        .sel(_T_208),
        .a(2'h3),
        .b(_T_213)
    );
    wire [1:0] _T_215;
    MUX_UNSIGNED #(.width(2)) u_mux_903 (
        .y(_T_215),
        .sel(_T_200),
        .a(_T_207),
        .b(_T_214)
    );
    wire [2:0] _T_216;
    CAT #(.width_a(1), .width_b(2)) cat_904 (
        .y(_T_216),
        .a(_T_200),
        .b(_T_215)
    );
    wire [3:0] _T_217;
    BITS #(.width(8), .high(7), .low(4)) bits_905 (
        .y(_T_217),
        .in(_T_194)
    );
    wire [3:0] _T_218;
    BITS #(.width(8), .high(3), .low(0)) bits_906 (
        .y(_T_218),
        .in(_T_194)
    );
    wire _T_220;
    wire [3:0] _WTEMP_119;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_907 (
        .y(_WTEMP_119),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_908 (
        .y(_T_220),
        .a(_T_217),
        .b(_WTEMP_119)
    );
    wire _T_221;
    BITS #(.width(4), .high(3), .low(3)) bits_909 (
        .y(_T_221),
        .in(_T_217)
    );
    wire _T_223;
    BITS #(.width(4), .high(2), .low(2)) bits_910 (
        .y(_T_223),
        .in(_T_217)
    );
    wire _T_225;
    BITS #(.width(4), .high(1), .low(1)) bits_911 (
        .y(_T_225),
        .in(_T_217)
    );
    wire [1:0] _T_226;
    wire [1:0] _WTEMP_120;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_912 (
        .y(_WTEMP_120),
        .in(_T_225)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_913 (
        .y(_T_226),
        .sel(_T_223),
        .a(2'h2),
        .b(_WTEMP_120)
    );
    wire [1:0] _T_227;
    MUX_UNSIGNED #(.width(2)) u_mux_914 (
        .y(_T_227),
        .sel(_T_221),
        .a(2'h3),
        .b(_T_226)
    );
    wire _T_228;
    BITS #(.width(4), .high(3), .low(3)) bits_915 (
        .y(_T_228),
        .in(_T_218)
    );
    wire _T_230;
    BITS #(.width(4), .high(2), .low(2)) bits_916 (
        .y(_T_230),
        .in(_T_218)
    );
    wire _T_232;
    BITS #(.width(4), .high(1), .low(1)) bits_917 (
        .y(_T_232),
        .in(_T_218)
    );
    wire [1:0] _T_233;
    wire [1:0] _WTEMP_121;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_918 (
        .y(_WTEMP_121),
        .in(_T_232)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_919 (
        .y(_T_233),
        .sel(_T_230),
        .a(2'h2),
        .b(_WTEMP_121)
    );
    wire [1:0] _T_234;
    MUX_UNSIGNED #(.width(2)) u_mux_920 (
        .y(_T_234),
        .sel(_T_228),
        .a(2'h3),
        .b(_T_233)
    );
    wire [1:0] _T_235;
    MUX_UNSIGNED #(.width(2)) u_mux_921 (
        .y(_T_235),
        .sel(_T_220),
        .a(_T_227),
        .b(_T_234)
    );
    wire [2:0] _T_236;
    CAT #(.width_a(1), .width_b(2)) cat_922 (
        .y(_T_236),
        .a(_T_220),
        .b(_T_235)
    );
    wire [2:0] _T_237;
    MUX_UNSIGNED #(.width(3)) u_mux_923 (
        .y(_T_237),
        .sel(_T_196),
        .a(_T_216),
        .b(_T_236)
    );
    wire [3:0] _T_238;
    CAT #(.width_a(1), .width_b(3)) cat_924 (
        .y(_T_238),
        .a(_T_196),
        .b(_T_237)
    );
    wire [3:0] _T_239;
    MUX_UNSIGNED #(.width(4)) u_mux_925 (
        .y(_T_239),
        .sel(_T_146),
        .a(_T_192),
        .b(_T_238)
    );
    wire [4:0] _T_240;
    CAT #(.width_a(1), .width_b(4)) cat_926 (
        .y(_T_240),
        .a(_T_146),
        .b(_T_239)
    );
    wire [4:0] _T_241;
    MUX_UNSIGNED #(.width(5)) u_mux_927 (
        .y(_T_241),
        .sel(_T_89),
        .a(_T_142),
        .b(_T_240)
    );
    wire [5:0] _T_242;
    CAT #(.width_a(1), .width_b(5)) cat_928 (
        .y(_T_242),
        .a(_T_89),
        .b(_T_241)
    );
    wire [7:0] _T_243;
    wire [6:0] _WTEMP_122;
    PAD_UNSIGNED #(.width(6), .n(7)) u_pad_929 (
        .y(_WTEMP_122),
        .in(_T_242)
    );
    SUB_UNSIGNED #(.width(7)) u_sub_930 (
        .y(_T_243),
        .a(7'h49),
        .b(_WTEMP_122)
    );
    wire [7:0] _T_244;
    ASUINT #(.width(8)) asuint_931 (
        .y(_T_244),
        .in(_T_243)
    );
    wire [6:0] estNormNeg_dist;
    TAIL #(.width(8), .n(1)) tail_932 (
        .y(estNormNeg_dist),
        .in(_T_244)
    );
    wire [15:0] _T_245;
    BITS #(.width(75), .high(33), .low(18)) bits_933 (
        .y(_T_245),
        .in(sigSum)
    );
    wire _T_247;
    wire [15:0] _WTEMP_123;
    PAD_UNSIGNED #(.width(1), .n(16)) u_pad_934 (
        .y(_WTEMP_123),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(16)) u_neq_935 (
        .y(_T_247),
        .a(_T_245),
        .b(_WTEMP_123)
    );
    wire [17:0] _T_248;
    BITS #(.width(75), .high(17), .low(0)) bits_936 (
        .y(_T_248),
        .in(sigSum)
    );
    wire _T_250;
    wire [17:0] _WTEMP_124;
    PAD_UNSIGNED #(.width(1), .n(18)) u_pad_937 (
        .y(_WTEMP_124),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(18)) u_neq_938 (
        .y(_T_250),
        .a(_T_248),
        .b(_WTEMP_124)
    );
    wire [1:0] firstReduceSigSum;
    CAT #(.width_a(1), .width_b(1)) cat_939 (
        .y(firstReduceSigSum),
        .a(_T_247),
        .b(_T_250)
    );
    wire [74:0] complSigSum;
    BITWISENOT #(.width(75)) bitwisenot_940 (
        .y(complSigSum),
        .in(sigSum)
    );
    wire [15:0] _T_251;
    BITS #(.width(75), .high(33), .low(18)) bits_941 (
        .y(_T_251),
        .in(complSigSum)
    );
    wire _T_253;
    wire [15:0] _WTEMP_125;
    PAD_UNSIGNED #(.width(1), .n(16)) u_pad_942 (
        .y(_WTEMP_125),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(16)) u_neq_943 (
        .y(_T_253),
        .a(_T_251),
        .b(_WTEMP_125)
    );
    wire [17:0] _T_254;
    BITS #(.width(75), .high(17), .low(0)) bits_944 (
        .y(_T_254),
        .in(complSigSum)
    );
    wire _T_256;
    wire [17:0] _WTEMP_126;
    PAD_UNSIGNED #(.width(1), .n(18)) u_pad_945 (
        .y(_WTEMP_126),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(18)) u_neq_946 (
        .y(_T_256),
        .a(_T_254),
        .b(_WTEMP_126)
    );
    wire [1:0] firstReduceComplSigSum;
    CAT #(.width_a(1), .width_b(1)) cat_947 (
        .y(firstReduceComplSigSum),
        .a(_T_253),
        .b(_T_256)
    );
    wire _T_257;
    BITWISEOR #(.width(1)) bitwiseor_948 (
        .y(_T_257),
        .a(io_fromPreMul_CAlignDist_0),
        .b(doSubMags)
    );
    wire [7:0] _T_259;
    wire [6:0] _WTEMP_127;
    PAD_UNSIGNED #(.width(1), .n(7)) u_pad_949 (
        .y(_WTEMP_127),
        .in(1'h1)
    );
    SUB_UNSIGNED #(.width(7)) u_sub_950 (
        .y(_T_259),
        .a(io_fromPreMul_CAlignDist),
        .b(_WTEMP_127)
    );
    wire [7:0] _T_260;
    ASUINT #(.width(8)) asuint_951 (
        .y(_T_260),
        .in(_T_259)
    );
    wire [6:0] _T_261;
    TAIL #(.width(8), .n(1)) tail_952 (
        .y(_T_261),
        .in(_T_260)
    );
    wire [4:0] _T_262;
    BITS #(.width(7), .high(4), .low(0)) bits_953 (
        .y(_T_262),
        .in(_T_261)
    );
    wire [6:0] CDom_estNormDist;
    wire [6:0] _WTEMP_128;
    PAD_UNSIGNED #(.width(5), .n(7)) u_pad_954 (
        .y(_WTEMP_128),
        .in(_T_262)
    );
    MUX_UNSIGNED #(.width(7)) u_mux_955 (
        .y(CDom_estNormDist),
        .sel(_T_257),
        .a(io_fromPreMul_CAlignDist),
        .b(_WTEMP_128)
    );
    wire _T_264;
    EQ_UNSIGNED #(.width(1)) u_eq_956 (
        .y(_T_264),
        .a(doSubMags),
        .b(1'h0)
    );
    wire _T_265;
    BITS #(.width(7), .high(4), .low(4)) bits_957 (
        .y(_T_265),
        .in(CDom_estNormDist)
    );
    wire _T_267;
    EQ_UNSIGNED #(.width(1)) u_eq_958 (
        .y(_T_267),
        .a(_T_265),
        .b(1'h0)
    );
    wire _T_268;
    BITWISEAND #(.width(1)) bitwiseand_959 (
        .y(_T_268),
        .a(_T_264),
        .b(_T_267)
    );
    wire [40:0] _T_269;
    BITS #(.width(75), .high(74), .low(34)) bits_960 (
        .y(_T_269),
        .in(sigSum)
    );
    wire _T_271;
    wire [1:0] _WTEMP_129;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_961 (
        .y(_WTEMP_129),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(2)) u_neq_962 (
        .y(_T_271),
        .a(firstReduceSigSum),
        .b(_WTEMP_129)
    );
    wire [41:0] _T_272;
    CAT #(.width_a(41), .width_b(1)) cat_963 (
        .y(_T_272),
        .a(_T_269),
        .b(_T_271)
    );
    wire [41:0] _T_274;
    wire [41:0] _WTEMP_130;
    PAD_UNSIGNED #(.width(1), .n(42)) u_pad_964 (
        .y(_WTEMP_130),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(42)) u_mux_965 (
        .y(_T_274),
        .sel(_T_268),
        .a(_T_272),
        .b(_WTEMP_130)
    );
    wire _T_276;
    EQ_UNSIGNED #(.width(1)) u_eq_966 (
        .y(_T_276),
        .a(doSubMags),
        .b(1'h0)
    );
    wire _T_277;
    BITS #(.width(7), .high(4), .low(4)) bits_967 (
        .y(_T_277),
        .in(CDom_estNormDist)
    );
    wire _T_278;
    BITWISEAND #(.width(1)) bitwiseand_968 (
        .y(_T_278),
        .a(_T_276),
        .b(_T_277)
    );
    wire [40:0] _T_279;
    BITS #(.width(75), .high(58), .low(18)) bits_969 (
        .y(_T_279),
        .in(sigSum)
    );
    wire _T_280;
    BITS #(.width(2), .high(0), .low(0)) bits_970 (
        .y(_T_280),
        .in(firstReduceSigSum)
    );
    wire [41:0] _T_281;
    CAT #(.width_a(41), .width_b(1)) cat_971 (
        .y(_T_281),
        .a(_T_279),
        .b(_T_280)
    );
    wire [41:0] _T_283;
    wire [41:0] _WTEMP_131;
    PAD_UNSIGNED #(.width(1), .n(42)) u_pad_972 (
        .y(_WTEMP_131),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(42)) u_mux_973 (
        .y(_T_283),
        .sel(_T_278),
        .a(_T_281),
        .b(_WTEMP_131)
    );
    wire [41:0] _T_284;
    BITWISEOR #(.width(42)) bitwiseor_974 (
        .y(_T_284),
        .a(_T_274),
        .b(_T_283)
    );
    wire _T_285;
    BITS #(.width(7), .high(4), .low(4)) bits_975 (
        .y(_T_285),
        .in(CDom_estNormDist)
    );
    wire _T_287;
    EQ_UNSIGNED #(.width(1)) u_eq_976 (
        .y(_T_287),
        .a(_T_285),
        .b(1'h0)
    );
    wire _T_288;
    BITWISEAND #(.width(1)) bitwiseand_977 (
        .y(_T_288),
        .a(doSubMags),
        .b(_T_287)
    );
    wire [40:0] _T_289;
    BITS #(.width(75), .high(74), .low(34)) bits_978 (
        .y(_T_289),
        .in(complSigSum)
    );
    wire _T_291;
    wire [1:0] _WTEMP_132;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_979 (
        .y(_WTEMP_132),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(2)) u_neq_980 (
        .y(_T_291),
        .a(firstReduceComplSigSum),
        .b(_WTEMP_132)
    );
    wire [41:0] _T_292;
    CAT #(.width_a(41), .width_b(1)) cat_981 (
        .y(_T_292),
        .a(_T_289),
        .b(_T_291)
    );
    wire [41:0] _T_294;
    wire [41:0] _WTEMP_133;
    PAD_UNSIGNED #(.width(1), .n(42)) u_pad_982 (
        .y(_WTEMP_133),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(42)) u_mux_983 (
        .y(_T_294),
        .sel(_T_288),
        .a(_T_292),
        .b(_WTEMP_133)
    );
    wire [41:0] _T_295;
    BITWISEOR #(.width(42)) bitwiseor_984 (
        .y(_T_295),
        .a(_T_284),
        .b(_T_294)
    );
    wire _T_296;
    BITS #(.width(7), .high(4), .low(4)) bits_985 (
        .y(_T_296),
        .in(CDom_estNormDist)
    );
    wire _T_297;
    BITWISEAND #(.width(1)) bitwiseand_986 (
        .y(_T_297),
        .a(doSubMags),
        .b(_T_296)
    );
    wire [40:0] _T_298;
    BITS #(.width(75), .high(58), .low(18)) bits_987 (
        .y(_T_298),
        .in(complSigSum)
    );
    wire _T_299;
    BITS #(.width(2), .high(0), .low(0)) bits_988 (
        .y(_T_299),
        .in(firstReduceComplSigSum)
    );
    wire [41:0] _T_300;
    CAT #(.width_a(41), .width_b(1)) cat_989 (
        .y(_T_300),
        .a(_T_298),
        .b(_T_299)
    );
    wire [41:0] _T_302;
    wire [41:0] _WTEMP_134;
    PAD_UNSIGNED #(.width(1), .n(42)) u_pad_990 (
        .y(_WTEMP_134),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(42)) u_mux_991 (
        .y(_T_302),
        .sel(_T_297),
        .a(_T_300),
        .b(_WTEMP_134)
    );
    wire [41:0] CDom_firstNormAbsSigSum;
    BITWISEOR #(.width(42)) bitwiseor_992 (
        .y(CDom_firstNormAbsSigSum),
        .a(_T_295),
        .b(_T_302)
    );
    wire [32:0] _T_303;
    BITS #(.width(75), .high(50), .low(18)) bits_993 (
        .y(_T_303),
        .in(sigSum)
    );
    wire _T_304;
    BITS #(.width(2), .high(0), .low(0)) bits_994 (
        .y(_T_304),
        .in(firstReduceComplSigSum)
    );
    wire _T_306;
    EQ_UNSIGNED #(.width(1)) u_eq_995 (
        .y(_T_306),
        .a(_T_304),
        .b(1'h0)
    );
    wire _T_307;
    BITS #(.width(2), .high(0), .low(0)) bits_996 (
        .y(_T_307),
        .in(firstReduceSigSum)
    );
    wire _T_308;
    MUX_UNSIGNED #(.width(1)) u_mux_997 (
        .y(_T_308),
        .sel(doSubMags),
        .a(_T_306),
        .b(_T_307)
    );
    wire [33:0] _T_309;
    CAT #(.width_a(33), .width_b(1)) cat_998 (
        .y(_T_309),
        .a(_T_303),
        .b(_T_308)
    );
    wire [41:0] _T_310;
    BITS #(.width(75), .high(42), .low(1)) bits_999 (
        .y(_T_310),
        .in(sigSum)
    );
    wire _T_311;
    BITS #(.width(7), .high(5), .low(5)) bits_1000 (
        .y(_T_311),
        .in(estNormNeg_dist)
    );
    wire _T_312;
    BITS #(.width(7), .high(4), .low(4)) bits_1001 (
        .y(_T_312),
        .in(estNormNeg_dist)
    );
    wire [25:0] _T_313;
    BITS #(.width(75), .high(26), .low(1)) bits_1002 (
        .y(_T_313),
        .in(sigSum)
    );
    wire _T_314;
    BITS #(.width(1), .high(0), .low(0)) bits_1003 (
        .y(_T_314),
        .in(doSubMags)
    );
    wire [15:0] _T_317;
    MUX_UNSIGNED #(.width(16)) u_mux_1004 (
        .y(_T_317),
        .sel(_T_314),
        .a(16'hFFFF),
        .b(16'h0)
    );
    wire [41:0] _T_318;
    CAT #(.width_a(26), .width_b(16)) cat_1005 (
        .y(_T_318),
        .a(_T_313),
        .b(_T_317)
    );
    wire [41:0] _T_319;
    MUX_UNSIGNED #(.width(42)) u_mux_1006 (
        .y(_T_319),
        .sel(_T_312),
        .a(_T_318),
        .b(_T_310)
    );
    wire _T_320;
    BITS #(.width(7), .high(4), .low(4)) bits_1007 (
        .y(_T_320),
        .in(estNormNeg_dist)
    );
    wire [9:0] _T_321;
    BITS #(.width(75), .high(10), .low(1)) bits_1008 (
        .y(_T_321),
        .in(sigSum)
    );
    wire _T_322;
    BITS #(.width(1), .high(0), .low(0)) bits_1009 (
        .y(_T_322),
        .in(doSubMags)
    );
    wire [31:0] _T_325;
    MUX_UNSIGNED #(.width(32)) u_mux_1010 (
        .y(_T_325),
        .sel(_T_322),
        .a(32'hFFFFFFFF),
        .b(32'h0)
    );
    wire [41:0] _T_326;
    CAT #(.width_a(10), .width_b(32)) cat_1011 (
        .y(_T_326),
        .a(_T_321),
        .b(_T_325)
    );
    wire [41:0] _T_327;
    wire [41:0] _WTEMP_135;
    PAD_UNSIGNED #(.width(34), .n(42)) u_pad_1012 (
        .y(_WTEMP_135),
        .in(_T_309)
    );
    MUX_UNSIGNED #(.width(42)) u_mux_1013 (
        .y(_T_327),
        .sel(_T_320),
        .a(_WTEMP_135),
        .b(_T_326)
    );
    wire [41:0] notCDom_pos_firstNormAbsSigSum;
    MUX_UNSIGNED #(.width(42)) u_mux_1014 (
        .y(notCDom_pos_firstNormAbsSigSum),
        .sel(_T_311),
        .a(_T_319),
        .b(_T_327)
    );
    wire [31:0] _T_328;
    BITS #(.width(75), .high(49), .low(18)) bits_1015 (
        .y(_T_328),
        .in(complSigSum)
    );
    wire _T_329;
    BITS #(.width(2), .high(0), .low(0)) bits_1016 (
        .y(_T_329),
        .in(firstReduceComplSigSum)
    );
    wire [32:0] _T_330;
    CAT #(.width_a(32), .width_b(1)) cat_1017 (
        .y(_T_330),
        .a(_T_328),
        .b(_T_329)
    );
    wire [41:0] _T_331;
    BITS #(.width(75), .high(42), .low(1)) bits_1018 (
        .y(_T_331),
        .in(complSigSum)
    );
    wire _T_332;
    BITS #(.width(7), .high(5), .low(5)) bits_1019 (
        .y(_T_332),
        .in(estNormNeg_dist)
    );
    wire _T_333;
    BITS #(.width(7), .high(4), .low(4)) bits_1020 (
        .y(_T_333),
        .in(estNormNeg_dist)
    );
    wire [26:0] _T_334;
    BITS #(.width(75), .high(27), .low(1)) bits_1021 (
        .y(_T_334),
        .in(complSigSum)
    );
    wire [42:0] _T_335;
    SHL_UNSIGNED #(.width(27), .n(16)) u_shl_1022 (
        .y(_T_335),
        .in(_T_334)
    );
    wire [42:0] _T_336;
    wire [42:0] _WTEMP_136;
    PAD_UNSIGNED #(.width(42), .n(43)) u_pad_1023 (
        .y(_WTEMP_136),
        .in(_T_331)
    );
    MUX_UNSIGNED #(.width(43)) u_mux_1024 (
        .y(_T_336),
        .sel(_T_333),
        .a(_T_335),
        .b(_WTEMP_136)
    );
    wire _T_337;
    BITS #(.width(7), .high(4), .low(4)) bits_1025 (
        .y(_T_337),
        .in(estNormNeg_dist)
    );
    wire [10:0] _T_338;
    BITS #(.width(75), .high(11), .low(1)) bits_1026 (
        .y(_T_338),
        .in(complSigSum)
    );
    wire [42:0] _T_339;
    SHL_UNSIGNED #(.width(11), .n(32)) u_shl_1027 (
        .y(_T_339),
        .in(_T_338)
    );
    wire [42:0] _T_340;
    wire [42:0] _WTEMP_137;
    PAD_UNSIGNED #(.width(33), .n(43)) u_pad_1028 (
        .y(_WTEMP_137),
        .in(_T_330)
    );
    MUX_UNSIGNED #(.width(43)) u_mux_1029 (
        .y(_T_340),
        .sel(_T_337),
        .a(_WTEMP_137),
        .b(_T_339)
    );
    wire [42:0] notCDom_neg_cFirstNormAbsSigSum;
    MUX_UNSIGNED #(.width(43)) u_mux_1030 (
        .y(notCDom_neg_cFirstNormAbsSigSum),
        .sel(_T_332),
        .a(_T_336),
        .b(_T_340)
    );
    wire notCDom_signSigSum;
    BITS #(.width(75), .high(51), .low(51)) bits_1031 (
        .y(notCDom_signSigSum),
        .in(sigSum)
    );
    wire _T_342;
    EQ_UNSIGNED #(.width(1)) u_eq_1032 (
        .y(_T_342),
        .a(isZeroC),
        .b(1'h0)
    );
    wire _T_343;
    BITWISEAND #(.width(1)) bitwiseand_1033 (
        .y(_T_343),
        .a(doSubMags),
        .b(_T_342)
    );
    wire doNegSignSum;
    MUX_UNSIGNED #(.width(1)) u_mux_1034 (
        .y(doNegSignSum),
        .sel(io_fromPreMul_isCDominant),
        .a(_T_343),
        .b(notCDom_signSigSum)
    );
    wire [6:0] _T_344;
    assign _T_344 = estNormNeg_dist;
    wire [6:0] estNormDist;
    MUX_UNSIGNED #(.width(7)) u_mux_1035 (
        .y(estNormDist),
        .sel(io_fromPreMul_isCDominant),
        .a(CDom_estNormDist),
        .b(_T_344)
    );
    wire [42:0] _T_345;
    wire [42:0] _WTEMP_138;
    PAD_UNSIGNED #(.width(42), .n(43)) u_pad_1036 (
        .y(_WTEMP_138),
        .in(CDom_firstNormAbsSigSum)
    );
    MUX_UNSIGNED #(.width(43)) u_mux_1037 (
        .y(_T_345),
        .sel(io_fromPreMul_isCDominant),
        .a(_WTEMP_138),
        .b(notCDom_neg_cFirstNormAbsSigSum)
    );
    wire [41:0] _T_346;
    MUX_UNSIGNED #(.width(42)) u_mux_1038 (
        .y(_T_346),
        .sel(io_fromPreMul_isCDominant),
        .a(CDom_firstNormAbsSigSum),
        .b(notCDom_pos_firstNormAbsSigSum)
    );
    wire [42:0] cFirstNormAbsSigSum;
    wire [42:0] _WTEMP_139;
    PAD_UNSIGNED #(.width(42), .n(43)) u_pad_1039 (
        .y(_WTEMP_139),
        .in(_T_346)
    );
    MUX_UNSIGNED #(.width(43)) u_mux_1040 (
        .y(cFirstNormAbsSigSum),
        .sel(notCDom_signSigSum),
        .a(_T_345),
        .b(_WTEMP_139)
    );
    wire _T_348;
    EQ_UNSIGNED #(.width(1)) u_eq_1041 (
        .y(_T_348),
        .a(io_fromPreMul_isCDominant),
        .b(1'h0)
    );
    wire _T_350;
    EQ_UNSIGNED #(.width(1)) u_eq_1042 (
        .y(_T_350),
        .a(notCDom_signSigSum),
        .b(1'h0)
    );
    wire _T_351;
    BITWISEAND #(.width(1)) bitwiseand_1043 (
        .y(_T_351),
        .a(_T_348),
        .b(_T_350)
    );
    wire doIncrSig;
    BITWISEAND #(.width(1)) bitwiseand_1044 (
        .y(doIncrSig),
        .a(_T_351),
        .b(doSubMags)
    );
    wire [3:0] estNormDist_5;
    BITS #(.width(7), .high(3), .low(0)) bits_1045 (
        .y(estNormDist_5),
        .in(estNormDist)
    );
    wire [3:0] normTo2ShiftDist;
    BITWISENOT #(.width(4)) bitwisenot_1046 (
        .y(normTo2ShiftDist),
        .in(estNormDist_5)
    );
    wire [16:0] _T_353;
    DSHR_SIGNED #(.width_in(17), .width_n(4)) s_dshr_1047 (
        .y(_T_353),
        .in(-17'sh10000),
        .n(normTo2ShiftDist)
    );
    wire [14:0] _T_354;
    BITS #(.width(17), .high(15), .low(1)) bits_1048 (
        .y(_T_354),
        .in(_T_353)
    );
    wire [7:0] _T_355;
    BITS #(.width(15), .high(7), .low(0)) bits_1049 (
        .y(_T_355),
        .in(_T_354)
    );
    wire [7:0] _T_358;
    assign _T_358 = 8'hF0;
    wire [7:0] _T_359;
    assign _T_359 = 8'hF;
    wire [3:0] _T_360;
    SHR_UNSIGNED #(.width(8), .n(4)) u_shr_1050 (
        .y(_T_360),
        .in(_T_355)
    );
    wire [7:0] _T_361;
    wire [7:0] _WTEMP_140;
    PAD_UNSIGNED #(.width(4), .n(8)) u_pad_1051 (
        .y(_WTEMP_140),
        .in(_T_360)
    );
    BITWISEAND #(.width(8)) bitwiseand_1052 (
        .y(_T_361),
        .a(_WTEMP_140),
        .b(_T_359)
    );
    wire [3:0] _T_362;
    BITS #(.width(8), .high(3), .low(0)) bits_1053 (
        .y(_T_362),
        .in(_T_355)
    );
    wire [7:0] _T_363;
    SHL_UNSIGNED #(.width(4), .n(4)) u_shl_1054 (
        .y(_T_363),
        .in(_T_362)
    );
    wire [7:0] _T_364;
    assign _T_364 = 8'hF0;
    wire [7:0] _T_365;
    BITWISEAND #(.width(8)) bitwiseand_1055 (
        .y(_T_365),
        .a(_T_363),
        .b(_T_364)
    );
    wire [7:0] _T_366;
    BITWISEOR #(.width(8)) bitwiseor_1056 (
        .y(_T_366),
        .a(_T_361),
        .b(_T_365)
    );
    wire [5:0] _T_367;
    assign _T_367 = 6'hF;
    wire [7:0] _T_368;
    assign _T_368 = 8'h3C;
    wire [7:0] _T_369;
    assign _T_369 = 8'h33;
    wire [5:0] _T_370;
    SHR_UNSIGNED #(.width(8), .n(2)) u_shr_1057 (
        .y(_T_370),
        .in(_T_366)
    );
    wire [7:0] _T_371;
    wire [7:0] _WTEMP_141;
    PAD_UNSIGNED #(.width(6), .n(8)) u_pad_1058 (
        .y(_WTEMP_141),
        .in(_T_370)
    );
    BITWISEAND #(.width(8)) bitwiseand_1059 (
        .y(_T_371),
        .a(_WTEMP_141),
        .b(_T_369)
    );
    wire [5:0] _T_372;
    BITS #(.width(8), .high(5), .low(0)) bits_1060 (
        .y(_T_372),
        .in(_T_366)
    );
    wire [7:0] _T_373;
    SHL_UNSIGNED #(.width(6), .n(2)) u_shl_1061 (
        .y(_T_373),
        .in(_T_372)
    );
    wire [7:0] _T_374;
    assign _T_374 = 8'hCC;
    wire [7:0] _T_375;
    BITWISEAND #(.width(8)) bitwiseand_1062 (
        .y(_T_375),
        .a(_T_373),
        .b(_T_374)
    );
    wire [7:0] _T_376;
    BITWISEOR #(.width(8)) bitwiseor_1063 (
        .y(_T_376),
        .a(_T_371),
        .b(_T_375)
    );
    wire [6:0] _T_377;
    assign _T_377 = 7'h33;
    wire [7:0] _T_378;
    assign _T_378 = 8'h66;
    wire [7:0] _T_379;
    assign _T_379 = 8'h55;
    wire [6:0] _T_380;
    SHR_UNSIGNED #(.width(8), .n(1)) u_shr_1064 (
        .y(_T_380),
        .in(_T_376)
    );
    wire [7:0] _T_381;
    wire [7:0] _WTEMP_142;
    PAD_UNSIGNED #(.width(7), .n(8)) u_pad_1065 (
        .y(_WTEMP_142),
        .in(_T_380)
    );
    BITWISEAND #(.width(8)) bitwiseand_1066 (
        .y(_T_381),
        .a(_WTEMP_142),
        .b(_T_379)
    );
    wire [6:0] _T_382;
    BITS #(.width(8), .high(6), .low(0)) bits_1067 (
        .y(_T_382),
        .in(_T_376)
    );
    wire [7:0] _T_383;
    SHL_UNSIGNED #(.width(7), .n(1)) u_shl_1068 (
        .y(_T_383),
        .in(_T_382)
    );
    wire [7:0] _T_384;
    assign _T_384 = 8'hAA;
    wire [7:0] _T_385;
    BITWISEAND #(.width(8)) bitwiseand_1069 (
        .y(_T_385),
        .a(_T_383),
        .b(_T_384)
    );
    wire [7:0] _T_386;
    BITWISEOR #(.width(8)) bitwiseor_1070 (
        .y(_T_386),
        .a(_T_381),
        .b(_T_385)
    );
    wire [6:0] _T_387;
    BITS #(.width(15), .high(14), .low(8)) bits_1071 (
        .y(_T_387),
        .in(_T_354)
    );
    wire [3:0] _T_388;
    BITS #(.width(7), .high(3), .low(0)) bits_1072 (
        .y(_T_388),
        .in(_T_387)
    );
    wire [1:0] _T_389;
    BITS #(.width(4), .high(1), .low(0)) bits_1073 (
        .y(_T_389),
        .in(_T_388)
    );
    wire _T_390;
    BITS #(.width(2), .high(0), .low(0)) bits_1074 (
        .y(_T_390),
        .in(_T_389)
    );
    wire _T_391;
    BITS #(.width(2), .high(1), .low(1)) bits_1075 (
        .y(_T_391),
        .in(_T_389)
    );
    wire [1:0] _T_392;
    CAT #(.width_a(1), .width_b(1)) cat_1076 (
        .y(_T_392),
        .a(_T_390),
        .b(_T_391)
    );
    wire [1:0] _T_393;
    BITS #(.width(4), .high(3), .low(2)) bits_1077 (
        .y(_T_393),
        .in(_T_388)
    );
    wire _T_394;
    BITS #(.width(2), .high(0), .low(0)) bits_1078 (
        .y(_T_394),
        .in(_T_393)
    );
    wire _T_395;
    BITS #(.width(2), .high(1), .low(1)) bits_1079 (
        .y(_T_395),
        .in(_T_393)
    );
    wire [1:0] _T_396;
    CAT #(.width_a(1), .width_b(1)) cat_1080 (
        .y(_T_396),
        .a(_T_394),
        .b(_T_395)
    );
    wire [3:0] _T_397;
    CAT #(.width_a(2), .width_b(2)) cat_1081 (
        .y(_T_397),
        .a(_T_392),
        .b(_T_396)
    );
    wire [2:0] _T_398;
    BITS #(.width(7), .high(6), .low(4)) bits_1082 (
        .y(_T_398),
        .in(_T_387)
    );
    wire [1:0] _T_399;
    BITS #(.width(3), .high(1), .low(0)) bits_1083 (
        .y(_T_399),
        .in(_T_398)
    );
    wire _T_400;
    BITS #(.width(2), .high(0), .low(0)) bits_1084 (
        .y(_T_400),
        .in(_T_399)
    );
    wire _T_401;
    BITS #(.width(2), .high(1), .low(1)) bits_1085 (
        .y(_T_401),
        .in(_T_399)
    );
    wire [1:0] _T_402;
    CAT #(.width_a(1), .width_b(1)) cat_1086 (
        .y(_T_402),
        .a(_T_400),
        .b(_T_401)
    );
    wire _T_403;
    BITS #(.width(3), .high(2), .low(2)) bits_1087 (
        .y(_T_403),
        .in(_T_398)
    );
    wire [2:0] _T_404;
    CAT #(.width_a(2), .width_b(1)) cat_1088 (
        .y(_T_404),
        .a(_T_402),
        .b(_T_403)
    );
    wire [6:0] _T_405;
    CAT #(.width_a(4), .width_b(3)) cat_1089 (
        .y(_T_405),
        .a(_T_397),
        .b(_T_404)
    );
    wire [14:0] _T_406;
    CAT #(.width_a(8), .width_b(7)) cat_1090 (
        .y(_T_406),
        .a(_T_386),
        .b(_T_405)
    );
    wire [15:0] absSigSumExtraMask;
    CAT #(.width_a(15), .width_b(1)) cat_1091 (
        .y(absSigSumExtraMask),
        .a(_T_406),
        .b(1'h1)
    );
    wire [41:0] _T_408;
    BITS #(.width(43), .high(42), .low(1)) bits_1092 (
        .y(_T_408),
        .in(cFirstNormAbsSigSum)
    );
    wire [41:0] _T_409;
    DSHR_UNSIGNED #(.width_in(42), .width_n(4)) u_dshr_1093 (
        .y(_T_409),
        .in(_T_408),
        .n(normTo2ShiftDist)
    );
    wire [15:0] _T_410;
    BITS #(.width(43), .high(15), .low(0)) bits_1094 (
        .y(_T_410),
        .in(cFirstNormAbsSigSum)
    );
    wire [15:0] _T_411;
    BITWISENOT #(.width(16)) bitwisenot_1095 (
        .y(_T_411),
        .in(_T_410)
    );
    wire [15:0] _T_412;
    BITWISEAND #(.width(16)) bitwiseand_1096 (
        .y(_T_412),
        .a(_T_411),
        .b(absSigSumExtraMask)
    );
    wire _T_414;
    wire [15:0] _WTEMP_143;
    PAD_UNSIGNED #(.width(1), .n(16)) u_pad_1097 (
        .y(_WTEMP_143),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(16)) u_eq_1098 (
        .y(_T_414),
        .a(_T_412),
        .b(_WTEMP_143)
    );
    wire [15:0] _T_415;
    BITS #(.width(43), .high(15), .low(0)) bits_1099 (
        .y(_T_415),
        .in(cFirstNormAbsSigSum)
    );
    wire [15:0] _T_416;
    BITWISEAND #(.width(16)) bitwiseand_1100 (
        .y(_T_416),
        .a(_T_415),
        .b(absSigSumExtraMask)
    );
    wire _T_418;
    wire [15:0] _WTEMP_144;
    PAD_UNSIGNED #(.width(1), .n(16)) u_pad_1101 (
        .y(_WTEMP_144),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(16)) u_neq_1102 (
        .y(_T_418),
        .a(_T_416),
        .b(_WTEMP_144)
    );
    wire _T_419;
    MUX_UNSIGNED #(.width(1)) u_mux_1103 (
        .y(_T_419),
        .sel(doIncrSig),
        .a(_T_414),
        .b(_T_418)
    );
    wire [42:0] _T_420;
    CAT #(.width_a(42), .width_b(1)) cat_1104 (
        .y(_T_420),
        .a(_T_409),
        .b(_T_419)
    );
    wire [27:0] sigX3;
    BITS #(.width(43), .high(27), .low(0)) bits_1105 (
        .y(sigX3),
        .in(_T_420)
    );
    wire [1:0] _T_421;
    BITS #(.width(28), .high(27), .low(26)) bits_1106 (
        .y(_T_421),
        .in(sigX3)
    );
    wire sigX3Shift1;
    wire [1:0] _WTEMP_145;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_1107 (
        .y(_WTEMP_145),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(2)) u_eq_1108 (
        .y(sigX3Shift1),
        .a(_T_421),
        .b(_WTEMP_145)
    );
    wire [11:0] _T_423;
    wire [10:0] _WTEMP_146;
    PAD_UNSIGNED #(.width(7), .n(11)) u_pad_1109 (
        .y(_WTEMP_146),
        .in(estNormDist)
    );
    SUB_UNSIGNED #(.width(11)) u_sub_1110 (
        .y(_T_423),
        .a(io_fromPreMul_sExpSum),
        .b(_WTEMP_146)
    );
    wire [11:0] _T_424;
    ASUINT #(.width(12)) asuint_1111 (
        .y(_T_424),
        .in(_T_423)
    );
    wire [10:0] sExpX3;
    TAIL #(.width(12), .n(1)) tail_1112 (
        .y(sExpX3),
        .in(_T_424)
    );
    wire [2:0] _T_425;
    BITS #(.width(28), .high(27), .low(25)) bits_1113 (
        .y(_T_425),
        .in(sigX3)
    );
    wire isZeroY;
    wire [2:0] _WTEMP_147;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_1114 (
        .y(_WTEMP_147),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(3)) u_eq_1115 (
        .y(isZeroY),
        .a(_T_425),
        .b(_WTEMP_147)
    );
    wire _T_427;
    BITWISEXOR #(.width(1)) bitwisexor_1116 (
        .y(_T_427),
        .a(io_fromPreMul_signProd),
        .b(doNegSignSum)
    );
    wire signY;
    MUX_UNSIGNED #(.width(1)) u_mux_1117 (
        .y(signY),
        .sel(isZeroY),
        .a(signZeroNotEqOpSigns),
        .b(_T_427)
    );
    wire [9:0] sExpX3_13;
    BITS #(.width(11), .high(9), .low(0)) bits_1118 (
        .y(sExpX3_13),
        .in(sExpX3)
    );
    wire _T_428;
    BITS #(.width(11), .high(10), .low(10)) bits_1119 (
        .y(_T_428),
        .in(sExpX3)
    );
    wire _T_429;
    BITS #(.width(1), .high(0), .low(0)) bits_1120 (
        .y(_T_429),
        .in(_T_428)
    );
    wire [26:0] _T_432;
    MUX_UNSIGNED #(.width(27)) u_mux_1121 (
        .y(_T_432),
        .sel(_T_429),
        .a(27'h7FFFFFF),
        .b(27'h0)
    );
    wire [9:0] _T_433;
    BITWISENOT #(.width(10)) bitwisenot_1122 (
        .y(_T_433),
        .in(sExpX3_13)
    );
    wire _T_434;
    BITS #(.width(10), .high(9), .low(9)) bits_1123 (
        .y(_T_434),
        .in(_T_433)
    );
    wire [8:0] _T_435;
    BITS #(.width(10), .high(8), .low(0)) bits_1124 (
        .y(_T_435),
        .in(_T_433)
    );
    wire _T_436;
    BITS #(.width(9), .high(8), .low(8)) bits_1125 (
        .y(_T_436),
        .in(_T_435)
    );
    wire [7:0] _T_437;
    BITS #(.width(9), .high(7), .low(0)) bits_1126 (
        .y(_T_437),
        .in(_T_435)
    );
    wire _T_438;
    BITS #(.width(8), .high(7), .low(7)) bits_1127 (
        .y(_T_438),
        .in(_T_437)
    );
    wire [6:0] _T_439;
    BITS #(.width(8), .high(6), .low(0)) bits_1128 (
        .y(_T_439),
        .in(_T_437)
    );
    wire _T_440;
    BITS #(.width(7), .high(6), .low(6)) bits_1129 (
        .y(_T_440),
        .in(_T_439)
    );
    wire [5:0] _T_441;
    BITS #(.width(7), .high(5), .low(0)) bits_1130 (
        .y(_T_441),
        .in(_T_439)
    );
    wire [64:0] _T_444;
    DSHR_SIGNED #(.width_in(65), .width_n(6)) s_dshr_1131 (
        .y(_T_444),
        .in(-65'sh10000000000000000),
        .n(_T_441)
    );
    wire [20:0] _T_445;
    BITS #(.width(65), .high(63), .low(43)) bits_1132 (
        .y(_T_445),
        .in(_T_444)
    );
    wire [15:0] _T_446;
    BITS #(.width(21), .high(15), .low(0)) bits_1133 (
        .y(_T_446),
        .in(_T_445)
    );
    wire [15:0] _T_449;
    assign _T_449 = 16'hFF00;
    wire [15:0] _T_450;
    assign _T_450 = 16'hFF;
    wire [7:0] _T_451;
    SHR_UNSIGNED #(.width(16), .n(8)) u_shr_1134 (
        .y(_T_451),
        .in(_T_446)
    );
    wire [15:0] _T_452;
    wire [15:0] _WTEMP_148;
    PAD_UNSIGNED #(.width(8), .n(16)) u_pad_1135 (
        .y(_WTEMP_148),
        .in(_T_451)
    );
    BITWISEAND #(.width(16)) bitwiseand_1136 (
        .y(_T_452),
        .a(_WTEMP_148),
        .b(_T_450)
    );
    wire [7:0] _T_453;
    BITS #(.width(16), .high(7), .low(0)) bits_1137 (
        .y(_T_453),
        .in(_T_446)
    );
    wire [15:0] _T_454;
    SHL_UNSIGNED #(.width(8), .n(8)) u_shl_1138 (
        .y(_T_454),
        .in(_T_453)
    );
    wire [15:0] _T_455;
    assign _T_455 = 16'hFF00;
    wire [15:0] _T_456;
    BITWISEAND #(.width(16)) bitwiseand_1139 (
        .y(_T_456),
        .a(_T_454),
        .b(_T_455)
    );
    wire [15:0] _T_457;
    BITWISEOR #(.width(16)) bitwiseor_1140 (
        .y(_T_457),
        .a(_T_452),
        .b(_T_456)
    );
    wire [11:0] _T_458;
    assign _T_458 = 12'hFF;
    wire [15:0] _T_459;
    assign _T_459 = 16'hFF0;
    wire [15:0] _T_460;
    assign _T_460 = 16'hF0F;
    wire [11:0] _T_461;
    SHR_UNSIGNED #(.width(16), .n(4)) u_shr_1141 (
        .y(_T_461),
        .in(_T_457)
    );
    wire [15:0] _T_462;
    wire [15:0] _WTEMP_149;
    PAD_UNSIGNED #(.width(12), .n(16)) u_pad_1142 (
        .y(_WTEMP_149),
        .in(_T_461)
    );
    BITWISEAND #(.width(16)) bitwiseand_1143 (
        .y(_T_462),
        .a(_WTEMP_149),
        .b(_T_460)
    );
    wire [11:0] _T_463;
    BITS #(.width(16), .high(11), .low(0)) bits_1144 (
        .y(_T_463),
        .in(_T_457)
    );
    wire [15:0] _T_464;
    SHL_UNSIGNED #(.width(12), .n(4)) u_shl_1145 (
        .y(_T_464),
        .in(_T_463)
    );
    wire [15:0] _T_465;
    assign _T_465 = 16'hF0F0;
    wire [15:0] _T_466;
    BITWISEAND #(.width(16)) bitwiseand_1146 (
        .y(_T_466),
        .a(_T_464),
        .b(_T_465)
    );
    wire [15:0] _T_467;
    BITWISEOR #(.width(16)) bitwiseor_1147 (
        .y(_T_467),
        .a(_T_462),
        .b(_T_466)
    );
    wire [13:0] _T_468;
    assign _T_468 = 14'hF0F;
    wire [15:0] _T_469;
    assign _T_469 = 16'h3C3C;
    wire [15:0] _T_470;
    assign _T_470 = 16'h3333;
    wire [13:0] _T_471;
    SHR_UNSIGNED #(.width(16), .n(2)) u_shr_1148 (
        .y(_T_471),
        .in(_T_467)
    );
    wire [15:0] _T_472;
    wire [15:0] _WTEMP_150;
    PAD_UNSIGNED #(.width(14), .n(16)) u_pad_1149 (
        .y(_WTEMP_150),
        .in(_T_471)
    );
    BITWISEAND #(.width(16)) bitwiseand_1150 (
        .y(_T_472),
        .a(_WTEMP_150),
        .b(_T_470)
    );
    wire [13:0] _T_473;
    BITS #(.width(16), .high(13), .low(0)) bits_1151 (
        .y(_T_473),
        .in(_T_467)
    );
    wire [15:0] _T_474;
    SHL_UNSIGNED #(.width(14), .n(2)) u_shl_1152 (
        .y(_T_474),
        .in(_T_473)
    );
    wire [15:0] _T_475;
    assign _T_475 = 16'hCCCC;
    wire [15:0] _T_476;
    BITWISEAND #(.width(16)) bitwiseand_1153 (
        .y(_T_476),
        .a(_T_474),
        .b(_T_475)
    );
    wire [15:0] _T_477;
    BITWISEOR #(.width(16)) bitwiseor_1154 (
        .y(_T_477),
        .a(_T_472),
        .b(_T_476)
    );
    wire [14:0] _T_478;
    assign _T_478 = 15'h3333;
    wire [15:0] _T_479;
    assign _T_479 = 16'h6666;
    wire [15:0] _T_480;
    assign _T_480 = 16'h5555;
    wire [14:0] _T_481;
    SHR_UNSIGNED #(.width(16), .n(1)) u_shr_1155 (
        .y(_T_481),
        .in(_T_477)
    );
    wire [15:0] _T_482;
    wire [15:0] _WTEMP_151;
    PAD_UNSIGNED #(.width(15), .n(16)) u_pad_1156 (
        .y(_WTEMP_151),
        .in(_T_481)
    );
    BITWISEAND #(.width(16)) bitwiseand_1157 (
        .y(_T_482),
        .a(_WTEMP_151),
        .b(_T_480)
    );
    wire [14:0] _T_483;
    BITS #(.width(16), .high(14), .low(0)) bits_1158 (
        .y(_T_483),
        .in(_T_477)
    );
    wire [15:0] _T_484;
    SHL_UNSIGNED #(.width(15), .n(1)) u_shl_1159 (
        .y(_T_484),
        .in(_T_483)
    );
    wire [15:0] _T_485;
    assign _T_485 = 16'hAAAA;
    wire [15:0] _T_486;
    BITWISEAND #(.width(16)) bitwiseand_1160 (
        .y(_T_486),
        .a(_T_484),
        .b(_T_485)
    );
    wire [15:0] _T_487;
    BITWISEOR #(.width(16)) bitwiseor_1161 (
        .y(_T_487),
        .a(_T_482),
        .b(_T_486)
    );
    wire [4:0] _T_488;
    BITS #(.width(21), .high(20), .low(16)) bits_1162 (
        .y(_T_488),
        .in(_T_445)
    );
    wire [3:0] _T_489;
    BITS #(.width(5), .high(3), .low(0)) bits_1163 (
        .y(_T_489),
        .in(_T_488)
    );
    wire [1:0] _T_490;
    BITS #(.width(4), .high(1), .low(0)) bits_1164 (
        .y(_T_490),
        .in(_T_489)
    );
    wire _T_491;
    BITS #(.width(2), .high(0), .low(0)) bits_1165 (
        .y(_T_491),
        .in(_T_490)
    );
    wire _T_492;
    BITS #(.width(2), .high(1), .low(1)) bits_1166 (
        .y(_T_492),
        .in(_T_490)
    );
    wire [1:0] _T_493;
    CAT #(.width_a(1), .width_b(1)) cat_1167 (
        .y(_T_493),
        .a(_T_491),
        .b(_T_492)
    );
    wire [1:0] _T_494;
    BITS #(.width(4), .high(3), .low(2)) bits_1168 (
        .y(_T_494),
        .in(_T_489)
    );
    wire _T_495;
    BITS #(.width(2), .high(0), .low(0)) bits_1169 (
        .y(_T_495),
        .in(_T_494)
    );
    wire _T_496;
    BITS #(.width(2), .high(1), .low(1)) bits_1170 (
        .y(_T_496),
        .in(_T_494)
    );
    wire [1:0] _T_497;
    CAT #(.width_a(1), .width_b(1)) cat_1171 (
        .y(_T_497),
        .a(_T_495),
        .b(_T_496)
    );
    wire [3:0] _T_498;
    CAT #(.width_a(2), .width_b(2)) cat_1172 (
        .y(_T_498),
        .a(_T_493),
        .b(_T_497)
    );
    wire _T_499;
    BITS #(.width(5), .high(4), .low(4)) bits_1173 (
        .y(_T_499),
        .in(_T_488)
    );
    wire [4:0] _T_500;
    CAT #(.width_a(4), .width_b(1)) cat_1174 (
        .y(_T_500),
        .a(_T_498),
        .b(_T_499)
    );
    wire [20:0] _T_501;
    CAT #(.width_a(16), .width_b(5)) cat_1175 (
        .y(_T_501),
        .a(_T_487),
        .b(_T_500)
    );
    wire [20:0] _T_502;
    BITWISENOT #(.width(21)) bitwisenot_1176 (
        .y(_T_502),
        .in(_T_501)
    );
    wire [20:0] _T_503;
    wire [20:0] _WTEMP_152;
    PAD_UNSIGNED #(.width(1), .n(21)) u_pad_1177 (
        .y(_WTEMP_152),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(21)) u_mux_1178 (
        .y(_T_503),
        .sel(_T_440),
        .a(_WTEMP_152),
        .b(_T_502)
    );
    wire [20:0] _T_504;
    BITWISENOT #(.width(21)) bitwisenot_1179 (
        .y(_T_504),
        .in(_T_503)
    );
    wire [24:0] _T_506;
    CAT #(.width_a(21), .width_b(4)) cat_1180 (
        .y(_T_506),
        .a(_T_504),
        .b(4'hF)
    );
    wire _T_507;
    BITS #(.width(7), .high(6), .low(6)) bits_1181 (
        .y(_T_507),
        .in(_T_439)
    );
    wire [5:0] _T_508;
    BITS #(.width(7), .high(5), .low(0)) bits_1182 (
        .y(_T_508),
        .in(_T_439)
    );
    wire [64:0] _T_510;
    DSHR_SIGNED #(.width_in(65), .width_n(6)) s_dshr_1183 (
        .y(_T_510),
        .in(-65'sh10000000000000000),
        .n(_T_508)
    );
    wire [3:0] _T_511;
    BITS #(.width(65), .high(3), .low(0)) bits_1184 (
        .y(_T_511),
        .in(_T_510)
    );
    wire [1:0] _T_512;
    BITS #(.width(4), .high(1), .low(0)) bits_1185 (
        .y(_T_512),
        .in(_T_511)
    );
    wire _T_513;
    BITS #(.width(2), .high(0), .low(0)) bits_1186 (
        .y(_T_513),
        .in(_T_512)
    );
    wire _T_514;
    BITS #(.width(2), .high(1), .low(1)) bits_1187 (
        .y(_T_514),
        .in(_T_512)
    );
    wire [1:0] _T_515;
    CAT #(.width_a(1), .width_b(1)) cat_1188 (
        .y(_T_515),
        .a(_T_513),
        .b(_T_514)
    );
    wire [1:0] _T_516;
    BITS #(.width(4), .high(3), .low(2)) bits_1189 (
        .y(_T_516),
        .in(_T_511)
    );
    wire _T_517;
    BITS #(.width(2), .high(0), .low(0)) bits_1190 (
        .y(_T_517),
        .in(_T_516)
    );
    wire _T_518;
    BITS #(.width(2), .high(1), .low(1)) bits_1191 (
        .y(_T_518),
        .in(_T_516)
    );
    wire [1:0] _T_519;
    CAT #(.width_a(1), .width_b(1)) cat_1192 (
        .y(_T_519),
        .a(_T_517),
        .b(_T_518)
    );
    wire [3:0] _T_520;
    CAT #(.width_a(2), .width_b(2)) cat_1193 (
        .y(_T_520),
        .a(_T_515),
        .b(_T_519)
    );
    wire [3:0] _T_522;
    wire [3:0] _WTEMP_153;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1194 (
        .y(_WTEMP_153),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(4)) u_mux_1195 (
        .y(_T_522),
        .sel(_T_507),
        .a(_T_520),
        .b(_WTEMP_153)
    );
    wire [24:0] _T_523;
    wire [24:0] _WTEMP_154;
    PAD_UNSIGNED #(.width(4), .n(25)) u_pad_1196 (
        .y(_WTEMP_154),
        .in(_T_522)
    );
    MUX_UNSIGNED #(.width(25)) u_mux_1197 (
        .y(_T_523),
        .sel(_T_438),
        .a(_T_506),
        .b(_WTEMP_154)
    );
    wire [24:0] _T_525;
    wire [24:0] _WTEMP_155;
    PAD_UNSIGNED #(.width(1), .n(25)) u_pad_1198 (
        .y(_WTEMP_155),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(25)) u_mux_1199 (
        .y(_T_525),
        .sel(_T_436),
        .a(_T_523),
        .b(_WTEMP_155)
    );
    wire [24:0] _T_527;
    wire [24:0] _WTEMP_156;
    PAD_UNSIGNED #(.width(1), .n(25)) u_pad_1200 (
        .y(_WTEMP_156),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(25)) u_mux_1201 (
        .y(_T_527),
        .sel(_T_434),
        .a(_T_525),
        .b(_WTEMP_156)
    );
    wire _T_528;
    BITS #(.width(28), .high(26), .low(26)) bits_1202 (
        .y(_T_528),
        .in(sigX3)
    );
    wire [24:0] _T_529;
    wire [24:0] _WTEMP_157;
    PAD_UNSIGNED #(.width(1), .n(25)) u_pad_1203 (
        .y(_WTEMP_157),
        .in(_T_528)
    );
    BITWISEOR #(.width(25)) bitwiseor_1204 (
        .y(_T_529),
        .a(_T_527),
        .b(_WTEMP_157)
    );
    wire [26:0] _T_531;
    CAT #(.width_a(25), .width_b(2)) cat_1205 (
        .y(_T_531),
        .a(_T_529),
        .b(2'h3)
    );
    wire [26:0] roundMask;
    BITWISEOR #(.width(27)) bitwiseor_1206 (
        .y(roundMask),
        .a(_T_432),
        .b(_T_531)
    );
    wire [25:0] _T_532;
    SHR_UNSIGNED #(.width(27), .n(1)) u_shr_1207 (
        .y(_T_532),
        .in(roundMask)
    );
    wire [25:0] _T_533;
    BITWISENOT #(.width(26)) bitwisenot_1208 (
        .y(_T_533),
        .in(_T_532)
    );
    wire [26:0] roundPosMask;
    wire [26:0] _WTEMP_158;
    PAD_UNSIGNED #(.width(26), .n(27)) u_pad_1209 (
        .y(_WTEMP_158),
        .in(_T_533)
    );
    BITWISEAND #(.width(27)) bitwiseand_1210 (
        .y(roundPosMask),
        .a(_WTEMP_158),
        .b(roundMask)
    );
    wire [27:0] _T_534;
    wire [27:0] _WTEMP_159;
    PAD_UNSIGNED #(.width(27), .n(28)) u_pad_1211 (
        .y(_WTEMP_159),
        .in(roundPosMask)
    );
    BITWISEAND #(.width(28)) bitwiseand_1212 (
        .y(_T_534),
        .a(sigX3),
        .b(_WTEMP_159)
    );
    wire roundPosBit;
    wire [27:0] _WTEMP_160;
    PAD_UNSIGNED #(.width(1), .n(28)) u_pad_1213 (
        .y(_WTEMP_160),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(28)) u_neq_1214 (
        .y(roundPosBit),
        .a(_T_534),
        .b(_WTEMP_160)
    );
    wire [25:0] _T_536;
    SHR_UNSIGNED #(.width(27), .n(1)) u_shr_1215 (
        .y(_T_536),
        .in(roundMask)
    );
    wire [27:0] _T_537;
    wire [27:0] _WTEMP_161;
    PAD_UNSIGNED #(.width(26), .n(28)) u_pad_1216 (
        .y(_WTEMP_161),
        .in(_T_536)
    );
    BITWISEAND #(.width(28)) bitwiseand_1217 (
        .y(_T_537),
        .a(sigX3),
        .b(_WTEMP_161)
    );
    wire anyRoundExtra;
    wire [27:0] _WTEMP_162;
    PAD_UNSIGNED #(.width(1), .n(28)) u_pad_1218 (
        .y(_WTEMP_162),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(28)) u_neq_1219 (
        .y(anyRoundExtra),
        .a(_T_537),
        .b(_WTEMP_162)
    );
    wire [27:0] _T_539;
    BITWISENOT #(.width(28)) bitwisenot_1220 (
        .y(_T_539),
        .in(sigX3)
    );
    wire [25:0] _T_540;
    SHR_UNSIGNED #(.width(27), .n(1)) u_shr_1221 (
        .y(_T_540),
        .in(roundMask)
    );
    wire [27:0] _T_541;
    wire [27:0] _WTEMP_163;
    PAD_UNSIGNED #(.width(26), .n(28)) u_pad_1222 (
        .y(_WTEMP_163),
        .in(_T_540)
    );
    BITWISEAND #(.width(28)) bitwiseand_1223 (
        .y(_T_541),
        .a(_T_539),
        .b(_WTEMP_163)
    );
    wire allRoundExtra;
    wire [27:0] _WTEMP_164;
    PAD_UNSIGNED #(.width(1), .n(28)) u_pad_1224 (
        .y(_WTEMP_164),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(28)) u_eq_1225 (
        .y(allRoundExtra),
        .a(_T_541),
        .b(_WTEMP_164)
    );
    wire anyRound;
    BITWISEOR #(.width(1)) bitwiseor_1226 (
        .y(anyRound),
        .a(roundPosBit),
        .b(anyRoundExtra)
    );
    wire allRound;
    BITWISEAND #(.width(1)) bitwiseand_1227 (
        .y(allRound),
        .a(roundPosBit),
        .b(allRoundExtra)
    );
    wire roundDirectUp;
    MUX_UNSIGNED #(.width(1)) u_mux_1228 (
        .y(roundDirectUp),
        .sel(signY),
        .a(roundingMode_min),
        .b(roundingMode_max)
    );
    wire _T_544;
    EQ_UNSIGNED #(.width(1)) u_eq_1229 (
        .y(_T_544),
        .a(doIncrSig),
        .b(1'h0)
    );
    wire _T_545;
    BITWISEAND #(.width(1)) bitwiseand_1230 (
        .y(_T_545),
        .a(_T_544),
        .b(roundingMode_nearest_even)
    );
    wire _T_546;
    BITWISEAND #(.width(1)) bitwiseand_1231 (
        .y(_T_546),
        .a(_T_545),
        .b(roundPosBit)
    );
    wire _T_547;
    BITWISEAND #(.width(1)) bitwiseand_1232 (
        .y(_T_547),
        .a(_T_546),
        .b(anyRoundExtra)
    );
    wire _T_549;
    EQ_UNSIGNED #(.width(1)) u_eq_1233 (
        .y(_T_549),
        .a(doIncrSig),
        .b(1'h0)
    );
    wire _T_550;
    BITWISEAND #(.width(1)) bitwiseand_1234 (
        .y(_T_550),
        .a(_T_549),
        .b(roundDirectUp)
    );
    wire _T_551;
    BITWISEAND #(.width(1)) bitwiseand_1235 (
        .y(_T_551),
        .a(_T_550),
        .b(anyRound)
    );
    wire _T_552;
    BITWISEOR #(.width(1)) bitwiseor_1236 (
        .y(_T_552),
        .a(_T_547),
        .b(_T_551)
    );
    wire _T_553;
    BITWISEAND #(.width(1)) bitwiseand_1237 (
        .y(_T_553),
        .a(doIncrSig),
        .b(allRound)
    );
    wire _T_554;
    BITWISEOR #(.width(1)) bitwiseor_1238 (
        .y(_T_554),
        .a(_T_552),
        .b(_T_553)
    );
    wire _T_555;
    BITWISEAND #(.width(1)) bitwiseand_1239 (
        .y(_T_555),
        .a(doIncrSig),
        .b(roundingMode_nearest_even)
    );
    wire _T_556;
    BITWISEAND #(.width(1)) bitwiseand_1240 (
        .y(_T_556),
        .a(_T_555),
        .b(roundPosBit)
    );
    wire _T_557;
    BITWISEOR #(.width(1)) bitwiseor_1241 (
        .y(_T_557),
        .a(_T_554),
        .b(_T_556)
    );
    wire _T_558;
    BITWISEAND #(.width(1)) bitwiseand_1242 (
        .y(_T_558),
        .a(doIncrSig),
        .b(roundDirectUp)
    );
    wire _T_560;
    BITWISEAND #(.width(1)) bitwiseand_1243 (
        .y(_T_560),
        .a(_T_558),
        .b(1'h1)
    );
    wire roundUp;
    BITWISEOR #(.width(1)) bitwiseor_1244 (
        .y(roundUp),
        .a(_T_557),
        .b(_T_560)
    );
    wire _T_562;
    EQ_UNSIGNED #(.width(1)) u_eq_1245 (
        .y(_T_562),
        .a(roundPosBit),
        .b(1'h0)
    );
    wire _T_563;
    BITWISEAND #(.width(1)) bitwiseand_1246 (
        .y(_T_563),
        .a(roundingMode_nearest_even),
        .b(_T_562)
    );
    wire _T_564;
    BITWISEAND #(.width(1)) bitwiseand_1247 (
        .y(_T_564),
        .a(_T_563),
        .b(allRoundExtra)
    );
    wire _T_565;
    BITWISEAND #(.width(1)) bitwiseand_1248 (
        .y(_T_565),
        .a(roundingMode_nearest_even),
        .b(roundPosBit)
    );
    wire _T_567;
    EQ_UNSIGNED #(.width(1)) u_eq_1249 (
        .y(_T_567),
        .a(anyRoundExtra),
        .b(1'h0)
    );
    wire _T_568;
    BITWISEAND #(.width(1)) bitwiseand_1250 (
        .y(_T_568),
        .a(_T_565),
        .b(_T_567)
    );
    wire roundEven;
    MUX_UNSIGNED #(.width(1)) u_mux_1251 (
        .y(roundEven),
        .sel(doIncrSig),
        .a(_T_564),
        .b(_T_568)
    );
    wire _T_570;
    EQ_UNSIGNED #(.width(1)) u_eq_1252 (
        .y(_T_570),
        .a(allRound),
        .b(1'h0)
    );
    wire inexactY;
    MUX_UNSIGNED #(.width(1)) u_mux_1253 (
        .y(inexactY),
        .sel(doIncrSig),
        .a(_T_570),
        .b(anyRound)
    );
    wire [27:0] _T_571;
    wire [27:0] _WTEMP_165;
    PAD_UNSIGNED #(.width(27), .n(28)) u_pad_1254 (
        .y(_WTEMP_165),
        .in(roundMask)
    );
    BITWISEOR #(.width(28)) bitwiseor_1255 (
        .y(_T_571),
        .a(sigX3),
        .b(_WTEMP_165)
    );
    wire [25:0] _T_572;
    SHR_UNSIGNED #(.width(28), .n(2)) u_shr_1256 (
        .y(_T_572),
        .in(_T_571)
    );
    wire [26:0] _T_574;
    wire [25:0] _WTEMP_166;
    PAD_UNSIGNED #(.width(1), .n(26)) u_pad_1257 (
        .y(_WTEMP_166),
        .in(1'h1)
    );
    ADD_UNSIGNED #(.width(26)) u_add_1258 (
        .y(_T_574),
        .a(_T_572),
        .b(_WTEMP_166)
    );
    wire [25:0] _T_575;
    TAIL #(.width(27), .n(1)) tail_1259 (
        .y(_T_575),
        .in(_T_574)
    );
    wire [25:0] roundUp_sigY3;
    BITS #(.width(26), .high(25), .low(0)) bits_1260 (
        .y(roundUp_sigY3),
        .in(_T_575)
    );
    wire _T_577;
    EQ_UNSIGNED #(.width(1)) u_eq_1261 (
        .y(_T_577),
        .a(roundUp),
        .b(1'h0)
    );
    wire _T_579;
    EQ_UNSIGNED #(.width(1)) u_eq_1262 (
        .y(_T_579),
        .a(roundEven),
        .b(1'h0)
    );
    wire _T_580;
    BITWISEAND #(.width(1)) bitwiseand_1263 (
        .y(_T_580),
        .a(_T_577),
        .b(_T_579)
    );
    wire [26:0] _T_581;
    BITWISENOT #(.width(27)) bitwisenot_1264 (
        .y(_T_581),
        .in(roundMask)
    );
    wire [27:0] _T_582;
    wire [27:0] _WTEMP_167;
    PAD_UNSIGNED #(.width(27), .n(28)) u_pad_1265 (
        .y(_WTEMP_167),
        .in(_T_581)
    );
    BITWISEAND #(.width(28)) bitwiseand_1266 (
        .y(_T_582),
        .a(sigX3),
        .b(_WTEMP_167)
    );
    wire [25:0] _T_583;
    SHR_UNSIGNED #(.width(28), .n(2)) u_shr_1267 (
        .y(_T_583),
        .in(_T_582)
    );
    wire [25:0] _T_585;
    wire [25:0] _WTEMP_168;
    PAD_UNSIGNED #(.width(1), .n(26)) u_pad_1268 (
        .y(_WTEMP_168),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(26)) u_mux_1269 (
        .y(_T_585),
        .sel(_T_580),
        .a(_T_583),
        .b(_WTEMP_168)
    );
    wire [25:0] _T_587;
    wire [25:0] _WTEMP_169;
    PAD_UNSIGNED #(.width(1), .n(26)) u_pad_1270 (
        .y(_WTEMP_169),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(26)) u_mux_1271 (
        .y(_T_587),
        .sel(roundUp),
        .a(roundUp_sigY3),
        .b(_WTEMP_169)
    );
    wire [25:0] _T_588;
    BITWISEOR #(.width(26)) bitwiseor_1272 (
        .y(_T_588),
        .a(_T_585),
        .b(_T_587)
    );
    wire [25:0] _T_589;
    SHR_UNSIGNED #(.width(27), .n(1)) u_shr_1273 (
        .y(_T_589),
        .in(roundMask)
    );
    wire [25:0] _T_590;
    BITWISENOT #(.width(26)) bitwisenot_1274 (
        .y(_T_590),
        .in(_T_589)
    );
    wire [25:0] _T_591;
    BITWISEAND #(.width(26)) bitwiseand_1275 (
        .y(_T_591),
        .a(roundUp_sigY3),
        .b(_T_590)
    );
    wire [25:0] _T_593;
    wire [25:0] _WTEMP_170;
    PAD_UNSIGNED #(.width(1), .n(26)) u_pad_1276 (
        .y(_WTEMP_170),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(26)) u_mux_1277 (
        .y(_T_593),
        .sel(roundEven),
        .a(_T_591),
        .b(_WTEMP_170)
    );
    wire [25:0] sigY3;
    BITWISEOR #(.width(26)) bitwiseor_1278 (
        .y(sigY3),
        .a(_T_588),
        .b(_T_593)
    );
    wire _T_594;
    BITS #(.width(26), .high(25), .low(25)) bits_1279 (
        .y(_T_594),
        .in(sigY3)
    );
    wire [11:0] _T_596;
    wire [10:0] _WTEMP_171;
    PAD_UNSIGNED #(.width(1), .n(11)) u_pad_1280 (
        .y(_WTEMP_171),
        .in(1'h1)
    );
    ADD_UNSIGNED #(.width(11)) u_add_1281 (
        .y(_T_596),
        .a(sExpX3),
        .b(_WTEMP_171)
    );
    wire [10:0] _T_597;
    TAIL #(.width(12), .n(1)) tail_1282 (
        .y(_T_597),
        .in(_T_596)
    );
    wire [10:0] _T_599;
    wire [10:0] _WTEMP_172;
    PAD_UNSIGNED #(.width(1), .n(11)) u_pad_1283 (
        .y(_WTEMP_172),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(11)) u_mux_1284 (
        .y(_T_599),
        .sel(_T_594),
        .a(_T_597),
        .b(_WTEMP_172)
    );
    wire _T_600;
    BITS #(.width(26), .high(24), .low(24)) bits_1285 (
        .y(_T_600),
        .in(sigY3)
    );
    wire [10:0] _T_602;
    wire [10:0] _WTEMP_173;
    PAD_UNSIGNED #(.width(1), .n(11)) u_pad_1286 (
        .y(_WTEMP_173),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(11)) u_mux_1287 (
        .y(_T_602),
        .sel(_T_600),
        .a(sExpX3),
        .b(_WTEMP_173)
    );
    wire [10:0] _T_603;
    BITWISEOR #(.width(11)) bitwiseor_1288 (
        .y(_T_603),
        .a(_T_599),
        .b(_T_602)
    );
    wire [1:0] _T_604;
    BITS #(.width(26), .high(25), .low(24)) bits_1289 (
        .y(_T_604),
        .in(sigY3)
    );
    wire _T_606;
    wire [1:0] _WTEMP_174;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_1290 (
        .y(_WTEMP_174),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(2)) u_eq_1291 (
        .y(_T_606),
        .a(_T_604),
        .b(_WTEMP_174)
    );
    wire [11:0] _T_608;
    wire [10:0] _WTEMP_175;
    PAD_UNSIGNED #(.width(1), .n(11)) u_pad_1292 (
        .y(_WTEMP_175),
        .in(1'h1)
    );
    SUB_UNSIGNED #(.width(11)) u_sub_1293 (
        .y(_T_608),
        .a(sExpX3),
        .b(_WTEMP_175)
    );
    wire [11:0] _T_609;
    ASUINT #(.width(12)) asuint_1294 (
        .y(_T_609),
        .in(_T_608)
    );
    wire [10:0] _T_610;
    TAIL #(.width(12), .n(1)) tail_1295 (
        .y(_T_610),
        .in(_T_609)
    );
    wire [10:0] _T_612;
    wire [10:0] _WTEMP_176;
    PAD_UNSIGNED #(.width(1), .n(11)) u_pad_1296 (
        .y(_WTEMP_176),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(11)) u_mux_1297 (
        .y(_T_612),
        .sel(_T_606),
        .a(_T_610),
        .b(_WTEMP_176)
    );
    wire [10:0] sExpY;
    BITWISEOR #(.width(11)) bitwiseor_1298 (
        .y(sExpY),
        .a(_T_603),
        .b(_T_612)
    );
    wire [8:0] expY;
    BITS #(.width(11), .high(8), .low(0)) bits_1299 (
        .y(expY),
        .in(sExpY)
    );
    wire [22:0] _T_613;
    BITS #(.width(26), .high(22), .low(0)) bits_1300 (
        .y(_T_613),
        .in(sigY3)
    );
    wire [22:0] _T_614;
    BITS #(.width(26), .high(23), .low(1)) bits_1301 (
        .y(_T_614),
        .in(sigY3)
    );
    wire [22:0] fractY;
    MUX_UNSIGNED #(.width(23)) u_mux_1302 (
        .y(fractY),
        .sel(sigX3Shift1),
        .a(_T_613),
        .b(_T_614)
    );
    wire [2:0] _T_615;
    BITS #(.width(11), .high(9), .low(7)) bits_1303 (
        .y(_T_615),
        .in(sExpY)
    );
    wire overflowY;
    wire [2:0] _WTEMP_177;
    PAD_UNSIGNED #(.width(2), .n(3)) u_pad_1304 (
        .y(_WTEMP_177),
        .in(2'h3)
    );
    EQ_UNSIGNED #(.width(3)) u_eq_1305 (
        .y(overflowY),
        .a(_T_615),
        .b(_WTEMP_177)
    );
    wire _T_618;
    EQ_UNSIGNED #(.width(1)) u_eq_1306 (
        .y(_T_618),
        .a(isZeroY),
        .b(1'h0)
    );
    wire _T_619;
    BITS #(.width(11), .high(9), .low(9)) bits_1307 (
        .y(_T_619),
        .in(sExpY)
    );
    wire [8:0] _T_620;
    BITS #(.width(11), .high(8), .low(0)) bits_1308 (
        .y(_T_620),
        .in(sExpY)
    );
    wire _T_622;
    wire [8:0] _WTEMP_178;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_1309 (
        .y(_WTEMP_178),
        .in(7'h6B)
    );
    LT_UNSIGNED #(.width(9)) u_lt_1310 (
        .y(_T_622),
        .a(_T_620),
        .b(_WTEMP_178)
    );
    wire _T_623;
    BITWISEOR #(.width(1)) bitwiseor_1311 (
        .y(_T_623),
        .a(_T_619),
        .b(_T_622)
    );
    wire totalUnderflowY;
    BITWISEAND #(.width(1)) bitwiseand_1312 (
        .y(totalUnderflowY),
        .a(_T_618),
        .b(_T_623)
    );
    wire _T_624;
    BITS #(.width(11), .high(10), .low(10)) bits_1313 (
        .y(_T_624),
        .in(sExpX3)
    );
    wire [7:0] _T_627;
    MUX_UNSIGNED #(.width(8)) u_mux_1314 (
        .y(_T_627),
        .sel(sigX3Shift1),
        .a(8'h82),
        .b(8'h81)
    );
    wire _T_628;
    wire [9:0] _WTEMP_179;
    PAD_UNSIGNED #(.width(8), .n(10)) u_pad_1315 (
        .y(_WTEMP_179),
        .in(_T_627)
    );
    LEQ_UNSIGNED #(.width(10)) u_leq_1316 (
        .y(_T_628),
        .a(sExpX3_13),
        .b(_WTEMP_179)
    );
    wire _T_629;
    BITWISEOR #(.width(1)) bitwiseor_1317 (
        .y(_T_629),
        .a(_T_624),
        .b(_T_628)
    );
    wire underflowY;
    BITWISEAND #(.width(1)) bitwiseand_1318 (
        .y(underflowY),
        .a(inexactY),
        .b(_T_629)
    );
    wire _T_630;
    BITWISEAND #(.width(1)) bitwiseand_1319 (
        .y(_T_630),
        .a(roundingMode_min),
        .b(signY)
    );
    wire _T_632;
    EQ_UNSIGNED #(.width(1)) u_eq_1320 (
        .y(_T_632),
        .a(signY),
        .b(1'h0)
    );
    wire _T_633;
    BITWISEAND #(.width(1)) bitwiseand_1321 (
        .y(_T_633),
        .a(roundingMode_max),
        .b(_T_632)
    );
    wire roundMagUp;
    BITWISEOR #(.width(1)) bitwiseor_1322 (
        .y(roundMagUp),
        .a(_T_630),
        .b(_T_633)
    );
    wire overflowY_roundMagUp;
    BITWISEOR #(.width(1)) bitwiseor_1323 (
        .y(overflowY_roundMagUp),
        .a(roundingMode_nearest_even),
        .b(roundMagUp)
    );
    wire mulSpecial;
    BITWISEOR #(.width(1)) bitwiseor_1324 (
        .y(mulSpecial),
        .a(isSpecialA),
        .b(isSpecialB)
    );
    wire addSpecial;
    BITWISEOR #(.width(1)) bitwiseor_1325 (
        .y(addSpecial),
        .a(mulSpecial),
        .b(isSpecialC)
    );
    wire notSpecial_addZeros;
    BITWISEAND #(.width(1)) bitwiseand_1326 (
        .y(notSpecial_addZeros),
        .a(io_fromPreMul_isZeroProd),
        .b(isZeroC)
    );
    wire _T_635;
    EQ_UNSIGNED #(.width(1)) u_eq_1327 (
        .y(_T_635),
        .a(addSpecial),
        .b(1'h0)
    );
    wire _T_637;
    EQ_UNSIGNED #(.width(1)) u_eq_1328 (
        .y(_T_637),
        .a(notSpecial_addZeros),
        .b(1'h0)
    );
    wire commonCase;
    BITWISEAND #(.width(1)) bitwiseand_1329 (
        .y(commonCase),
        .a(_T_635),
        .b(_T_637)
    );
    wire _T_638;
    BITWISEAND #(.width(1)) bitwiseand_1330 (
        .y(_T_638),
        .a(isInfA),
        .b(isZeroB)
    );
    wire _T_639;
    BITWISEAND #(.width(1)) bitwiseand_1331 (
        .y(_T_639),
        .a(isZeroA),
        .b(isInfB)
    );
    wire _T_640;
    BITWISEOR #(.width(1)) bitwiseor_1332 (
        .y(_T_640),
        .a(_T_638),
        .b(_T_639)
    );
    wire _T_642;
    EQ_UNSIGNED #(.width(1)) u_eq_1333 (
        .y(_T_642),
        .a(isNaNA),
        .b(1'h0)
    );
    wire _T_644;
    EQ_UNSIGNED #(.width(1)) u_eq_1334 (
        .y(_T_644),
        .a(isNaNB),
        .b(1'h0)
    );
    wire _T_645;
    BITWISEAND #(.width(1)) bitwiseand_1335 (
        .y(_T_645),
        .a(_T_642),
        .b(_T_644)
    );
    wire _T_646;
    BITWISEOR #(.width(1)) bitwiseor_1336 (
        .y(_T_646),
        .a(isInfA),
        .b(isInfB)
    );
    wire _T_647;
    BITWISEAND #(.width(1)) bitwiseand_1337 (
        .y(_T_647),
        .a(_T_645),
        .b(_T_646)
    );
    wire _T_648;
    BITWISEAND #(.width(1)) bitwiseand_1338 (
        .y(_T_648),
        .a(_T_647),
        .b(isInfC)
    );
    wire _T_649;
    BITWISEAND #(.width(1)) bitwiseand_1339 (
        .y(_T_649),
        .a(_T_648),
        .b(doSubMags)
    );
    wire notSigNaN_invalid;
    BITWISEOR #(.width(1)) bitwiseor_1340 (
        .y(notSigNaN_invalid),
        .a(_T_640),
        .b(_T_649)
    );
    wire _T_650;
    BITWISEOR #(.width(1)) bitwiseor_1341 (
        .y(_T_650),
        .a(isSigNaNA),
        .b(isSigNaNB)
    );
    wire _T_651;
    BITWISEOR #(.width(1)) bitwiseor_1342 (
        .y(_T_651),
        .a(_T_650),
        .b(isSigNaNC)
    );
    wire invalid;
    BITWISEOR #(.width(1)) bitwiseor_1343 (
        .y(invalid),
        .a(_T_651),
        .b(notSigNaN_invalid)
    );
    wire overflow;
    BITWISEAND #(.width(1)) bitwiseand_1344 (
        .y(overflow),
        .a(commonCase),
        .b(overflowY)
    );
    wire underflow;
    BITWISEAND #(.width(1)) bitwiseand_1345 (
        .y(underflow),
        .a(commonCase),
        .b(underflowY)
    );
    wire _T_652;
    BITWISEAND #(.width(1)) bitwiseand_1346 (
        .y(_T_652),
        .a(commonCase),
        .b(inexactY)
    );
    wire inexact;
    BITWISEOR #(.width(1)) bitwiseor_1347 (
        .y(inexact),
        .a(overflow),
        .b(_T_652)
    );
    wire _T_653;
    BITWISEOR #(.width(1)) bitwiseor_1348 (
        .y(_T_653),
        .a(notSpecial_addZeros),
        .b(isZeroY)
    );
    wire notSpecial_isZeroOut;
    BITWISEOR #(.width(1)) bitwiseor_1349 (
        .y(notSpecial_isZeroOut),
        .a(_T_653),
        .b(totalUnderflowY)
    );
    wire _T_654;
    BITWISEAND #(.width(1)) bitwiseand_1350 (
        .y(_T_654),
        .a(commonCase),
        .b(totalUnderflowY)
    );
    wire pegMinFiniteMagOut;
    BITWISEAND #(.width(1)) bitwiseand_1351 (
        .y(pegMinFiniteMagOut),
        .a(_T_654),
        .b(roundMagUp)
    );
    wire _T_656;
    EQ_UNSIGNED #(.width(1)) u_eq_1352 (
        .y(_T_656),
        .a(overflowY_roundMagUp),
        .b(1'h0)
    );
    wire pegMaxFiniteMagOut;
    BITWISEAND #(.width(1)) bitwiseand_1353 (
        .y(pegMaxFiniteMagOut),
        .a(overflow),
        .b(_T_656)
    );
    wire _T_657;
    BITWISEOR #(.width(1)) bitwiseor_1354 (
        .y(_T_657),
        .a(isInfA),
        .b(isInfB)
    );
    wire _T_658;
    BITWISEOR #(.width(1)) bitwiseor_1355 (
        .y(_T_658),
        .a(_T_657),
        .b(isInfC)
    );
    wire _T_659;
    BITWISEAND #(.width(1)) bitwiseand_1356 (
        .y(_T_659),
        .a(overflow),
        .b(overflowY_roundMagUp)
    );
    wire notNaN_isInfOut;
    BITWISEOR #(.width(1)) bitwiseor_1357 (
        .y(notNaN_isInfOut),
        .a(_T_658),
        .b(_T_659)
    );
    wire _T_660;
    BITWISEOR #(.width(1)) bitwiseor_1358 (
        .y(_T_660),
        .a(isNaNA),
        .b(isNaNB)
    );
    wire _T_661;
    BITWISEOR #(.width(1)) bitwiseor_1359 (
        .y(_T_661),
        .a(_T_660),
        .b(isNaNC)
    );
    wire isNaNOut;
    BITWISEOR #(.width(1)) bitwiseor_1360 (
        .y(isNaNOut),
        .a(_T_661),
        .b(notSigNaN_invalid)
    );
    wire _T_663;
    EQ_UNSIGNED #(.width(1)) u_eq_1361 (
        .y(_T_663),
        .a(doSubMags),
        .b(1'h0)
    );
    wire _T_664;
    BITWISEAND #(.width(1)) bitwiseand_1362 (
        .y(_T_664),
        .a(_T_663),
        .b(io_fromPreMul_opSignC)
    );
    wire _T_666;
    EQ_UNSIGNED #(.width(1)) u_eq_1363 (
        .y(_T_666),
        .a(isSpecialC),
        .b(1'h0)
    );
    wire _T_667;
    BITWISEAND #(.width(1)) bitwiseand_1364 (
        .y(_T_667),
        .a(mulSpecial),
        .b(_T_666)
    );
    wire _T_668;
    BITWISEAND #(.width(1)) bitwiseand_1365 (
        .y(_T_668),
        .a(_T_667),
        .b(io_fromPreMul_signProd)
    );
    wire _T_669;
    BITWISEOR #(.width(1)) bitwiseor_1366 (
        .y(_T_669),
        .a(_T_664),
        .b(_T_668)
    );
    wire _T_671;
    EQ_UNSIGNED #(.width(1)) u_eq_1367 (
        .y(_T_671),
        .a(mulSpecial),
        .b(1'h0)
    );
    wire _T_672;
    BITWISEAND #(.width(1)) bitwiseand_1368 (
        .y(_T_672),
        .a(_T_671),
        .b(isSpecialC)
    );
    wire _T_673;
    BITWISEAND #(.width(1)) bitwiseand_1369 (
        .y(_T_673),
        .a(_T_672),
        .b(io_fromPreMul_opSignC)
    );
    wire _T_674;
    BITWISEOR #(.width(1)) bitwiseor_1370 (
        .y(_T_674),
        .a(_T_669),
        .b(_T_673)
    );
    wire _T_676;
    EQ_UNSIGNED #(.width(1)) u_eq_1371 (
        .y(_T_676),
        .a(mulSpecial),
        .b(1'h0)
    );
    wire _T_677;
    BITWISEAND #(.width(1)) bitwiseand_1372 (
        .y(_T_677),
        .a(_T_676),
        .b(notSpecial_addZeros)
    );
    wire _T_678;
    BITWISEAND #(.width(1)) bitwiseand_1373 (
        .y(_T_678),
        .a(_T_677),
        .b(doSubMags)
    );
    wire _T_679;
    BITWISEAND #(.width(1)) bitwiseand_1374 (
        .y(_T_679),
        .a(_T_678),
        .b(signZeroNotEqOpSigns)
    );
    wire uncommonCaseSignOut;
    BITWISEOR #(.width(1)) bitwiseor_1375 (
        .y(uncommonCaseSignOut),
        .a(_T_674),
        .b(_T_679)
    );
    wire _T_681;
    EQ_UNSIGNED #(.width(1)) u_eq_1376 (
        .y(_T_681),
        .a(isNaNOut),
        .b(1'h0)
    );
    wire _T_682;
    BITWISEAND #(.width(1)) bitwiseand_1377 (
        .y(_T_682),
        .a(_T_681),
        .b(uncommonCaseSignOut)
    );
    wire _T_683;
    BITWISEAND #(.width(1)) bitwiseand_1378 (
        .y(_T_683),
        .a(commonCase),
        .b(signY)
    );
    wire signOut;
    BITWISEOR #(.width(1)) bitwiseor_1379 (
        .y(signOut),
        .a(_T_682),
        .b(_T_683)
    );
    wire [8:0] _T_686;
    MUX_UNSIGNED #(.width(9)) u_mux_1380 (
        .y(_T_686),
        .sel(notSpecial_isZeroOut),
        .a(9'h1C0),
        .b(9'h0)
    );
    wire [8:0] _T_687;
    BITWISENOT #(.width(9)) bitwisenot_1381 (
        .y(_T_687),
        .in(_T_686)
    );
    wire [8:0] _T_688;
    BITWISEAND #(.width(9)) bitwiseand_1382 (
        .y(_T_688),
        .a(expY),
        .b(_T_687)
    );
    wire [8:0] _T_690;
    assign _T_690 = 9'h194;
    wire [8:0] _T_692;
    MUX_UNSIGNED #(.width(9)) u_mux_1383 (
        .y(_T_692),
        .sel(pegMinFiniteMagOut),
        .a(_T_690),
        .b(9'h0)
    );
    wire [8:0] _T_693;
    BITWISENOT #(.width(9)) bitwisenot_1384 (
        .y(_T_693),
        .in(_T_692)
    );
    wire [8:0] _T_694;
    BITWISEAND #(.width(9)) bitwiseand_1385 (
        .y(_T_694),
        .a(_T_688),
        .b(_T_693)
    );
    wire [8:0] _T_697;
    MUX_UNSIGNED #(.width(9)) u_mux_1386 (
        .y(_T_697),
        .sel(pegMaxFiniteMagOut),
        .a(9'h80),
        .b(9'h0)
    );
    wire [8:0] _T_698;
    BITWISENOT #(.width(9)) bitwisenot_1387 (
        .y(_T_698),
        .in(_T_697)
    );
    wire [8:0] _T_699;
    BITWISEAND #(.width(9)) bitwiseand_1388 (
        .y(_T_699),
        .a(_T_694),
        .b(_T_698)
    );
    wire [8:0] _T_702;
    wire [8:0] _WTEMP_180;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_1389 (
        .y(_WTEMP_180),
        .in(7'h40)
    );
    MUX_UNSIGNED #(.width(9)) u_mux_1390 (
        .y(_T_702),
        .sel(notNaN_isInfOut),
        .a(_WTEMP_180),
        .b(9'h0)
    );
    wire [8:0] _T_703;
    BITWISENOT #(.width(9)) bitwisenot_1391 (
        .y(_T_703),
        .in(_T_702)
    );
    wire [8:0] _T_704;
    BITWISEAND #(.width(9)) bitwiseand_1392 (
        .y(_T_704),
        .a(_T_699),
        .b(_T_703)
    );
    wire [8:0] _T_707;
    wire [8:0] _WTEMP_181;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_1393 (
        .y(_WTEMP_181),
        .in(7'h6B)
    );
    MUX_UNSIGNED #(.width(9)) u_mux_1394 (
        .y(_T_707),
        .sel(pegMinFiniteMagOut),
        .a(_WTEMP_181),
        .b(9'h0)
    );
    wire [8:0] _T_708;
    BITWISEOR #(.width(9)) bitwiseor_1395 (
        .y(_T_708),
        .a(_T_704),
        .b(_T_707)
    );
    wire [8:0] _T_711;
    MUX_UNSIGNED #(.width(9)) u_mux_1396 (
        .y(_T_711),
        .sel(pegMaxFiniteMagOut),
        .a(9'h17F),
        .b(9'h0)
    );
    wire [8:0] _T_712;
    BITWISEOR #(.width(9)) bitwiseor_1397 (
        .y(_T_712),
        .a(_T_708),
        .b(_T_711)
    );
    wire [8:0] _T_715;
    MUX_UNSIGNED #(.width(9)) u_mux_1398 (
        .y(_T_715),
        .sel(notNaN_isInfOut),
        .a(9'h180),
        .b(9'h0)
    );
    wire [8:0] _T_716;
    BITWISEOR #(.width(9)) bitwiseor_1399 (
        .y(_T_716),
        .a(_T_712),
        .b(_T_715)
    );
    wire [8:0] _T_719;
    MUX_UNSIGNED #(.width(9)) u_mux_1400 (
        .y(_T_719),
        .sel(isNaNOut),
        .a(9'h1C0),
        .b(9'h0)
    );
    wire [8:0] expOut;
    BITWISEOR #(.width(9)) bitwiseor_1401 (
        .y(expOut),
        .a(_T_716),
        .b(_T_719)
    );
    wire _T_720;
    BITWISEAND #(.width(1)) bitwiseand_1402 (
        .y(_T_720),
        .a(totalUnderflowY),
        .b(roundMagUp)
    );
    wire _T_721;
    BITWISEOR #(.width(1)) bitwiseor_1403 (
        .y(_T_721),
        .a(_T_720),
        .b(isNaNOut)
    );
    wire [22:0] _T_723;
    assign _T_723 = 23'h400000;
    wire [22:0] _T_725;
    wire [22:0] _WTEMP_182;
    PAD_UNSIGNED #(.width(1), .n(23)) u_pad_1404 (
        .y(_WTEMP_182),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(23)) u_mux_1405 (
        .y(_T_725),
        .sel(isNaNOut),
        .a(_T_723),
        .b(_WTEMP_182)
    );
    wire [22:0] _T_726;
    MUX_UNSIGNED #(.width(23)) u_mux_1406 (
        .y(_T_726),
        .sel(_T_721),
        .a(_T_725),
        .b(fractY)
    );
    wire _T_727;
    BITS #(.width(1), .high(0), .low(0)) bits_1407 (
        .y(_T_727),
        .in(pegMaxFiniteMagOut)
    );
    wire [22:0] _T_730;
    MUX_UNSIGNED #(.width(23)) u_mux_1408 (
        .y(_T_730),
        .sel(_T_727),
        .a(23'h7FFFFF),
        .b(23'h0)
    );
    wire [22:0] fractOut;
    BITWISEOR #(.width(23)) bitwiseor_1409 (
        .y(fractOut),
        .a(_T_726),
        .b(_T_730)
    );
    wire [9:0] _T_731;
    CAT #(.width_a(1), .width_b(9)) cat_1410 (
        .y(_T_731),
        .a(signOut),
        .b(expOut)
    );
    wire [32:0] _T_732;
    CAT #(.width_a(10), .width_b(23)) cat_1411 (
        .y(_T_732),
        .a(_T_731),
        .b(fractOut)
    );
    wire [1:0] _T_734;
    CAT #(.width_a(1), .width_b(1)) cat_1412 (
        .y(_T_734),
        .a(underflow),
        .b(inexact)
    );
    wire [1:0] _T_735;
    CAT #(.width_a(1), .width_b(1)) cat_1413 (
        .y(_T_735),
        .a(invalid),
        .b(1'h0)
    );
    wire [2:0] _T_736;
    CAT #(.width_a(2), .width_b(1)) cat_1414 (
        .y(_T_736),
        .a(_T_735),
        .b(overflow)
    );
    wire [4:0] _T_737;
    CAT #(.width_a(3), .width_b(2)) cat_1415 (
        .y(_T_737),
        .a(_T_736),
        .b(_T_734)
    );
    assign io_exceptionFlags = _T_737;
    assign io_out = _T_732;
endmodule //MulAddRecFN_postMul
module DSHR_UNSIGNED(y, in, n);
    parameter width_in = 4;
    parameter width_n = 2;
    output [width_in-1:0] y;
    input [width_in-1:0] in;
    input [width_n-1:0] n;
    assign y = in >> n;
endmodule // DSHR_UNSIGNED
module LEQ_UNSIGNED(y, a, b);
    parameter width = 4;
    output y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a <= b;
endmodule // LEQ_UNSIGNED
module MUL2_UNSIGNED(y, a, b);
    parameter width_a = 4;
    parameter width_b = 4;
    output [width_a+width_b-1:0] y;
    input [width_a-1:0] a;
    input [width_b-1:0] b;
    assign y = a * b;
endmodule // MUL2_UNSIGNED
module FPToInt(
    input clock,
    input reset,
    input io_in_valid,
    input [4:0] io_in_bits_cmd,
    input io_in_bits_ldst,
    input io_in_bits_wen,
    input io_in_bits_ren1,
    input io_in_bits_ren2,
    input io_in_bits_ren3,
    input io_in_bits_swap12,
    input io_in_bits_swap23,
    input io_in_bits_single,
    input io_in_bits_fromint,
    input io_in_bits_toint,
    input io_in_bits_fastpipe,
    input io_in_bits_fma,
    input io_in_bits_div,
    input io_in_bits_sqrt,
    input io_in_bits_wflags,
    input [2:0] io_in_bits_rm,
    input [1:0] io_in_bits_typ,
    input [64:0] io_in_bits_in1,
    input [64:0] io_in_bits_in2,
    input [64:0] io_in_bits_in3,
    output [4:0] io_as_double_cmd,
    output io_as_double_ldst,
    output io_as_double_wen,
    output io_as_double_ren1,
    output io_as_double_ren2,
    output io_as_double_ren3,
    output io_as_double_swap12,
    output io_as_double_swap23,
    output io_as_double_single,
    output io_as_double_fromint,
    output io_as_double_toint,
    output io_as_double_fastpipe,
    output io_as_double_fma,
    output io_as_double_div,
    output io_as_double_sqrt,
    output io_as_double_wflags,
    output [2:0] io_as_double_rm,
    output [1:0] io_as_double_typ,
    output [64:0] io_as_double_in1,
    output [64:0] io_as_double_in2,
    output [64:0] io_as_double_in3,
    output io_out_valid,
    output io_out_bits_lt,
    output [63:0] io_out_bits_store,
    output [63:0] io_out_bits_toint,
    output [4:0] io_out_bits_exc
);
    wire [4:0] _in_cmd__q;
    wire [4:0] _in_cmd__d;
    DFF_POSCLK #(.width(5)) in_cmd (
        .q(_in_cmd__q),
        .d(_in_cmd__d),
        .clk(clock)
    );
    wire _in_ldst__q;
    wire _in_ldst__d;
    DFF_POSCLK #(.width(1)) in_ldst (
        .q(_in_ldst__q),
        .d(_in_ldst__d),
        .clk(clock)
    );
    wire _in_wen__q;
    wire _in_wen__d;
    DFF_POSCLK #(.width(1)) in_wen (
        .q(_in_wen__q),
        .d(_in_wen__d),
        .clk(clock)
    );
    wire _in_ren1__q;
    wire _in_ren1__d;
    DFF_POSCLK #(.width(1)) in_ren1 (
        .q(_in_ren1__q),
        .d(_in_ren1__d),
        .clk(clock)
    );
    wire _in_ren2__q;
    wire _in_ren2__d;
    DFF_POSCLK #(.width(1)) in_ren2 (
        .q(_in_ren2__q),
        .d(_in_ren2__d),
        .clk(clock)
    );
    wire _in_ren3__q;
    wire _in_ren3__d;
    DFF_POSCLK #(.width(1)) in_ren3 (
        .q(_in_ren3__q),
        .d(_in_ren3__d),
        .clk(clock)
    );
    wire _in_swap12__q;
    wire _in_swap12__d;
    DFF_POSCLK #(.width(1)) in_swap12 (
        .q(_in_swap12__q),
        .d(_in_swap12__d),
        .clk(clock)
    );
    wire _in_swap23__q;
    wire _in_swap23__d;
    DFF_POSCLK #(.width(1)) in_swap23 (
        .q(_in_swap23__q),
        .d(_in_swap23__d),
        .clk(clock)
    );
    wire _in_single__q;
    wire _in_single__d;
    DFF_POSCLK #(.width(1)) in_single (
        .q(_in_single__q),
        .d(_in_single__d),
        .clk(clock)
    );
    wire _in_fromint__q;
    wire _in_fromint__d;
    DFF_POSCLK #(.width(1)) in_fromint (
        .q(_in_fromint__q),
        .d(_in_fromint__d),
        .clk(clock)
    );
    wire _in_toint__q;
    wire _in_toint__d;
    DFF_POSCLK #(.width(1)) in_toint (
        .q(_in_toint__q),
        .d(_in_toint__d),
        .clk(clock)
    );
    wire _in_fastpipe__q;
    wire _in_fastpipe__d;
    DFF_POSCLK #(.width(1)) in_fastpipe (
        .q(_in_fastpipe__q),
        .d(_in_fastpipe__d),
        .clk(clock)
    );
    wire _in_fma__q;
    wire _in_fma__d;
    DFF_POSCLK #(.width(1)) in_fma (
        .q(_in_fma__q),
        .d(_in_fma__d),
        .clk(clock)
    );
    wire _in_div__q;
    wire _in_div__d;
    DFF_POSCLK #(.width(1)) in_div (
        .q(_in_div__q),
        .d(_in_div__d),
        .clk(clock)
    );
    wire _in_sqrt__q;
    wire _in_sqrt__d;
    DFF_POSCLK #(.width(1)) in_sqrt (
        .q(_in_sqrt__q),
        .d(_in_sqrt__d),
        .clk(clock)
    );
    wire _in_wflags__q;
    wire _in_wflags__d;
    DFF_POSCLK #(.width(1)) in_wflags (
        .q(_in_wflags__q),
        .d(_in_wflags__d),
        .clk(clock)
    );
    wire [2:0] _in_rm__q;
    wire [2:0] _in_rm__d;
    DFF_POSCLK #(.width(3)) in_rm (
        .q(_in_rm__q),
        .d(_in_rm__d),
        .clk(clock)
    );
    wire [1:0] _in_typ__q;
    wire [1:0] _in_typ__d;
    DFF_POSCLK #(.width(2)) in_typ (
        .q(_in_typ__q),
        .d(_in_typ__d),
        .clk(clock)
    );
    wire [64:0] _in_in1__q;
    wire [64:0] _in_in1__d;
    DFF_POSCLK #(.width(65)) in_in1 (
        .q(_in_in1__q),
        .d(_in_in1__d),
        .clk(clock)
    );
    wire [64:0] _in_in2__q;
    wire [64:0] _in_in2__d;
    DFF_POSCLK #(.width(65)) in_in2 (
        .q(_in_in2__q),
        .d(_in_in2__d),
        .clk(clock)
    );
    wire [64:0] _in_in3__q;
    wire [64:0] _in_in3__d;
    DFF_POSCLK #(.width(65)) in_in3 (
        .q(_in_in3__q),
        .d(_in_in3__d),
        .clk(clock)
    );
    wire _valid__q;
    wire _valid__d;
    DFF_POSCLK #(.width(1)) valid (
        .q(_valid__q),
        .d(_valid__d),
        .clk(clock)
    );
    wire _T_224;
    EQ_UNSIGNED #(.width(1)) u_eq_1457 (
        .y(_T_224),
        .a(io_in_bits_ldst),
        .b(1'h0)
    );
    wire _T_225;
    BITWISEAND #(.width(1)) bitwiseand_1458 (
        .y(_T_225),
        .a(io_in_bits_single),
        .b(_T_224)
    );
    wire [4:0] _T_228;
    wire [4:0] _WTEMP_187;
    PAD_UNSIGNED #(.width(4), .n(5)) u_pad_1459 (
        .y(_WTEMP_187),
        .in(4'hC)
    );
    BITWISEAND #(.width(5)) bitwiseand_1460 (
        .y(_T_228),
        .a(io_in_bits_cmd),
        .b(_WTEMP_187)
    );
    wire _T_229;
    wire [4:0] _WTEMP_188;
    PAD_UNSIGNED #(.width(4), .n(5)) u_pad_1461 (
        .y(_WTEMP_188),
        .in(4'hC)
    );
    EQ_UNSIGNED #(.width(5)) u_eq_1462 (
        .y(_T_229),
        .a(_WTEMP_188),
        .b(_T_228)
    );
    wire _T_231;
    EQ_UNSIGNED #(.width(1)) u_eq_1463 (
        .y(_T_231),
        .a(_T_229),
        .b(1'h0)
    );
    wire _T_232;
    BITWISEAND #(.width(1)) bitwiseand_1464 (
        .y(_T_232),
        .a(_T_225),
        .b(_T_231)
    );
    wire _T_233;
    BITS #(.width(65), .high(32), .low(32)) bits_1465 (
        .y(_T_233),
        .in(io_in_bits_in1)
    );
    wire [22:0] _T_234;
    BITS #(.width(65), .high(22), .low(0)) bits_1466 (
        .y(_T_234),
        .in(io_in_bits_in1)
    );
    wire [8:0] _T_235;
    BITS #(.width(65), .high(31), .low(23)) bits_1467 (
        .y(_T_235),
        .in(io_in_bits_in1)
    );
    wire [75:0] _T_236;
    SHL_UNSIGNED #(.width(23), .n(53)) u_shl_1468 (
        .y(_T_236),
        .in(_T_234)
    );
    wire [51:0] _T_237;
    SHR_UNSIGNED #(.width(76), .n(24)) u_shr_1469 (
        .y(_T_237),
        .in(_T_236)
    );
    wire [2:0] _T_238;
    BITS #(.width(9), .high(8), .low(6)) bits_1470 (
        .y(_T_238),
        .in(_T_235)
    );
    wire [12:0] _T_240;
    wire [11:0] _WTEMP_189;
    PAD_UNSIGNED #(.width(9), .n(12)) u_pad_1471 (
        .y(_WTEMP_189),
        .in(_T_235)
    );
    ADD_UNSIGNED #(.width(12)) u_add_1472 (
        .y(_T_240),
        .a(_WTEMP_189),
        .b(12'h800)
    );
    wire [11:0] _T_241;
    TAIL #(.width(13), .n(1)) tail_1473 (
        .y(_T_241),
        .in(_T_240)
    );
    wire [12:0] _T_243;
    wire [11:0] _WTEMP_190;
    PAD_UNSIGNED #(.width(9), .n(12)) u_pad_1474 (
        .y(_WTEMP_190),
        .in(9'h100)
    );
    SUB_UNSIGNED #(.width(12)) u_sub_1475 (
        .y(_T_243),
        .a(_T_241),
        .b(_WTEMP_190)
    );
    wire [12:0] _T_244;
    ASUINT #(.width(13)) asuint_1476 (
        .y(_T_244),
        .in(_T_243)
    );
    wire [11:0] _T_245;
    TAIL #(.width(13), .n(1)) tail_1477 (
        .y(_T_245),
        .in(_T_244)
    );
    wire _T_247;
    wire [2:0] _WTEMP_191;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_1478 (
        .y(_WTEMP_191),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(3)) u_eq_1479 (
        .y(_T_247),
        .a(_T_238),
        .b(_WTEMP_191)
    );
    wire _T_249;
    GEQ_UNSIGNED #(.width(3)) u_geq_1480 (
        .y(_T_249),
        .a(_T_238),
        .b(3'h6)
    );
    wire _T_250;
    BITWISEOR #(.width(1)) bitwiseor_1481 (
        .y(_T_250),
        .a(_T_247),
        .b(_T_249)
    );
    wire [8:0] _T_251;
    BITS #(.width(12), .high(8), .low(0)) bits_1482 (
        .y(_T_251),
        .in(_T_245)
    );
    wire [11:0] _T_252;
    CAT #(.width_a(3), .width_b(9)) cat_1483 (
        .y(_T_252),
        .a(_T_238),
        .b(_T_251)
    );
    wire [11:0] _T_253;
    BITS #(.width(12), .high(11), .low(0)) bits_1484 (
        .y(_T_253),
        .in(_T_245)
    );
    wire [11:0] _T_254;
    MUX_UNSIGNED #(.width(12)) u_mux_1485 (
        .y(_T_254),
        .sel(_T_250),
        .a(_T_252),
        .b(_T_253)
    );
    wire [12:0] _T_255;
    CAT #(.width_a(1), .width_b(12)) cat_1486 (
        .y(_T_255),
        .a(_T_233),
        .b(_T_254)
    );
    wire [64:0] _T_256;
    CAT #(.width_a(13), .width_b(52)) cat_1487 (
        .y(_T_256),
        .a(_T_255),
        .b(_T_237)
    );
    wire _T_257;
    BITS #(.width(65), .high(32), .low(32)) bits_1488 (
        .y(_T_257),
        .in(io_in_bits_in2)
    );
    wire [22:0] _T_258;
    BITS #(.width(65), .high(22), .low(0)) bits_1489 (
        .y(_T_258),
        .in(io_in_bits_in2)
    );
    wire [8:0] _T_259;
    BITS #(.width(65), .high(31), .low(23)) bits_1490 (
        .y(_T_259),
        .in(io_in_bits_in2)
    );
    wire [75:0] _T_260;
    SHL_UNSIGNED #(.width(23), .n(53)) u_shl_1491 (
        .y(_T_260),
        .in(_T_258)
    );
    wire [51:0] _T_261;
    SHR_UNSIGNED #(.width(76), .n(24)) u_shr_1492 (
        .y(_T_261),
        .in(_T_260)
    );
    wire [2:0] _T_262;
    BITS #(.width(9), .high(8), .low(6)) bits_1493 (
        .y(_T_262),
        .in(_T_259)
    );
    wire [12:0] _T_264;
    wire [11:0] _WTEMP_192;
    PAD_UNSIGNED #(.width(9), .n(12)) u_pad_1494 (
        .y(_WTEMP_192),
        .in(_T_259)
    );
    ADD_UNSIGNED #(.width(12)) u_add_1495 (
        .y(_T_264),
        .a(_WTEMP_192),
        .b(12'h800)
    );
    wire [11:0] _T_265;
    TAIL #(.width(13), .n(1)) tail_1496 (
        .y(_T_265),
        .in(_T_264)
    );
    wire [12:0] _T_267;
    wire [11:0] _WTEMP_193;
    PAD_UNSIGNED #(.width(9), .n(12)) u_pad_1497 (
        .y(_WTEMP_193),
        .in(9'h100)
    );
    SUB_UNSIGNED #(.width(12)) u_sub_1498 (
        .y(_T_267),
        .a(_T_265),
        .b(_WTEMP_193)
    );
    wire [12:0] _T_268;
    ASUINT #(.width(13)) asuint_1499 (
        .y(_T_268),
        .in(_T_267)
    );
    wire [11:0] _T_269;
    TAIL #(.width(13), .n(1)) tail_1500 (
        .y(_T_269),
        .in(_T_268)
    );
    wire _T_271;
    wire [2:0] _WTEMP_194;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_1501 (
        .y(_WTEMP_194),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(3)) u_eq_1502 (
        .y(_T_271),
        .a(_T_262),
        .b(_WTEMP_194)
    );
    wire _T_273;
    GEQ_UNSIGNED #(.width(3)) u_geq_1503 (
        .y(_T_273),
        .a(_T_262),
        .b(3'h6)
    );
    wire _T_274;
    BITWISEOR #(.width(1)) bitwiseor_1504 (
        .y(_T_274),
        .a(_T_271),
        .b(_T_273)
    );
    wire [8:0] _T_275;
    BITS #(.width(12), .high(8), .low(0)) bits_1505 (
        .y(_T_275),
        .in(_T_269)
    );
    wire [11:0] _T_276;
    CAT #(.width_a(3), .width_b(9)) cat_1506 (
        .y(_T_276),
        .a(_T_262),
        .b(_T_275)
    );
    wire [11:0] _T_277;
    BITS #(.width(12), .high(11), .low(0)) bits_1507 (
        .y(_T_277),
        .in(_T_269)
    );
    wire [11:0] _T_278;
    MUX_UNSIGNED #(.width(12)) u_mux_1508 (
        .y(_T_278),
        .sel(_T_274),
        .a(_T_276),
        .b(_T_277)
    );
    wire [12:0] _T_279;
    CAT #(.width_a(1), .width_b(12)) cat_1509 (
        .y(_T_279),
        .a(_T_257),
        .b(_T_278)
    );
    wire [64:0] _T_280;
    CAT #(.width_a(13), .width_b(52)) cat_1510 (
        .y(_T_280),
        .a(_T_279),
        .b(_T_261)
    );
    wire [64:0] _node_17;
    MUX_UNSIGNED #(.width(65)) u_mux_1511 (
        .y(_node_17),
        .sel(_T_232),
        .a(_T_256),
        .b(io_in_bits_in1)
    );
    wire [64:0] _node_18;
    MUX_UNSIGNED #(.width(65)) u_mux_1512 (
        .y(_node_18),
        .sel(_T_232),
        .a(_T_280),
        .b(io_in_bits_in2)
    );
    wire _T_281;
    BITS #(.width(65), .high(32), .low(32)) bits_1513 (
        .y(_T_281),
        .in(_in_in1__q)
    );
    wire [8:0] _T_282;
    BITS #(.width(65), .high(31), .low(23)) bits_1514 (
        .y(_T_282),
        .in(_in_in1__q)
    );
    wire [22:0] _T_283;
    BITS #(.width(65), .high(22), .low(0)) bits_1515 (
        .y(_T_283),
        .in(_in_in1__q)
    );
    wire [6:0] _T_284;
    BITS #(.width(9), .high(6), .low(0)) bits_1516 (
        .y(_T_284),
        .in(_T_282)
    );
    wire _T_286;
    wire [6:0] _WTEMP_195;
    PAD_UNSIGNED #(.width(2), .n(7)) u_pad_1517 (
        .y(_WTEMP_195),
        .in(2'h2)
    );
    LT_UNSIGNED #(.width(7)) u_lt_1518 (
        .y(_T_286),
        .a(_T_284),
        .b(_WTEMP_195)
    );
    wire [2:0] _T_287;
    BITS #(.width(9), .high(8), .low(6)) bits_1519 (
        .y(_T_287),
        .in(_T_282)
    );
    wire _T_289;
    wire [2:0] _WTEMP_196;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_1520 (
        .y(_WTEMP_196),
        .in(1'h1)
    );
    EQ_UNSIGNED #(.width(3)) u_eq_1521 (
        .y(_T_289),
        .a(_T_287),
        .b(_WTEMP_196)
    );
    wire [1:0] _T_290;
    BITS #(.width(9), .high(8), .low(7)) bits_1522 (
        .y(_T_290),
        .in(_T_282)
    );
    wire _T_292;
    wire [1:0] _WTEMP_197;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_1523 (
        .y(_WTEMP_197),
        .in(1'h1)
    );
    EQ_UNSIGNED #(.width(2)) u_eq_1524 (
        .y(_T_292),
        .a(_T_290),
        .b(_WTEMP_197)
    );
    wire _T_293;
    BITWISEAND #(.width(1)) bitwiseand_1525 (
        .y(_T_293),
        .a(_T_292),
        .b(_T_286)
    );
    wire _T_294;
    BITWISEOR #(.width(1)) bitwiseor_1526 (
        .y(_T_294),
        .a(_T_289),
        .b(_T_293)
    );
    wire [1:0] _T_295;
    BITS #(.width(9), .high(8), .low(7)) bits_1527 (
        .y(_T_295),
        .in(_T_282)
    );
    wire _T_297;
    wire [1:0] _WTEMP_198;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_1528 (
        .y(_WTEMP_198),
        .in(1'h1)
    );
    EQ_UNSIGNED #(.width(2)) u_eq_1529 (
        .y(_T_297),
        .a(_T_295),
        .b(_WTEMP_198)
    );
    wire _T_299;
    EQ_UNSIGNED #(.width(1)) u_eq_1530 (
        .y(_T_299),
        .a(_T_286),
        .b(1'h0)
    );
    wire _T_300;
    BITWISEAND #(.width(1)) bitwiseand_1531 (
        .y(_T_300),
        .a(_T_297),
        .b(_T_299)
    );
    wire [1:0] _T_301;
    BITS #(.width(9), .high(8), .low(7)) bits_1532 (
        .y(_T_301),
        .in(_T_282)
    );
    wire _T_303;
    EQ_UNSIGNED #(.width(2)) u_eq_1533 (
        .y(_T_303),
        .a(_T_301),
        .b(2'h2)
    );
    wire _T_304;
    BITWISEOR #(.width(1)) bitwiseor_1534 (
        .y(_T_304),
        .a(_T_300),
        .b(_T_303)
    );
    wire [1:0] _T_305;
    BITS #(.width(9), .high(8), .low(7)) bits_1535 (
        .y(_T_305),
        .in(_T_282)
    );
    wire _T_307;
    EQ_UNSIGNED #(.width(2)) u_eq_1536 (
        .y(_T_307),
        .a(_T_305),
        .b(2'h3)
    );
    wire _T_308;
    BITS #(.width(9), .high(6), .low(6)) bits_1537 (
        .y(_T_308),
        .in(_T_282)
    );
    wire _T_309;
    BITWISEAND #(.width(1)) bitwiseand_1538 (
        .y(_T_309),
        .a(_T_307),
        .b(_T_308)
    );
    wire [4:0] _T_311;
    BITS #(.width(9), .high(4), .low(0)) bits_1539 (
        .y(_T_311),
        .in(_T_282)
    );
    wire [5:0] _T_312;
    wire [4:0] _WTEMP_199;
    PAD_UNSIGNED #(.width(2), .n(5)) u_pad_1540 (
        .y(_WTEMP_199),
        .in(2'h2)
    );
    SUB_UNSIGNED #(.width(5)) u_sub_1541 (
        .y(_T_312),
        .a(_WTEMP_199),
        .b(_T_311)
    );
    wire [5:0] _T_313;
    ASUINT #(.width(6)) asuint_1542 (
        .y(_T_313),
        .in(_T_312)
    );
    wire [4:0] _T_314;
    TAIL #(.width(6), .n(1)) tail_1543 (
        .y(_T_314),
        .in(_T_313)
    );
    wire [23:0] _T_316;
    CAT #(.width_a(1), .width_b(23)) cat_1544 (
        .y(_T_316),
        .a(1'h1),
        .b(_T_283)
    );
    wire [23:0] _T_317;
    DSHR_UNSIGNED #(.width_in(24), .width_n(5)) u_dshr_1545 (
        .y(_T_317),
        .in(_T_316),
        .n(_T_314)
    );
    wire [22:0] _T_318;
    BITS #(.width(24), .high(22), .low(0)) bits_1546 (
        .y(_T_318),
        .in(_T_317)
    );
    wire [7:0] _T_319;
    BITS #(.width(9), .high(7), .low(0)) bits_1547 (
        .y(_T_319),
        .in(_T_282)
    );
    wire [8:0] _T_321;
    SUB_UNSIGNED #(.width(8)) u_sub_1548 (
        .y(_T_321),
        .a(_T_319),
        .b(8'h81)
    );
    wire [8:0] _T_322;
    ASUINT #(.width(9)) asuint_1549 (
        .y(_T_322),
        .in(_T_321)
    );
    wire [7:0] _T_323;
    TAIL #(.width(9), .n(1)) tail_1550 (
        .y(_T_323),
        .in(_T_322)
    );
    wire _T_324;
    BITS #(.width(1), .high(0), .low(0)) bits_1551 (
        .y(_T_324),
        .in(_T_307)
    );
    wire [7:0] _T_327;
    MUX_UNSIGNED #(.width(8)) u_mux_1552 (
        .y(_T_327),
        .sel(_T_324),
        .a(8'hFF),
        .b(8'h0)
    );
    wire [7:0] _T_328;
    MUX_UNSIGNED #(.width(8)) u_mux_1553 (
        .y(_T_328),
        .sel(_T_304),
        .a(_T_323),
        .b(_T_327)
    );
    wire _T_329;
    BITWISEOR #(.width(1)) bitwiseor_1554 (
        .y(_T_329),
        .a(_T_304),
        .b(_T_309)
    );
    wire [22:0] _T_331;
    wire [22:0] _WTEMP_200;
    PAD_UNSIGNED #(.width(1), .n(23)) u_pad_1555 (
        .y(_WTEMP_200),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(23)) u_mux_1556 (
        .y(_T_331),
        .sel(_T_294),
        .a(_T_318),
        .b(_WTEMP_200)
    );
    wire [22:0] _T_332;
    MUX_UNSIGNED #(.width(23)) u_mux_1557 (
        .y(_T_332),
        .sel(_T_329),
        .a(_T_283),
        .b(_T_331)
    );
    wire [8:0] _T_333;
    CAT #(.width_a(1), .width_b(8)) cat_1558 (
        .y(_T_333),
        .a(_T_281),
        .b(_T_328)
    );
    wire [31:0] _T_334;
    CAT #(.width_a(9), .width_b(23)) cat_1559 (
        .y(_T_334),
        .a(_T_333),
        .b(_T_332)
    );
    wire _T_335;
    BITS #(.width(32), .high(31), .low(31)) bits_1560 (
        .y(_T_335),
        .in(_T_334)
    );
    wire _T_336;
    BITS #(.width(1), .high(0), .low(0)) bits_1561 (
        .y(_T_336),
        .in(_T_335)
    );
    wire [31:0] _T_339;
    MUX_UNSIGNED #(.width(32)) u_mux_1562 (
        .y(_T_339),
        .sel(_T_336),
        .a(32'hFFFFFFFF),
        .b(32'h0)
    );
    wire [63:0] unrec_s;
    CAT #(.width_a(32), .width_b(32)) cat_1563 (
        .y(unrec_s),
        .a(_T_339),
        .b(_T_334)
    );
    wire _T_340;
    BITS #(.width(65), .high(64), .low(64)) bits_1564 (
        .y(_T_340),
        .in(_in_in1__q)
    );
    wire [11:0] _T_341;
    BITS #(.width(65), .high(63), .low(52)) bits_1565 (
        .y(_T_341),
        .in(_in_in1__q)
    );
    wire [51:0] _T_342;
    BITS #(.width(65), .high(51), .low(0)) bits_1566 (
        .y(_T_342),
        .in(_in_in1__q)
    );
    wire [9:0] _T_343;
    BITS #(.width(12), .high(9), .low(0)) bits_1567 (
        .y(_T_343),
        .in(_T_341)
    );
    wire _T_345;
    wire [9:0] _WTEMP_201;
    PAD_UNSIGNED #(.width(2), .n(10)) u_pad_1568 (
        .y(_WTEMP_201),
        .in(2'h2)
    );
    LT_UNSIGNED #(.width(10)) u_lt_1569 (
        .y(_T_345),
        .a(_T_343),
        .b(_WTEMP_201)
    );
    wire [2:0] _T_346;
    BITS #(.width(12), .high(11), .low(9)) bits_1570 (
        .y(_T_346),
        .in(_T_341)
    );
    wire _T_348;
    wire [2:0] _WTEMP_202;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_1571 (
        .y(_WTEMP_202),
        .in(1'h1)
    );
    EQ_UNSIGNED #(.width(3)) u_eq_1572 (
        .y(_T_348),
        .a(_T_346),
        .b(_WTEMP_202)
    );
    wire [1:0] _T_349;
    BITS #(.width(12), .high(11), .low(10)) bits_1573 (
        .y(_T_349),
        .in(_T_341)
    );
    wire _T_351;
    wire [1:0] _WTEMP_203;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_1574 (
        .y(_WTEMP_203),
        .in(1'h1)
    );
    EQ_UNSIGNED #(.width(2)) u_eq_1575 (
        .y(_T_351),
        .a(_T_349),
        .b(_WTEMP_203)
    );
    wire _T_352;
    BITWISEAND #(.width(1)) bitwiseand_1576 (
        .y(_T_352),
        .a(_T_351),
        .b(_T_345)
    );
    wire _T_353;
    BITWISEOR #(.width(1)) bitwiseor_1577 (
        .y(_T_353),
        .a(_T_348),
        .b(_T_352)
    );
    wire [1:0] _T_354;
    BITS #(.width(12), .high(11), .low(10)) bits_1578 (
        .y(_T_354),
        .in(_T_341)
    );
    wire _T_356;
    wire [1:0] _WTEMP_204;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_1579 (
        .y(_WTEMP_204),
        .in(1'h1)
    );
    EQ_UNSIGNED #(.width(2)) u_eq_1580 (
        .y(_T_356),
        .a(_T_354),
        .b(_WTEMP_204)
    );
    wire _T_358;
    EQ_UNSIGNED #(.width(1)) u_eq_1581 (
        .y(_T_358),
        .a(_T_345),
        .b(1'h0)
    );
    wire _T_359;
    BITWISEAND #(.width(1)) bitwiseand_1582 (
        .y(_T_359),
        .a(_T_356),
        .b(_T_358)
    );
    wire [1:0] _T_360;
    BITS #(.width(12), .high(11), .low(10)) bits_1583 (
        .y(_T_360),
        .in(_T_341)
    );
    wire _T_362;
    EQ_UNSIGNED #(.width(2)) u_eq_1584 (
        .y(_T_362),
        .a(_T_360),
        .b(2'h2)
    );
    wire _T_363;
    BITWISEOR #(.width(1)) bitwiseor_1585 (
        .y(_T_363),
        .a(_T_359),
        .b(_T_362)
    );
    wire [1:0] _T_364;
    BITS #(.width(12), .high(11), .low(10)) bits_1586 (
        .y(_T_364),
        .in(_T_341)
    );
    wire _T_366;
    EQ_UNSIGNED #(.width(2)) u_eq_1587 (
        .y(_T_366),
        .a(_T_364),
        .b(2'h3)
    );
    wire _T_367;
    BITS #(.width(12), .high(9), .low(9)) bits_1588 (
        .y(_T_367),
        .in(_T_341)
    );
    wire _T_368;
    BITWISEAND #(.width(1)) bitwiseand_1589 (
        .y(_T_368),
        .a(_T_366),
        .b(_T_367)
    );
    wire [5:0] _T_370;
    BITS #(.width(12), .high(5), .low(0)) bits_1590 (
        .y(_T_370),
        .in(_T_341)
    );
    wire [6:0] _T_371;
    wire [5:0] _WTEMP_205;
    PAD_UNSIGNED #(.width(2), .n(6)) u_pad_1591 (
        .y(_WTEMP_205),
        .in(2'h2)
    );
    SUB_UNSIGNED #(.width(6)) u_sub_1592 (
        .y(_T_371),
        .a(_WTEMP_205),
        .b(_T_370)
    );
    wire [6:0] _T_372;
    ASUINT #(.width(7)) asuint_1593 (
        .y(_T_372),
        .in(_T_371)
    );
    wire [5:0] _T_373;
    TAIL #(.width(7), .n(1)) tail_1594 (
        .y(_T_373),
        .in(_T_372)
    );
    wire [52:0] _T_375;
    CAT #(.width_a(1), .width_b(52)) cat_1595 (
        .y(_T_375),
        .a(1'h1),
        .b(_T_342)
    );
    wire [52:0] _T_376;
    DSHR_UNSIGNED #(.width_in(53), .width_n(6)) u_dshr_1596 (
        .y(_T_376),
        .in(_T_375),
        .n(_T_373)
    );
    wire [51:0] _T_377;
    BITS #(.width(53), .high(51), .low(0)) bits_1597 (
        .y(_T_377),
        .in(_T_376)
    );
    wire [10:0] _T_378;
    BITS #(.width(12), .high(10), .low(0)) bits_1598 (
        .y(_T_378),
        .in(_T_341)
    );
    wire [11:0] _T_380;
    SUB_UNSIGNED #(.width(11)) u_sub_1599 (
        .y(_T_380),
        .a(_T_378),
        .b(11'h401)
    );
    wire [11:0] _T_381;
    ASUINT #(.width(12)) asuint_1600 (
        .y(_T_381),
        .in(_T_380)
    );
    wire [10:0] _T_382;
    TAIL #(.width(12), .n(1)) tail_1601 (
        .y(_T_382),
        .in(_T_381)
    );
    wire _T_383;
    BITS #(.width(1), .high(0), .low(0)) bits_1602 (
        .y(_T_383),
        .in(_T_366)
    );
    wire [10:0] _T_386;
    MUX_UNSIGNED #(.width(11)) u_mux_1603 (
        .y(_T_386),
        .sel(_T_383),
        .a(11'h7FF),
        .b(11'h0)
    );
    wire [10:0] _T_387;
    MUX_UNSIGNED #(.width(11)) u_mux_1604 (
        .y(_T_387),
        .sel(_T_363),
        .a(_T_382),
        .b(_T_386)
    );
    wire _T_388;
    BITWISEOR #(.width(1)) bitwiseor_1605 (
        .y(_T_388),
        .a(_T_363),
        .b(_T_368)
    );
    wire [51:0] _T_390;
    wire [51:0] _WTEMP_206;
    PAD_UNSIGNED #(.width(1), .n(52)) u_pad_1606 (
        .y(_WTEMP_206),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(52)) u_mux_1607 (
        .y(_T_390),
        .sel(_T_353),
        .a(_T_377),
        .b(_WTEMP_206)
    );
    wire [51:0] _T_391;
    MUX_UNSIGNED #(.width(52)) u_mux_1608 (
        .y(_T_391),
        .sel(_T_388),
        .a(_T_342),
        .b(_T_390)
    );
    wire [11:0] _T_392;
    CAT #(.width_a(1), .width_b(11)) cat_1609 (
        .y(_T_392),
        .a(_T_340),
        .b(_T_387)
    );
    wire [63:0] _T_393;
    CAT #(.width_a(12), .width_b(52)) cat_1610 (
        .y(_T_393),
        .a(_T_392),
        .b(_T_391)
    );
    wire [63:0] unrec_int;
    MUX_UNSIGNED #(.width(64)) u_mux_1611 (
        .y(unrec_int),
        .sel(_in_single__q),
        .a(unrec_s),
        .b(_T_393)
    );
    wire _T_394;
    BITS #(.width(65), .high(32), .low(32)) bits_1612 (
        .y(_T_394),
        .in(_in_in1__q)
    );
    wire [8:0] _T_395;
    BITS #(.width(65), .high(31), .low(23)) bits_1613 (
        .y(_T_395),
        .in(_in_in1__q)
    );
    wire [22:0] _T_396;
    BITS #(.width(65), .high(22), .low(0)) bits_1614 (
        .y(_T_396),
        .in(_in_in1__q)
    );
    wire [2:0] _T_397;
    BITS #(.width(9), .high(8), .low(6)) bits_1615 (
        .y(_T_397),
        .in(_T_395)
    );
    wire [1:0] _T_398;
    BITS #(.width(3), .high(2), .low(1)) bits_1616 (
        .y(_T_398),
        .in(_T_397)
    );
    wire _T_400;
    EQ_UNSIGNED #(.width(2)) u_eq_1617 (
        .y(_T_400),
        .a(_T_398),
        .b(2'h3)
    );
    wire [6:0] _T_401;
    BITS #(.width(9), .high(6), .low(0)) bits_1618 (
        .y(_T_401),
        .in(_T_395)
    );
    wire _T_403;
    wire [6:0] _WTEMP_207;
    PAD_UNSIGNED #(.width(2), .n(7)) u_pad_1619 (
        .y(_WTEMP_207),
        .in(2'h2)
    );
    LT_UNSIGNED #(.width(7)) u_lt_1620 (
        .y(_T_403),
        .a(_T_401),
        .b(_WTEMP_207)
    );
    wire _T_405;
    wire [2:0] _WTEMP_208;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_1621 (
        .y(_WTEMP_208),
        .in(1'h1)
    );
    EQ_UNSIGNED #(.width(3)) u_eq_1622 (
        .y(_T_405),
        .a(_T_397),
        .b(_WTEMP_208)
    );
    wire _T_407;
    wire [1:0] _WTEMP_209;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_1623 (
        .y(_WTEMP_209),
        .in(1'h1)
    );
    EQ_UNSIGNED #(.width(2)) u_eq_1624 (
        .y(_T_407),
        .a(_T_398),
        .b(_WTEMP_209)
    );
    wire _T_408;
    BITWISEAND #(.width(1)) bitwiseand_1625 (
        .y(_T_408),
        .a(_T_407),
        .b(_T_403)
    );
    wire _T_409;
    BITWISEOR #(.width(1)) bitwiseor_1626 (
        .y(_T_409),
        .a(_T_405),
        .b(_T_408)
    );
    wire _T_411;
    wire [1:0] _WTEMP_210;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_1627 (
        .y(_WTEMP_210),
        .in(1'h1)
    );
    EQ_UNSIGNED #(.width(2)) u_eq_1628 (
        .y(_T_411),
        .a(_T_398),
        .b(_WTEMP_210)
    );
    wire _T_413;
    EQ_UNSIGNED #(.width(1)) u_eq_1629 (
        .y(_T_413),
        .a(_T_403),
        .b(1'h0)
    );
    wire _T_414;
    BITWISEAND #(.width(1)) bitwiseand_1630 (
        .y(_T_414),
        .a(_T_411),
        .b(_T_413)
    );
    wire _T_416;
    EQ_UNSIGNED #(.width(2)) u_eq_1631 (
        .y(_T_416),
        .a(_T_398),
        .b(2'h2)
    );
    wire _T_417;
    BITWISEOR #(.width(1)) bitwiseor_1632 (
        .y(_T_417),
        .a(_T_414),
        .b(_T_416)
    );
    wire _T_419;
    wire [2:0] _WTEMP_211;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_1633 (
        .y(_WTEMP_211),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(3)) u_eq_1634 (
        .y(_T_419),
        .a(_T_397),
        .b(_WTEMP_211)
    );
    wire _T_420;
    BITS #(.width(9), .high(6), .low(6)) bits_1635 (
        .y(_T_420),
        .in(_T_395)
    );
    wire _T_422;
    EQ_UNSIGNED #(.width(1)) u_eq_1636 (
        .y(_T_422),
        .a(_T_420),
        .b(1'h0)
    );
    wire _T_423;
    BITWISEAND #(.width(1)) bitwiseand_1637 (
        .y(_T_423),
        .a(_T_400),
        .b(_T_422)
    );
    wire [2:0] _T_424;
    BITWISENOT #(.width(3)) bitwisenot_1638 (
        .y(_T_424),
        .in(_T_397)
    );
    wire _T_426;
    wire [2:0] _WTEMP_212;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_1639 (
        .y(_WTEMP_212),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(3)) u_eq_1640 (
        .y(_T_426),
        .a(_T_424),
        .b(_WTEMP_212)
    );
    wire _T_427;
    BITS #(.width(23), .high(22), .low(22)) bits_1641 (
        .y(_T_427),
        .in(_T_396)
    );
    wire _T_429;
    EQ_UNSIGNED #(.width(1)) u_eq_1642 (
        .y(_T_429),
        .a(_T_427),
        .b(1'h0)
    );
    wire _T_430;
    BITWISEAND #(.width(1)) bitwiseand_1643 (
        .y(_T_430),
        .a(_T_426),
        .b(_T_429)
    );
    wire _T_431;
    BITS #(.width(23), .high(22), .low(22)) bits_1644 (
        .y(_T_431),
        .in(_T_396)
    );
    wire _T_432;
    BITWISEAND #(.width(1)) bitwiseand_1645 (
        .y(_T_432),
        .a(_T_426),
        .b(_T_431)
    );
    wire _T_434;
    EQ_UNSIGNED #(.width(1)) u_eq_1646 (
        .y(_T_434),
        .a(_T_394),
        .b(1'h0)
    );
    wire _T_435;
    BITWISEAND #(.width(1)) bitwiseand_1647 (
        .y(_T_435),
        .a(_T_423),
        .b(_T_434)
    );
    wire _T_437;
    EQ_UNSIGNED #(.width(1)) u_eq_1648 (
        .y(_T_437),
        .a(_T_394),
        .b(1'h0)
    );
    wire _T_438;
    BITWISEAND #(.width(1)) bitwiseand_1649 (
        .y(_T_438),
        .a(_T_417),
        .b(_T_437)
    );
    wire _T_440;
    EQ_UNSIGNED #(.width(1)) u_eq_1650 (
        .y(_T_440),
        .a(_T_394),
        .b(1'h0)
    );
    wire _T_441;
    BITWISEAND #(.width(1)) bitwiseand_1651 (
        .y(_T_441),
        .a(_T_409),
        .b(_T_440)
    );
    wire _T_443;
    EQ_UNSIGNED #(.width(1)) u_eq_1652 (
        .y(_T_443),
        .a(_T_394),
        .b(1'h0)
    );
    wire _T_444;
    BITWISEAND #(.width(1)) bitwiseand_1653 (
        .y(_T_444),
        .a(_T_419),
        .b(_T_443)
    );
    wire _T_445;
    BITWISEAND #(.width(1)) bitwiseand_1654 (
        .y(_T_445),
        .a(_T_419),
        .b(_T_394)
    );
    wire _T_446;
    BITWISEAND #(.width(1)) bitwiseand_1655 (
        .y(_T_446),
        .a(_T_409),
        .b(_T_394)
    );
    wire _T_447;
    BITWISEAND #(.width(1)) bitwiseand_1656 (
        .y(_T_447),
        .a(_T_417),
        .b(_T_394)
    );
    wire _T_448;
    BITWISEAND #(.width(1)) bitwiseand_1657 (
        .y(_T_448),
        .a(_T_423),
        .b(_T_394)
    );
    wire [1:0] _T_449;
    CAT #(.width_a(1), .width_b(1)) cat_1658 (
        .y(_T_449),
        .a(_T_447),
        .b(_T_448)
    );
    wire [1:0] _T_450;
    CAT #(.width_a(1), .width_b(1)) cat_1659 (
        .y(_T_450),
        .a(_T_444),
        .b(_T_445)
    );
    wire [2:0] _T_451;
    CAT #(.width_a(2), .width_b(1)) cat_1660 (
        .y(_T_451),
        .a(_T_450),
        .b(_T_446)
    );
    wire [4:0] _T_452;
    CAT #(.width_a(3), .width_b(2)) cat_1661 (
        .y(_T_452),
        .a(_T_451),
        .b(_T_449)
    );
    wire [1:0] _T_453;
    CAT #(.width_a(1), .width_b(1)) cat_1662 (
        .y(_T_453),
        .a(_T_438),
        .b(_T_441)
    );
    wire [1:0] _T_454;
    CAT #(.width_a(1), .width_b(1)) cat_1663 (
        .y(_T_454),
        .a(_T_432),
        .b(_T_430)
    );
    wire [2:0] _T_455;
    CAT #(.width_a(2), .width_b(1)) cat_1664 (
        .y(_T_455),
        .a(_T_454),
        .b(_T_435)
    );
    wire [4:0] _T_456;
    CAT #(.width_a(3), .width_b(2)) cat_1665 (
        .y(_T_456),
        .a(_T_455),
        .b(_T_453)
    );
    wire [9:0] classify_s;
    CAT #(.width_a(5), .width_b(5)) cat_1666 (
        .y(classify_s),
        .a(_T_456),
        .b(_T_452)
    );
    wire _T_457;
    BITS #(.width(65), .high(64), .low(64)) bits_1667 (
        .y(_T_457),
        .in(_in_in1__q)
    );
    wire [11:0] _T_458;
    BITS #(.width(65), .high(63), .low(52)) bits_1668 (
        .y(_T_458),
        .in(_in_in1__q)
    );
    wire [51:0] _T_459;
    BITS #(.width(65), .high(51), .low(0)) bits_1669 (
        .y(_T_459),
        .in(_in_in1__q)
    );
    wire [2:0] _T_460;
    BITS #(.width(12), .high(11), .low(9)) bits_1670 (
        .y(_T_460),
        .in(_T_458)
    );
    wire [1:0] _T_461;
    BITS #(.width(3), .high(2), .low(1)) bits_1671 (
        .y(_T_461),
        .in(_T_460)
    );
    wire _T_463;
    EQ_UNSIGNED #(.width(2)) u_eq_1672 (
        .y(_T_463),
        .a(_T_461),
        .b(2'h3)
    );
    wire [9:0] _T_464;
    BITS #(.width(12), .high(9), .low(0)) bits_1673 (
        .y(_T_464),
        .in(_T_458)
    );
    wire _T_466;
    wire [9:0] _WTEMP_213;
    PAD_UNSIGNED #(.width(2), .n(10)) u_pad_1674 (
        .y(_WTEMP_213),
        .in(2'h2)
    );
    LT_UNSIGNED #(.width(10)) u_lt_1675 (
        .y(_T_466),
        .a(_T_464),
        .b(_WTEMP_213)
    );
    wire _T_468;
    wire [2:0] _WTEMP_214;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_1676 (
        .y(_WTEMP_214),
        .in(1'h1)
    );
    EQ_UNSIGNED #(.width(3)) u_eq_1677 (
        .y(_T_468),
        .a(_T_460),
        .b(_WTEMP_214)
    );
    wire _T_470;
    wire [1:0] _WTEMP_215;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_1678 (
        .y(_WTEMP_215),
        .in(1'h1)
    );
    EQ_UNSIGNED #(.width(2)) u_eq_1679 (
        .y(_T_470),
        .a(_T_461),
        .b(_WTEMP_215)
    );
    wire _T_471;
    BITWISEAND #(.width(1)) bitwiseand_1680 (
        .y(_T_471),
        .a(_T_470),
        .b(_T_466)
    );
    wire _T_472;
    BITWISEOR #(.width(1)) bitwiseor_1681 (
        .y(_T_472),
        .a(_T_468),
        .b(_T_471)
    );
    wire _T_474;
    wire [1:0] _WTEMP_216;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_1682 (
        .y(_WTEMP_216),
        .in(1'h1)
    );
    EQ_UNSIGNED #(.width(2)) u_eq_1683 (
        .y(_T_474),
        .a(_T_461),
        .b(_WTEMP_216)
    );
    wire _T_476;
    EQ_UNSIGNED #(.width(1)) u_eq_1684 (
        .y(_T_476),
        .a(_T_466),
        .b(1'h0)
    );
    wire _T_477;
    BITWISEAND #(.width(1)) bitwiseand_1685 (
        .y(_T_477),
        .a(_T_474),
        .b(_T_476)
    );
    wire _T_479;
    EQ_UNSIGNED #(.width(2)) u_eq_1686 (
        .y(_T_479),
        .a(_T_461),
        .b(2'h2)
    );
    wire _T_480;
    BITWISEOR #(.width(1)) bitwiseor_1687 (
        .y(_T_480),
        .a(_T_477),
        .b(_T_479)
    );
    wire _T_482;
    wire [2:0] _WTEMP_217;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_1688 (
        .y(_WTEMP_217),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(3)) u_eq_1689 (
        .y(_T_482),
        .a(_T_460),
        .b(_WTEMP_217)
    );
    wire _T_483;
    BITS #(.width(12), .high(9), .low(9)) bits_1690 (
        .y(_T_483),
        .in(_T_458)
    );
    wire _T_485;
    EQ_UNSIGNED #(.width(1)) u_eq_1691 (
        .y(_T_485),
        .a(_T_483),
        .b(1'h0)
    );
    wire _T_486;
    BITWISEAND #(.width(1)) bitwiseand_1692 (
        .y(_T_486),
        .a(_T_463),
        .b(_T_485)
    );
    wire [2:0] _T_487;
    BITWISENOT #(.width(3)) bitwisenot_1693 (
        .y(_T_487),
        .in(_T_460)
    );
    wire _T_489;
    wire [2:0] _WTEMP_218;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_1694 (
        .y(_WTEMP_218),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(3)) u_eq_1695 (
        .y(_T_489),
        .a(_T_487),
        .b(_WTEMP_218)
    );
    wire _T_490;
    BITS #(.width(52), .high(51), .low(51)) bits_1696 (
        .y(_T_490),
        .in(_T_459)
    );
    wire _T_492;
    EQ_UNSIGNED #(.width(1)) u_eq_1697 (
        .y(_T_492),
        .a(_T_490),
        .b(1'h0)
    );
    wire _T_493;
    BITWISEAND #(.width(1)) bitwiseand_1698 (
        .y(_T_493),
        .a(_T_489),
        .b(_T_492)
    );
    wire _T_494;
    BITS #(.width(52), .high(51), .low(51)) bits_1699 (
        .y(_T_494),
        .in(_T_459)
    );
    wire _T_495;
    BITWISEAND #(.width(1)) bitwiseand_1700 (
        .y(_T_495),
        .a(_T_489),
        .b(_T_494)
    );
    wire _T_497;
    EQ_UNSIGNED #(.width(1)) u_eq_1701 (
        .y(_T_497),
        .a(_T_457),
        .b(1'h0)
    );
    wire _T_498;
    BITWISEAND #(.width(1)) bitwiseand_1702 (
        .y(_T_498),
        .a(_T_486),
        .b(_T_497)
    );
    wire _T_500;
    EQ_UNSIGNED #(.width(1)) u_eq_1703 (
        .y(_T_500),
        .a(_T_457),
        .b(1'h0)
    );
    wire _T_501;
    BITWISEAND #(.width(1)) bitwiseand_1704 (
        .y(_T_501),
        .a(_T_480),
        .b(_T_500)
    );
    wire _T_503;
    EQ_UNSIGNED #(.width(1)) u_eq_1705 (
        .y(_T_503),
        .a(_T_457),
        .b(1'h0)
    );
    wire _T_504;
    BITWISEAND #(.width(1)) bitwiseand_1706 (
        .y(_T_504),
        .a(_T_472),
        .b(_T_503)
    );
    wire _T_506;
    EQ_UNSIGNED #(.width(1)) u_eq_1707 (
        .y(_T_506),
        .a(_T_457),
        .b(1'h0)
    );
    wire _T_507;
    BITWISEAND #(.width(1)) bitwiseand_1708 (
        .y(_T_507),
        .a(_T_482),
        .b(_T_506)
    );
    wire _T_508;
    BITWISEAND #(.width(1)) bitwiseand_1709 (
        .y(_T_508),
        .a(_T_482),
        .b(_T_457)
    );
    wire _T_509;
    BITWISEAND #(.width(1)) bitwiseand_1710 (
        .y(_T_509),
        .a(_T_472),
        .b(_T_457)
    );
    wire _T_510;
    BITWISEAND #(.width(1)) bitwiseand_1711 (
        .y(_T_510),
        .a(_T_480),
        .b(_T_457)
    );
    wire _T_511;
    BITWISEAND #(.width(1)) bitwiseand_1712 (
        .y(_T_511),
        .a(_T_486),
        .b(_T_457)
    );
    wire [1:0] _T_512;
    CAT #(.width_a(1), .width_b(1)) cat_1713 (
        .y(_T_512),
        .a(_T_510),
        .b(_T_511)
    );
    wire [1:0] _T_513;
    CAT #(.width_a(1), .width_b(1)) cat_1714 (
        .y(_T_513),
        .a(_T_507),
        .b(_T_508)
    );
    wire [2:0] _T_514;
    CAT #(.width_a(2), .width_b(1)) cat_1715 (
        .y(_T_514),
        .a(_T_513),
        .b(_T_509)
    );
    wire [4:0] _T_515;
    CAT #(.width_a(3), .width_b(2)) cat_1716 (
        .y(_T_515),
        .a(_T_514),
        .b(_T_512)
    );
    wire [1:0] _T_516;
    CAT #(.width_a(1), .width_b(1)) cat_1717 (
        .y(_T_516),
        .a(_T_501),
        .b(_T_504)
    );
    wire [1:0] _T_517;
    CAT #(.width_a(1), .width_b(1)) cat_1718 (
        .y(_T_517),
        .a(_T_495),
        .b(_T_493)
    );
    wire [2:0] _T_518;
    CAT #(.width_a(2), .width_b(1)) cat_1719 (
        .y(_T_518),
        .a(_T_517),
        .b(_T_498)
    );
    wire [4:0] _T_519;
    CAT #(.width_a(3), .width_b(2)) cat_1720 (
        .y(_T_519),
        .a(_T_518),
        .b(_T_516)
    );
    wire [9:0] _T_520;
    CAT #(.width_a(5), .width_b(5)) cat_1721 (
        .y(_T_520),
        .a(_T_519),
        .b(_T_515)
    );
    wire [9:0] classify_out;
    MUX_UNSIGNED #(.width(10)) u_mux_1722 (
        .y(classify_out),
        .sel(_in_single__q),
        .a(classify_s),
        .b(_T_520)
    );
    wire _dcmp__clock;
    wire _dcmp__reset;
    wire [64:0] _dcmp__io_a;
    wire [64:0] _dcmp__io_b;
    wire _dcmp__io_signaling;
    wire _dcmp__io_lt;
    wire _dcmp__io_eq;
    wire _dcmp__io_gt;
    wire [4:0] _dcmp__io_exceptionFlags;
    CompareRecFN dcmp (
        .clock(_dcmp__clock),
        .reset(_dcmp__reset),
        .io_a(_dcmp__io_a),
        .io_b(_dcmp__io_b),
        .io_signaling(_dcmp__io_signaling),
        .io_lt(_dcmp__io_lt),
        .io_eq(_dcmp__io_eq),
        .io_gt(_dcmp__io_gt),
        .io_exceptionFlags(_dcmp__io_exceptionFlags)
    );
    wire _T_521;
    BITS #(.width(3), .high(1), .low(1)) bits_1806 (
        .y(_T_521),
        .in(_in_rm__q)
    );
    wire _T_523;
    EQ_UNSIGNED #(.width(1)) u_eq_1807 (
        .y(_T_523),
        .a(_T_521),
        .b(1'h0)
    );
    wire _T_524;
    BITS #(.width(3), .high(0), .low(0)) bits_1808 (
        .y(_T_524),
        .in(_in_rm__q)
    );
    wire [63:0] _T_525;
    wire [63:0] _WTEMP_221;
    PAD_UNSIGNED #(.width(10), .n(64)) u_pad_1809 (
        .y(_WTEMP_221),
        .in(classify_out)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_1810 (
        .y(_T_525),
        .sel(_T_524),
        .a(_WTEMP_221),
        .b(unrec_int)
    );
    wire [4:0] _T_529;
    wire [4:0] _WTEMP_222;
    PAD_UNSIGNED #(.width(4), .n(5)) u_pad_1811 (
        .y(_WTEMP_222),
        .in(4'hC)
    );
    BITWISEAND #(.width(5)) bitwiseand_1812 (
        .y(_T_529),
        .a(_in_cmd__q),
        .b(_WTEMP_222)
    );
    wire _T_530;
    wire [4:0] _WTEMP_223;
    PAD_UNSIGNED #(.width(3), .n(5)) u_pad_1813 (
        .y(_WTEMP_223),
        .in(3'h4)
    );
    EQ_UNSIGNED #(.width(5)) u_eq_1814 (
        .y(_T_530),
        .a(_WTEMP_223),
        .b(_T_529)
    );
    wire [2:0] _T_531;
    BITWISENOT #(.width(3)) bitwisenot_1815 (
        .y(_T_531),
        .in(_in_rm__q)
    );
    wire [1:0] _T_532;
    CAT #(.width_a(1), .width_b(1)) cat_1816 (
        .y(_T_532),
        .a(_dcmp__io_lt),
        .b(_dcmp__io_eq)
    );
    wire [2:0] _T_533;
    wire [2:0] _WTEMP_224;
    PAD_UNSIGNED #(.width(2), .n(3)) u_pad_1817 (
        .y(_WTEMP_224),
        .in(_T_532)
    );
    BITWISEAND #(.width(3)) bitwiseand_1818 (
        .y(_T_533),
        .a(_T_531),
        .b(_WTEMP_224)
    );
    wire _T_535;
    wire [2:0] _WTEMP_225;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_1819 (
        .y(_WTEMP_225),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(3)) u_neq_1820 (
        .y(_T_535),
        .a(_T_533),
        .b(_WTEMP_225)
    );
    wire [4:0] _T_538;
    wire [4:0] _WTEMP_226;
    PAD_UNSIGNED #(.width(4), .n(5)) u_pad_1821 (
        .y(_WTEMP_226),
        .in(4'hC)
    );
    BITWISEAND #(.width(5)) bitwiseand_1822 (
        .y(_T_538),
        .a(_in_cmd__q),
        .b(_WTEMP_226)
    );
    wire _T_539;
    wire [4:0] _WTEMP_227;
    PAD_UNSIGNED #(.width(4), .n(5)) u_pad_1823 (
        .y(_WTEMP_227),
        .in(4'h8)
    );
    EQ_UNSIGNED #(.width(5)) u_eq_1824 (
        .y(_T_539),
        .a(_WTEMP_227),
        .b(_T_538)
    );
    wire _RecFNToIN__clock;
    wire _RecFNToIN__reset;
    wire [64:0] _RecFNToIN__io_in;
    wire [1:0] _RecFNToIN__io_roundingMode;
    wire _RecFNToIN__io_signedOut;
    wire [31:0] _RecFNToIN__io_out;
    wire [2:0] _RecFNToIN__io_intExceptionFlags;
    RecFNToIN RecFNToIN (
        .clock(_RecFNToIN__clock),
        .reset(_RecFNToIN__reset),
        .io_in(_RecFNToIN__io_in),
        .io_roundingMode(_RecFNToIN__io_roundingMode),
        .io_signedOut(_RecFNToIN__io_signedOut),
        .io_out(_RecFNToIN__io_out),
        .io_intExceptionFlags(_RecFNToIN__io_intExceptionFlags)
    );
    wire _T_540;
    BITS #(.width(2), .high(0), .low(0)) bits_1950 (
        .y(_T_540),
        .in(_in_typ__q)
    );
    wire _T_541;
    BITWISENOT #(.width(1)) bitwisenot_1951 (
        .y(_T_541),
        .in(_T_540)
    );
    wire _T_542;
    BITS #(.width(2), .high(1), .low(1)) bits_1952 (
        .y(_T_542),
        .in(_in_typ__q)
    );
    wire _T_544;
    EQ_UNSIGNED #(.width(1)) u_eq_1953 (
        .y(_T_544),
        .a(_T_542),
        .b(1'h0)
    );
    wire _T_545;
    BITS #(.width(32), .high(31), .low(31)) bits_1954 (
        .y(_T_545),
        .in(_RecFNToIN__io_out)
    );
    wire _T_546;
    BITS #(.width(1), .high(0), .low(0)) bits_1955 (
        .y(_T_546),
        .in(_T_545)
    );
    wire [31:0] _T_549;
    MUX_UNSIGNED #(.width(32)) u_mux_1956 (
        .y(_T_549),
        .sel(_T_546),
        .a(32'hFFFFFFFF),
        .b(32'h0)
    );
    wire [63:0] _T_550;
    CAT #(.width_a(32), .width_b(32)) cat_1957 (
        .y(_T_550),
        .a(_T_549),
        .b(_RecFNToIN__io_out)
    );
    wire [1:0] _T_551;
    BITS #(.width(3), .high(2), .low(1)) bits_1958 (
        .y(_T_551),
        .in(_RecFNToIN__io_intExceptionFlags)
    );
    wire _T_553;
    wire [1:0] _WTEMP_248;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_1959 (
        .y(_WTEMP_248),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(2)) u_neq_1960 (
        .y(_T_553),
        .a(_T_551),
        .b(_WTEMP_248)
    );
    wire _T_555;
    BITS #(.width(3), .high(0), .low(0)) bits_1961 (
        .y(_T_555),
        .in(_RecFNToIN__io_intExceptionFlags)
    );
    wire [3:0] _T_556;
    CAT #(.width_a(1), .width_b(3)) cat_1962 (
        .y(_T_556),
        .a(_T_553),
        .b(3'h0)
    );
    wire [4:0] _T_557;
    CAT #(.width_a(4), .width_b(1)) cat_1963 (
        .y(_T_557),
        .a(_T_556),
        .b(_T_555)
    );
    wire [4:0] _node_19;
    wire [4:0] _WTEMP_249;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_1964 (
        .y(_WTEMP_249),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(5)) u_mux_1965 (
        .y(_node_19),
        .sel(_T_530),
        .a(_dcmp__io_exceptionFlags),
        .b(_WTEMP_249)
    );
    wire [63:0] _node_20;
    wire [63:0] _WTEMP_250;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_1966 (
        .y(_WTEMP_250),
        .in(_T_535)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_1967 (
        .y(_node_20),
        .sel(_T_530),
        .a(_WTEMP_250),
        .b(_T_525)
    );
    wire _RecFNToIN_1__clock;
    wire _RecFNToIN_1__reset;
    wire [64:0] _RecFNToIN_1__io_in;
    wire [1:0] _RecFNToIN_1__io_roundingMode;
    wire _RecFNToIN_1__io_signedOut;
    wire [63:0] _RecFNToIN_1__io_out;
    wire [2:0] _RecFNToIN_1__io_intExceptionFlags;
    RecFNToIN_1 RecFNToIN_1 (
        .clock(_RecFNToIN_1__clock),
        .reset(_RecFNToIN_1__reset),
        .io_in(_RecFNToIN_1__io_in),
        .io_roundingMode(_RecFNToIN_1__io_roundingMode),
        .io_signedOut(_RecFNToIN_1__io_signedOut),
        .io_out(_RecFNToIN_1__io_out),
        .io_intExceptionFlags(_RecFNToIN_1__io_intExceptionFlags)
    );
    wire _T_558;
    BITS #(.width(2), .high(0), .low(0)) bits_2093 (
        .y(_T_558),
        .in(_in_typ__q)
    );
    wire _T_559;
    BITWISENOT #(.width(1)) bitwisenot_2094 (
        .y(_T_559),
        .in(_T_558)
    );
    wire _T_560;
    BITS #(.width(2), .high(1), .low(1)) bits_2095 (
        .y(_T_560),
        .in(_in_typ__q)
    );
    wire _T_562;
    EQ_UNSIGNED #(.width(1)) u_eq_2096 (
        .y(_T_562),
        .a(_T_560),
        .b(1'h1)
    );
    wire [1:0] _T_563;
    BITS #(.width(3), .high(2), .low(1)) bits_2097 (
        .y(_T_563),
        .in(_RecFNToIN_1__io_intExceptionFlags)
    );
    wire _T_565;
    wire [1:0] _WTEMP_271;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2098 (
        .y(_WTEMP_271),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(2)) u_neq_2099 (
        .y(_T_565),
        .a(_T_563),
        .b(_WTEMP_271)
    );
    wire _T_567;
    BITS #(.width(3), .high(0), .low(0)) bits_2100 (
        .y(_T_567),
        .in(_RecFNToIN_1__io_intExceptionFlags)
    );
    wire [3:0] _T_568;
    CAT #(.width_a(1), .width_b(3)) cat_2101 (
        .y(_T_568),
        .a(_T_565),
        .b(3'h0)
    );
    wire [4:0] _T_569;
    CAT #(.width_a(4), .width_b(1)) cat_2102 (
        .y(_T_569),
        .a(_T_568),
        .b(_T_567)
    );
    wire [4:0] _node_21;
    MUX_UNSIGNED #(.width(5)) u_mux_2103 (
        .y(_node_21),
        .sel(_T_544),
        .a(_T_557),
        .b(_node_19)
    );
    wire [63:0] _node_22;
    MUX_UNSIGNED #(.width(64)) u_mux_2104 (
        .y(_node_22),
        .sel(_T_544),
        .a(_T_550),
        .b(_node_20)
    );
    wire [4:0] _node_23;
    MUX_UNSIGNED #(.width(5)) u_mux_2105 (
        .y(_node_23),
        .sel(_T_562),
        .a(_T_569),
        .b(_node_21)
    );
    wire [4:0] _node_24;
    wire [4:0] _WTEMP_272;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_2106 (
        .y(_WTEMP_272),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(5)) u_mux_2107 (
        .y(_node_24),
        .sel(_T_530),
        .a(_dcmp__io_exceptionFlags),
        .b(_WTEMP_272)
    );
    wire [63:0] _node_25;
    MUX_UNSIGNED #(.width(64)) u_mux_2108 (
        .y(_node_25),
        .sel(_T_562),
        .a(_RecFNToIN_1__io_out),
        .b(_node_22)
    );
    wire [63:0] _node_26;
    wire [63:0] _WTEMP_273;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_2109 (
        .y(_WTEMP_273),
        .in(_T_535)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_2110 (
        .y(_node_26),
        .sel(_T_530),
        .a(_WTEMP_273),
        .b(_T_525)
    );
    assign _RecFNToIN__clock = clock;
    assign _RecFNToIN__io_in = _in_in1__q;
    BITS #(.width(3), .high(1), .low(0)) bits_2111 (
        .y(_RecFNToIN__io_roundingMode),
        .in(_in_rm__q)
    );
    assign _RecFNToIN__io_signedOut = _T_541;
    assign _RecFNToIN__reset = reset;
    assign _RecFNToIN_1__clock = clock;
    assign _RecFNToIN_1__io_in = _in_in1__q;
    BITS #(.width(3), .high(1), .low(0)) bits_2112 (
        .y(_RecFNToIN_1__io_roundingMode),
        .in(_in_rm__q)
    );
    assign _RecFNToIN_1__io_signedOut = _T_559;
    assign _RecFNToIN_1__reset = reset;
    assign _dcmp__clock = clock;
    assign _dcmp__io_a = _in_in1__q;
    assign _dcmp__io_b = _in_in2__q;
    assign _dcmp__io_signaling = _T_523;
    assign _dcmp__reset = reset;
    MUX_UNSIGNED #(.width(5)) u_mux_2113 (
        .y(_in_cmd__d),
        .sel(io_in_valid),
        .a(io_in_bits_cmd),
        .b(_in_cmd__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_2114 (
        .y(_in_div__d),
        .sel(io_in_valid),
        .a(io_in_bits_div),
        .b(_in_div__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_2115 (
        .y(_in_fastpipe__d),
        .sel(io_in_valid),
        .a(io_in_bits_fastpipe),
        .b(_in_fastpipe__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_2116 (
        .y(_in_fma__d),
        .sel(io_in_valid),
        .a(io_in_bits_fma),
        .b(_in_fma__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_2117 (
        .y(_in_fromint__d),
        .sel(io_in_valid),
        .a(io_in_bits_fromint),
        .b(_in_fromint__q)
    );
    MUX_UNSIGNED #(.width(65)) u_mux_2118 (
        .y(_in_in1__d),
        .sel(io_in_valid),
        .a(_node_17),
        .b(_in_in1__q)
    );
    MUX_UNSIGNED #(.width(65)) u_mux_2119 (
        .y(_in_in2__d),
        .sel(io_in_valid),
        .a(_node_18),
        .b(_in_in2__q)
    );
    MUX_UNSIGNED #(.width(65)) u_mux_2120 (
        .y(_in_in3__d),
        .sel(io_in_valid),
        .a(io_in_bits_in3),
        .b(_in_in3__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_2121 (
        .y(_in_ldst__d),
        .sel(io_in_valid),
        .a(io_in_bits_ldst),
        .b(_in_ldst__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_2122 (
        .y(_in_ren1__d),
        .sel(io_in_valid),
        .a(io_in_bits_ren1),
        .b(_in_ren1__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_2123 (
        .y(_in_ren2__d),
        .sel(io_in_valid),
        .a(io_in_bits_ren2),
        .b(_in_ren2__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_2124 (
        .y(_in_ren3__d),
        .sel(io_in_valid),
        .a(io_in_bits_ren3),
        .b(_in_ren3__q)
    );
    MUX_UNSIGNED #(.width(3)) u_mux_2125 (
        .y(_in_rm__d),
        .sel(io_in_valid),
        .a(io_in_bits_rm),
        .b(_in_rm__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_2126 (
        .y(_in_single__d),
        .sel(io_in_valid),
        .a(io_in_bits_single),
        .b(_in_single__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_2127 (
        .y(_in_sqrt__d),
        .sel(io_in_valid),
        .a(io_in_bits_sqrt),
        .b(_in_sqrt__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_2128 (
        .y(_in_swap12__d),
        .sel(io_in_valid),
        .a(io_in_bits_swap12),
        .b(_in_swap12__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_2129 (
        .y(_in_swap23__d),
        .sel(io_in_valid),
        .a(io_in_bits_swap23),
        .b(_in_swap23__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_2130 (
        .y(_in_toint__d),
        .sel(io_in_valid),
        .a(io_in_bits_toint),
        .b(_in_toint__q)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_2131 (
        .y(_in_typ__d),
        .sel(io_in_valid),
        .a(io_in_bits_typ),
        .b(_in_typ__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_2132 (
        .y(_in_wen__d),
        .sel(io_in_valid),
        .a(io_in_bits_wen),
        .b(_in_wen__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_2133 (
        .y(_in_wflags__d),
        .sel(io_in_valid),
        .a(io_in_bits_wflags),
        .b(_in_wflags__q)
    );
    assign io_as_double_cmd = _in_cmd__q;
    assign io_as_double_div = _in_div__q;
    assign io_as_double_fastpipe = _in_fastpipe__q;
    assign io_as_double_fma = _in_fma__q;
    assign io_as_double_fromint = _in_fromint__q;
    assign io_as_double_in1 = _in_in1__q;
    assign io_as_double_in2 = _in_in2__q;
    assign io_as_double_in3 = _in_in3__q;
    assign io_as_double_ldst = _in_ldst__q;
    assign io_as_double_ren1 = _in_ren1__q;
    assign io_as_double_ren2 = _in_ren2__q;
    assign io_as_double_ren3 = _in_ren3__q;
    assign io_as_double_rm = _in_rm__q;
    assign io_as_double_single = _in_single__q;
    assign io_as_double_sqrt = _in_sqrt__q;
    assign io_as_double_swap12 = _in_swap12__q;
    assign io_as_double_swap23 = _in_swap23__q;
    assign io_as_double_toint = _in_toint__q;
    assign io_as_double_typ = _in_typ__q;
    assign io_as_double_wen = _in_wen__q;
    assign io_as_double_wflags = _in_wflags__q;
    MUX_UNSIGNED #(.width(5)) u_mux_2134 (
        .y(io_out_bits_exc),
        .sel(_T_539),
        .a(_node_23),
        .b(_node_24)
    );
    assign io_out_bits_lt = _dcmp__io_lt;
    assign io_out_bits_store = unrec_int;
    MUX_UNSIGNED #(.width(64)) u_mux_2135 (
        .y(io_out_bits_toint),
        .sel(_T_539),
        .a(_node_25),
        .b(_node_26)
    );
    assign io_out_valid = _valid__q;
    assign _valid__d = io_in_valid;
endmodule //FPToInt
module GEQ_UNSIGNED(y, a, b);
    parameter width = 4;
    output y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a >= b;
endmodule // GEQ_UNSIGNED
module CompareRecFN(
    input clock,
    input reset,
    input [64:0] io_a,
    input [64:0] io_b,
    input io_signaling,
    output io_lt,
    output io_eq,
    output io_gt,
    output [4:0] io_exceptionFlags
);
    wire [11:0] _T_16;
    BITS #(.width(65), .high(63), .low(52)) bits_1723 (
        .y(_T_16),
        .in(io_a)
    );
    wire [2:0] _T_17;
    BITS #(.width(12), .high(11), .low(9)) bits_1724 (
        .y(_T_17),
        .in(_T_16)
    );
    wire _T_19;
    wire [2:0] _WTEMP_219;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_1725 (
        .y(_WTEMP_219),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(3)) u_eq_1726 (
        .y(_T_19),
        .a(_T_17),
        .b(_WTEMP_219)
    );
    wire [1:0] _T_20;
    BITS #(.width(12), .high(11), .low(10)) bits_1727 (
        .y(_T_20),
        .in(_T_16)
    );
    wire _T_22;
    EQ_UNSIGNED #(.width(2)) u_eq_1728 (
        .y(_T_22),
        .a(_T_20),
        .b(2'h3)
    );
    wire rawA_sign;
    wire rawA_isNaN;
    wire rawA_isInf;
    wire rawA_isZero;
    wire [12:0] rawA_sExp;
    wire [55:0] rawA_sig;
    wire _T_36;
    BITS #(.width(65), .high(64), .low(64)) bits_1729 (
        .y(_T_36),
        .in(io_a)
    );
    wire _T_37;
    BITS #(.width(12), .high(9), .low(9)) bits_1730 (
        .y(_T_37),
        .in(_T_16)
    );
    wire _T_38;
    BITWISEAND #(.width(1)) bitwiseand_1731 (
        .y(_T_38),
        .a(_T_22),
        .b(_T_37)
    );
    wire _T_39;
    BITS #(.width(12), .high(9), .low(9)) bits_1732 (
        .y(_T_39),
        .in(_T_16)
    );
    wire _T_41;
    EQ_UNSIGNED #(.width(1)) u_eq_1733 (
        .y(_T_41),
        .a(_T_39),
        .b(1'h0)
    );
    wire _T_42;
    BITWISEAND #(.width(1)) bitwiseand_1734 (
        .y(_T_42),
        .a(_T_22),
        .b(_T_41)
    );
    wire [12:0] _T_43;
    CVT_UNSIGNED #(.width(12)) u_cvt_1735 (
        .y(_T_43),
        .in(_T_16)
    );
    wire _T_46;
    EQ_UNSIGNED #(.width(1)) u_eq_1736 (
        .y(_T_46),
        .a(_T_19),
        .b(1'h0)
    );
    wire [51:0] _T_47;
    BITS #(.width(65), .high(51), .low(0)) bits_1737 (
        .y(_T_47),
        .in(io_a)
    );
    wire [53:0] _T_49;
    CAT #(.width_a(52), .width_b(2)) cat_1738 (
        .y(_T_49),
        .a(_T_47),
        .b(2'h0)
    );
    wire [1:0] _T_50;
    CAT #(.width_a(1), .width_b(1)) cat_1739 (
        .y(_T_50),
        .a(1'h0),
        .b(_T_46)
    );
    wire [55:0] _T_51;
    CAT #(.width_a(2), .width_b(54)) cat_1740 (
        .y(_T_51),
        .a(_T_50),
        .b(_T_49)
    );
    wire [11:0] _T_52;
    BITS #(.width(65), .high(63), .low(52)) bits_1741 (
        .y(_T_52),
        .in(io_b)
    );
    wire [2:0] _T_53;
    BITS #(.width(12), .high(11), .low(9)) bits_1742 (
        .y(_T_53),
        .in(_T_52)
    );
    wire _T_55;
    wire [2:0] _WTEMP_220;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_1743 (
        .y(_WTEMP_220),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(3)) u_eq_1744 (
        .y(_T_55),
        .a(_T_53),
        .b(_WTEMP_220)
    );
    wire [1:0] _T_56;
    BITS #(.width(12), .high(11), .low(10)) bits_1745 (
        .y(_T_56),
        .in(_T_52)
    );
    wire _T_58;
    EQ_UNSIGNED #(.width(2)) u_eq_1746 (
        .y(_T_58),
        .a(_T_56),
        .b(2'h3)
    );
    wire rawB_sign;
    wire rawB_isNaN;
    wire rawB_isInf;
    wire rawB_isZero;
    wire [12:0] rawB_sExp;
    wire [55:0] rawB_sig;
    wire _T_72;
    BITS #(.width(65), .high(64), .low(64)) bits_1747 (
        .y(_T_72),
        .in(io_b)
    );
    wire _T_73;
    BITS #(.width(12), .high(9), .low(9)) bits_1748 (
        .y(_T_73),
        .in(_T_52)
    );
    wire _T_74;
    BITWISEAND #(.width(1)) bitwiseand_1749 (
        .y(_T_74),
        .a(_T_58),
        .b(_T_73)
    );
    wire _T_75;
    BITS #(.width(12), .high(9), .low(9)) bits_1750 (
        .y(_T_75),
        .in(_T_52)
    );
    wire _T_77;
    EQ_UNSIGNED #(.width(1)) u_eq_1751 (
        .y(_T_77),
        .a(_T_75),
        .b(1'h0)
    );
    wire _T_78;
    BITWISEAND #(.width(1)) bitwiseand_1752 (
        .y(_T_78),
        .a(_T_58),
        .b(_T_77)
    );
    wire [12:0] _T_79;
    CVT_UNSIGNED #(.width(12)) u_cvt_1753 (
        .y(_T_79),
        .in(_T_52)
    );
    wire _T_82;
    EQ_UNSIGNED #(.width(1)) u_eq_1754 (
        .y(_T_82),
        .a(_T_55),
        .b(1'h0)
    );
    wire [51:0] _T_83;
    BITS #(.width(65), .high(51), .low(0)) bits_1755 (
        .y(_T_83),
        .in(io_b)
    );
    wire [53:0] _T_85;
    CAT #(.width_a(52), .width_b(2)) cat_1756 (
        .y(_T_85),
        .a(_T_83),
        .b(2'h0)
    );
    wire [1:0] _T_86;
    CAT #(.width_a(1), .width_b(1)) cat_1757 (
        .y(_T_86),
        .a(1'h0),
        .b(_T_82)
    );
    wire [55:0] _T_87;
    CAT #(.width_a(2), .width_b(54)) cat_1758 (
        .y(_T_87),
        .a(_T_86),
        .b(_T_85)
    );
    wire _T_89;
    EQ_UNSIGNED #(.width(1)) u_eq_1759 (
        .y(_T_89),
        .a(rawA_isNaN),
        .b(1'h0)
    );
    wire _T_91;
    EQ_UNSIGNED #(.width(1)) u_eq_1760 (
        .y(_T_91),
        .a(rawB_isNaN),
        .b(1'h0)
    );
    wire ordered;
    BITWISEAND #(.width(1)) bitwiseand_1761 (
        .y(ordered),
        .a(_T_89),
        .b(_T_91)
    );
    wire bothInfs;
    BITWISEAND #(.width(1)) bitwiseand_1762 (
        .y(bothInfs),
        .a(rawA_isInf),
        .b(rawB_isInf)
    );
    wire bothZeros;
    BITWISEAND #(.width(1)) bitwiseand_1763 (
        .y(bothZeros),
        .a(rawA_isZero),
        .b(rawB_isZero)
    );
    wire eqExps;
    EQ_SIGNED #(.width(13)) s_eq_1764 (
        .y(eqExps),
        .a(rawA_sExp),
        .b(rawB_sExp)
    );
    wire _T_92;
    LT_SIGNED #(.width(13)) s_lt_1765 (
        .y(_T_92),
        .a(rawA_sExp),
        .b(rawB_sExp)
    );
    wire _T_93;
    LT_UNSIGNED #(.width(56)) u_lt_1766 (
        .y(_T_93),
        .a(rawA_sig),
        .b(rawB_sig)
    );
    wire _T_94;
    BITWISEAND #(.width(1)) bitwiseand_1767 (
        .y(_T_94),
        .a(eqExps),
        .b(_T_93)
    );
    wire common_ltMags;
    BITWISEOR #(.width(1)) bitwiseor_1768 (
        .y(common_ltMags),
        .a(_T_92),
        .b(_T_94)
    );
    wire _T_95;
    EQ_UNSIGNED #(.width(56)) u_eq_1769 (
        .y(_T_95),
        .a(rawA_sig),
        .b(rawB_sig)
    );
    wire common_eqMags;
    BITWISEAND #(.width(1)) bitwiseand_1770 (
        .y(common_eqMags),
        .a(eqExps),
        .b(_T_95)
    );
    wire _T_97;
    EQ_UNSIGNED #(.width(1)) u_eq_1771 (
        .y(_T_97),
        .a(bothZeros),
        .b(1'h0)
    );
    wire _T_99;
    EQ_UNSIGNED #(.width(1)) u_eq_1772 (
        .y(_T_99),
        .a(rawB_sign),
        .b(1'h0)
    );
    wire _T_100;
    BITWISEAND #(.width(1)) bitwiseand_1773 (
        .y(_T_100),
        .a(rawA_sign),
        .b(_T_99)
    );
    wire _T_102;
    EQ_UNSIGNED #(.width(1)) u_eq_1774 (
        .y(_T_102),
        .a(bothInfs),
        .b(1'h0)
    );
    wire _T_104;
    EQ_UNSIGNED #(.width(1)) u_eq_1775 (
        .y(_T_104),
        .a(common_ltMags),
        .b(1'h0)
    );
    wire _T_105;
    BITWISEAND #(.width(1)) bitwiseand_1776 (
        .y(_T_105),
        .a(rawA_sign),
        .b(_T_104)
    );
    wire _T_107;
    EQ_UNSIGNED #(.width(1)) u_eq_1777 (
        .y(_T_107),
        .a(common_eqMags),
        .b(1'h0)
    );
    wire _T_108;
    BITWISEAND #(.width(1)) bitwiseand_1778 (
        .y(_T_108),
        .a(_T_105),
        .b(_T_107)
    );
    wire _T_110;
    EQ_UNSIGNED #(.width(1)) u_eq_1779 (
        .y(_T_110),
        .a(rawB_sign),
        .b(1'h0)
    );
    wire _T_111;
    BITWISEAND #(.width(1)) bitwiseand_1780 (
        .y(_T_111),
        .a(_T_110),
        .b(common_ltMags)
    );
    wire _T_112;
    BITWISEOR #(.width(1)) bitwiseor_1781 (
        .y(_T_112),
        .a(_T_108),
        .b(_T_111)
    );
    wire _T_113;
    BITWISEAND #(.width(1)) bitwiseand_1782 (
        .y(_T_113),
        .a(_T_102),
        .b(_T_112)
    );
    wire _T_114;
    BITWISEOR #(.width(1)) bitwiseor_1783 (
        .y(_T_114),
        .a(_T_100),
        .b(_T_113)
    );
    wire ordered_lt;
    BITWISEAND #(.width(1)) bitwiseand_1784 (
        .y(ordered_lt),
        .a(_T_97),
        .b(_T_114)
    );
    wire _T_115;
    EQ_UNSIGNED #(.width(1)) u_eq_1785 (
        .y(_T_115),
        .a(rawA_sign),
        .b(rawB_sign)
    );
    wire _T_116;
    BITWISEOR #(.width(1)) bitwiseor_1786 (
        .y(_T_116),
        .a(bothInfs),
        .b(common_eqMags)
    );
    wire _T_117;
    BITWISEAND #(.width(1)) bitwiseand_1787 (
        .y(_T_117),
        .a(_T_115),
        .b(_T_116)
    );
    wire ordered_eq;
    BITWISEOR #(.width(1)) bitwiseor_1788 (
        .y(ordered_eq),
        .a(bothZeros),
        .b(_T_117)
    );
    wire _T_118;
    BITS #(.width(56), .high(53), .low(53)) bits_1789 (
        .y(_T_118),
        .in(rawA_sig)
    );
    wire _T_120;
    EQ_UNSIGNED #(.width(1)) u_eq_1790 (
        .y(_T_120),
        .a(_T_118),
        .b(1'h0)
    );
    wire _T_121;
    BITWISEAND #(.width(1)) bitwiseand_1791 (
        .y(_T_121),
        .a(rawA_isNaN),
        .b(_T_120)
    );
    wire _T_122;
    BITS #(.width(56), .high(53), .low(53)) bits_1792 (
        .y(_T_122),
        .in(rawB_sig)
    );
    wire _T_124;
    EQ_UNSIGNED #(.width(1)) u_eq_1793 (
        .y(_T_124),
        .a(_T_122),
        .b(1'h0)
    );
    wire _T_125;
    BITWISEAND #(.width(1)) bitwiseand_1794 (
        .y(_T_125),
        .a(rawB_isNaN),
        .b(_T_124)
    );
    wire _T_126;
    BITWISEOR #(.width(1)) bitwiseor_1795 (
        .y(_T_126),
        .a(_T_121),
        .b(_T_125)
    );
    wire _T_128;
    EQ_UNSIGNED #(.width(1)) u_eq_1796 (
        .y(_T_128),
        .a(ordered),
        .b(1'h0)
    );
    wire _T_129;
    BITWISEAND #(.width(1)) bitwiseand_1797 (
        .y(_T_129),
        .a(io_signaling),
        .b(_T_128)
    );
    wire invalid;
    BITWISEOR #(.width(1)) bitwiseor_1798 (
        .y(invalid),
        .a(_T_126),
        .b(_T_129)
    );
    wire _T_130;
    BITWISEAND #(.width(1)) bitwiseand_1799 (
        .y(_T_130),
        .a(ordered),
        .b(ordered_lt)
    );
    wire _T_131;
    BITWISEAND #(.width(1)) bitwiseand_1800 (
        .y(_T_131),
        .a(ordered),
        .b(ordered_eq)
    );
    wire _T_133;
    EQ_UNSIGNED #(.width(1)) u_eq_1801 (
        .y(_T_133),
        .a(ordered_lt),
        .b(1'h0)
    );
    wire _T_134;
    BITWISEAND #(.width(1)) bitwiseand_1802 (
        .y(_T_134),
        .a(ordered),
        .b(_T_133)
    );
    wire _T_136;
    EQ_UNSIGNED #(.width(1)) u_eq_1803 (
        .y(_T_136),
        .a(ordered_eq),
        .b(1'h0)
    );
    wire _T_137;
    BITWISEAND #(.width(1)) bitwiseand_1804 (
        .y(_T_137),
        .a(_T_134),
        .b(_T_136)
    );
    wire [4:0] _T_139;
    CAT #(.width_a(1), .width_b(4)) cat_1805 (
        .y(_T_139),
        .a(invalid),
        .b(4'h0)
    );
    assign io_eq = _T_131;
    assign io_exceptionFlags = _T_139;
    assign io_gt = _T_137;
    assign io_lt = _T_130;
    assign rawA_isInf = _T_42;
    assign rawA_isNaN = _T_38;
    assign rawA_isZero = _T_19;
    assign rawA_sExp = _T_43;
    assign rawA_sig = _T_51;
    assign rawA_sign = _T_36;
    assign rawB_isInf = _T_78;
    assign rawB_isNaN = _T_74;
    assign rawB_isZero = _T_55;
    assign rawB_sExp = _T_79;
    assign rawB_sig = _T_87;
    assign rawB_sign = _T_72;
endmodule //CompareRecFN
module CVT_UNSIGNED(y, in);
    parameter width = 4;
    output [width:0] y;
    input [width-1:0] in;
    assign y = $signed({1'b0, in});
endmodule // CVT_UNSIGNED
module EQ_SIGNED(y, a, b);
    parameter width = 4;
    output y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = $signed(a) == $signed(b);
endmodule // EQ_SIGNED
module LT_SIGNED(y, a, b);
    parameter width = 4;
    output y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = $signed(a) < $signed(b);
endmodule // LT_SIGNED
module RecFNToIN(
    input clock,
    input reset,
    input [64:0] io_in,
    input [1:0] io_roundingMode,
    input io_signedOut,
    output [31:0] io_out,
    output [2:0] io_intExceptionFlags
);
    wire sign;
    BITS #(.width(65), .high(64), .low(64)) bits_1825 (
        .y(sign),
        .in(io_in)
    );
    wire [11:0] exp;
    BITS #(.width(65), .high(63), .low(52)) bits_1826 (
        .y(exp),
        .in(io_in)
    );
    wire [51:0] fract;
    BITS #(.width(65), .high(51), .low(0)) bits_1827 (
        .y(fract),
        .in(io_in)
    );
    wire [2:0] _T_12;
    BITS #(.width(12), .high(11), .low(9)) bits_1828 (
        .y(_T_12),
        .in(exp)
    );
    wire isZero;
    wire [2:0] _WTEMP_228;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_1829 (
        .y(_WTEMP_228),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(3)) u_eq_1830 (
        .y(isZero),
        .a(_T_12),
        .b(_WTEMP_228)
    );
    wire [1:0] _T_14;
    BITS #(.width(12), .high(11), .low(10)) bits_1831 (
        .y(_T_14),
        .in(exp)
    );
    wire invalid;
    EQ_UNSIGNED #(.width(2)) u_eq_1832 (
        .y(invalid),
        .a(_T_14),
        .b(2'h3)
    );
    wire _T_16;
    BITS #(.width(12), .high(9), .low(9)) bits_1833 (
        .y(_T_16),
        .in(exp)
    );
    wire isNaN;
    BITWISEAND #(.width(1)) bitwiseand_1834 (
        .y(isNaN),
        .a(invalid),
        .b(_T_16)
    );
    wire notSpecial_magGeOne;
    BITS #(.width(12), .high(11), .low(11)) bits_1835 (
        .y(notSpecial_magGeOne),
        .in(exp)
    );
    wire [52:0] _T_17;
    CAT #(.width_a(1), .width_b(52)) cat_1836 (
        .y(_T_17),
        .a(notSpecial_magGeOne),
        .b(fract)
    );
    wire [4:0] _T_18;
    BITS #(.width(12), .high(4), .low(0)) bits_1837 (
        .y(_T_18),
        .in(exp)
    );
    wire [4:0] _T_20;
    wire [4:0] _WTEMP_229;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_1838 (
        .y(_WTEMP_229),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(5)) u_mux_1839 (
        .y(_T_20),
        .sel(notSpecial_magGeOne),
        .a(_T_18),
        .b(_WTEMP_229)
    );
    wire [83:0] shiftedSig;
    DSHL_UNSIGNED #(.width_in(53), .width_n(5)) u_dshl_1840 (
        .y(shiftedSig),
        .in(_T_17),
        .n(_T_20)
    );
    wire [31:0] unroundedInt;
    BITS #(.width(84), .high(83), .low(52)) bits_1841 (
        .y(unroundedInt),
        .in(shiftedSig)
    );
    wire [1:0] _T_21;
    BITS #(.width(84), .high(52), .low(51)) bits_1842 (
        .y(_T_21),
        .in(shiftedSig)
    );
    wire [50:0] _T_22;
    BITS #(.width(84), .high(50), .low(0)) bits_1843 (
        .y(_T_22),
        .in(shiftedSig)
    );
    wire _T_24;
    wire [50:0] _WTEMP_230;
    PAD_UNSIGNED #(.width(1), .n(51)) u_pad_1844 (
        .y(_WTEMP_230),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(51)) u_neq_1845 (
        .y(_T_24),
        .a(_T_22),
        .b(_WTEMP_230)
    );
    wire [2:0] roundBits;
    CAT #(.width_a(2), .width_b(1)) cat_1846 (
        .y(roundBits),
        .a(_T_21),
        .b(_T_24)
    );
    wire [1:0] _T_25;
    BITS #(.width(3), .high(1), .low(0)) bits_1847 (
        .y(_T_25),
        .in(roundBits)
    );
    wire _T_27;
    wire [1:0] _WTEMP_231;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_1848 (
        .y(_WTEMP_231),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(2)) u_neq_1849 (
        .y(_T_27),
        .a(_T_25),
        .b(_WTEMP_231)
    );
    wire _T_29;
    EQ_UNSIGNED #(.width(1)) u_eq_1850 (
        .y(_T_29),
        .a(isZero),
        .b(1'h0)
    );
    wire roundInexact;
    MUX_UNSIGNED #(.width(1)) u_mux_1851 (
        .y(roundInexact),
        .sel(notSpecial_magGeOne),
        .a(_T_27),
        .b(_T_29)
    );
    wire [1:0] _T_30;
    BITS #(.width(3), .high(2), .low(1)) bits_1852 (
        .y(_T_30),
        .in(roundBits)
    );
    wire [1:0] _T_31;
    BITWISENOT #(.width(2)) bitwisenot_1853 (
        .y(_T_31),
        .in(_T_30)
    );
    wire _T_33;
    wire [1:0] _WTEMP_232;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_1854 (
        .y(_WTEMP_232),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(2)) u_eq_1855 (
        .y(_T_33),
        .a(_T_31),
        .b(_WTEMP_232)
    );
    wire [1:0] _T_34;
    BITS #(.width(3), .high(1), .low(0)) bits_1856 (
        .y(_T_34),
        .in(roundBits)
    );
    wire [1:0] _T_35;
    BITWISENOT #(.width(2)) bitwisenot_1857 (
        .y(_T_35),
        .in(_T_34)
    );
    wire _T_37;
    wire [1:0] _WTEMP_233;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_1858 (
        .y(_WTEMP_233),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(2)) u_eq_1859 (
        .y(_T_37),
        .a(_T_35),
        .b(_WTEMP_233)
    );
    wire _T_38;
    BITWISEOR #(.width(1)) bitwiseor_1860 (
        .y(_T_38),
        .a(_T_33),
        .b(_T_37)
    );
    wire [10:0] _T_39;
    BITS #(.width(12), .high(10), .low(0)) bits_1861 (
        .y(_T_39),
        .in(exp)
    );
    wire [10:0] _T_40;
    BITWISENOT #(.width(11)) bitwisenot_1862 (
        .y(_T_40),
        .in(_T_39)
    );
    wire _T_42;
    wire [10:0] _WTEMP_234;
    PAD_UNSIGNED #(.width(1), .n(11)) u_pad_1863 (
        .y(_WTEMP_234),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(11)) u_eq_1864 (
        .y(_T_42),
        .a(_T_40),
        .b(_WTEMP_234)
    );
    wire [1:0] _T_43;
    BITS #(.width(3), .high(1), .low(0)) bits_1865 (
        .y(_T_43),
        .in(roundBits)
    );
    wire _T_45;
    wire [1:0] _WTEMP_235;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_1866 (
        .y(_WTEMP_235),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(2)) u_neq_1867 (
        .y(_T_45),
        .a(_T_43),
        .b(_WTEMP_235)
    );
    wire _T_47;
    MUX_UNSIGNED #(.width(1)) u_mux_1868 (
        .y(_T_47),
        .sel(_T_42),
        .a(_T_45),
        .b(1'h0)
    );
    wire roundIncr_nearestEven;
    MUX_UNSIGNED #(.width(1)) u_mux_1869 (
        .y(roundIncr_nearestEven),
        .sel(notSpecial_magGeOne),
        .a(_T_38),
        .b(_T_47)
    );
    wire _T_48;
    EQ_UNSIGNED #(.width(2)) u_eq_1870 (
        .y(_T_48),
        .a(io_roundingMode),
        .b(2'h0)
    );
    wire _T_49;
    BITWISEAND #(.width(1)) bitwiseand_1871 (
        .y(_T_49),
        .a(_T_48),
        .b(roundIncr_nearestEven)
    );
    wire _T_50;
    EQ_UNSIGNED #(.width(2)) u_eq_1872 (
        .y(_T_50),
        .a(io_roundingMode),
        .b(2'h2)
    );
    wire _T_51;
    BITWISEAND #(.width(1)) bitwiseand_1873 (
        .y(_T_51),
        .a(sign),
        .b(roundInexact)
    );
    wire _T_52;
    BITWISEAND #(.width(1)) bitwiseand_1874 (
        .y(_T_52),
        .a(_T_50),
        .b(_T_51)
    );
    wire _T_53;
    BITWISEOR #(.width(1)) bitwiseor_1875 (
        .y(_T_53),
        .a(_T_49),
        .b(_T_52)
    );
    wire _T_54;
    EQ_UNSIGNED #(.width(2)) u_eq_1876 (
        .y(_T_54),
        .a(io_roundingMode),
        .b(2'h3)
    );
    wire _T_56;
    EQ_UNSIGNED #(.width(1)) u_eq_1877 (
        .y(_T_56),
        .a(sign),
        .b(1'h0)
    );
    wire _T_57;
    BITWISEAND #(.width(1)) bitwiseand_1878 (
        .y(_T_57),
        .a(_T_56),
        .b(roundInexact)
    );
    wire _T_58;
    BITWISEAND #(.width(1)) bitwiseand_1879 (
        .y(_T_58),
        .a(_T_54),
        .b(_T_57)
    );
    wire roundIncr;
    BITWISEOR #(.width(1)) bitwiseor_1880 (
        .y(roundIncr),
        .a(_T_53),
        .b(_T_58)
    );
    wire [31:0] _T_59;
    BITWISENOT #(.width(32)) bitwisenot_1881 (
        .y(_T_59),
        .in(unroundedInt)
    );
    wire [31:0] complUnroundedInt;
    MUX_UNSIGNED #(.width(32)) u_mux_1882 (
        .y(complUnroundedInt),
        .sel(sign),
        .a(_T_59),
        .b(unroundedInt)
    );
    wire _T_60;
    BITWISEXOR #(.width(1)) bitwisexor_1883 (
        .y(_T_60),
        .a(roundIncr),
        .b(sign)
    );
    wire [32:0] _T_62;
    wire [31:0] _WTEMP_236;
    PAD_UNSIGNED #(.width(1), .n(32)) u_pad_1884 (
        .y(_WTEMP_236),
        .in(1'h1)
    );
    ADD_UNSIGNED #(.width(32)) u_add_1885 (
        .y(_T_62),
        .a(complUnroundedInt),
        .b(_WTEMP_236)
    );
    wire [31:0] _T_63;
    TAIL #(.width(33), .n(1)) tail_1886 (
        .y(_T_63),
        .in(_T_62)
    );
    wire [31:0] roundedInt;
    MUX_UNSIGNED #(.width(32)) u_mux_1887 (
        .y(roundedInt),
        .sel(_T_60),
        .a(_T_63),
        .b(complUnroundedInt)
    );
    wire [29:0] _T_64;
    BITS #(.width(32), .high(29), .low(0)) bits_1888 (
        .y(_T_64),
        .in(unroundedInt)
    );
    wire [29:0] _T_65;
    BITWISENOT #(.width(30)) bitwisenot_1889 (
        .y(_T_65),
        .in(_T_64)
    );
    wire _T_67;
    wire [29:0] _WTEMP_237;
    PAD_UNSIGNED #(.width(1), .n(30)) u_pad_1890 (
        .y(_WTEMP_237),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(30)) u_eq_1891 (
        .y(_T_67),
        .a(_T_65),
        .b(_WTEMP_237)
    );
    wire roundCarryBut2;
    BITWISEAND #(.width(1)) bitwiseand_1892 (
        .y(roundCarryBut2),
        .a(_T_67),
        .b(roundIncr)
    );
    wire [10:0] posExp;
    BITS #(.width(12), .high(10), .low(0)) bits_1893 (
        .y(posExp),
        .in(exp)
    );
    wire _T_69;
    wire [10:0] _WTEMP_238;
    PAD_UNSIGNED #(.width(6), .n(11)) u_pad_1894 (
        .y(_WTEMP_238),
        .in(6'h20)
    );
    GEQ_UNSIGNED #(.width(11)) u_geq_1895 (
        .y(_T_69),
        .a(posExp),
        .b(_WTEMP_238)
    );
    wire _T_71;
    wire [10:0] _WTEMP_239;
    PAD_UNSIGNED #(.width(5), .n(11)) u_pad_1896 (
        .y(_WTEMP_239),
        .in(5'h1F)
    );
    EQ_UNSIGNED #(.width(11)) u_eq_1897 (
        .y(_T_71),
        .a(posExp),
        .b(_WTEMP_239)
    );
    wire _T_73;
    EQ_UNSIGNED #(.width(1)) u_eq_1898 (
        .y(_T_73),
        .a(sign),
        .b(1'h0)
    );
    wire [30:0] _T_74;
    BITS #(.width(32), .high(30), .low(0)) bits_1899 (
        .y(_T_74),
        .in(unroundedInt)
    );
    wire _T_76;
    wire [30:0] _WTEMP_240;
    PAD_UNSIGNED #(.width(1), .n(31)) u_pad_1900 (
        .y(_WTEMP_240),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(31)) u_neq_1901 (
        .y(_T_76),
        .a(_T_74),
        .b(_WTEMP_240)
    );
    wire _T_77;
    BITWISEOR #(.width(1)) bitwiseor_1902 (
        .y(_T_77),
        .a(_T_73),
        .b(_T_76)
    );
    wire _T_78;
    BITWISEOR #(.width(1)) bitwiseor_1903 (
        .y(_T_78),
        .a(_T_77),
        .b(roundIncr)
    );
    wire _T_79;
    BITWISEAND #(.width(1)) bitwiseand_1904 (
        .y(_T_79),
        .a(_T_71),
        .b(_T_78)
    );
    wire _T_80;
    BITWISEOR #(.width(1)) bitwiseor_1905 (
        .y(_T_80),
        .a(_T_69),
        .b(_T_79)
    );
    wire _T_82;
    EQ_UNSIGNED #(.width(1)) u_eq_1906 (
        .y(_T_82),
        .a(sign),
        .b(1'h0)
    );
    wire _T_84;
    wire [10:0] _WTEMP_241;
    PAD_UNSIGNED #(.width(5), .n(11)) u_pad_1907 (
        .y(_WTEMP_241),
        .in(5'h1E)
    );
    EQ_UNSIGNED #(.width(11)) u_eq_1908 (
        .y(_T_84),
        .a(posExp),
        .b(_WTEMP_241)
    );
    wire _T_85;
    BITWISEAND #(.width(1)) bitwiseand_1909 (
        .y(_T_85),
        .a(_T_82),
        .b(_T_84)
    );
    wire _T_86;
    BITWISEAND #(.width(1)) bitwiseand_1910 (
        .y(_T_86),
        .a(_T_85),
        .b(roundCarryBut2)
    );
    wire _T_87;
    BITWISEOR #(.width(1)) bitwiseor_1911 (
        .y(_T_87),
        .a(_T_80),
        .b(_T_86)
    );
    wire overflow_signed;
    MUX_UNSIGNED #(.width(1)) u_mux_1912 (
        .y(overflow_signed),
        .sel(notSpecial_magGeOne),
        .a(_T_87),
        .b(1'h0)
    );
    wire _T_90;
    wire [10:0] _WTEMP_242;
    PAD_UNSIGNED #(.width(6), .n(11)) u_pad_1913 (
        .y(_WTEMP_242),
        .in(6'h20)
    );
    GEQ_UNSIGNED #(.width(11)) u_geq_1914 (
        .y(_T_90),
        .a(posExp),
        .b(_WTEMP_242)
    );
    wire _T_91;
    BITWISEOR #(.width(1)) bitwiseor_1915 (
        .y(_T_91),
        .a(sign),
        .b(_T_90)
    );
    wire _T_93;
    wire [10:0] _WTEMP_243;
    PAD_UNSIGNED #(.width(5), .n(11)) u_pad_1916 (
        .y(_WTEMP_243),
        .in(5'h1F)
    );
    EQ_UNSIGNED #(.width(11)) u_eq_1917 (
        .y(_T_93),
        .a(posExp),
        .b(_WTEMP_243)
    );
    wire _T_94;
    BITS #(.width(32), .high(30), .low(30)) bits_1918 (
        .y(_T_94),
        .in(unroundedInt)
    );
    wire _T_95;
    BITWISEAND #(.width(1)) bitwiseand_1919 (
        .y(_T_95),
        .a(_T_93),
        .b(_T_94)
    );
    wire _T_96;
    BITWISEAND #(.width(1)) bitwiseand_1920 (
        .y(_T_96),
        .a(_T_95),
        .b(roundCarryBut2)
    );
    wire _T_97;
    BITWISEOR #(.width(1)) bitwiseor_1921 (
        .y(_T_97),
        .a(_T_91),
        .b(_T_96)
    );
    wire _T_98;
    BITWISEAND #(.width(1)) bitwiseand_1922 (
        .y(_T_98),
        .a(sign),
        .b(roundIncr)
    );
    wire overflow_unsigned;
    MUX_UNSIGNED #(.width(1)) u_mux_1923 (
        .y(overflow_unsigned),
        .sel(notSpecial_magGeOne),
        .a(_T_97),
        .b(_T_98)
    );
    wire overflow;
    MUX_UNSIGNED #(.width(1)) u_mux_1924 (
        .y(overflow),
        .sel(io_signedOut),
        .a(overflow_signed),
        .b(overflow_unsigned)
    );
    wire _T_100;
    EQ_UNSIGNED #(.width(1)) u_eq_1925 (
        .y(_T_100),
        .a(isNaN),
        .b(1'h0)
    );
    wire excSign;
    BITWISEAND #(.width(1)) bitwiseand_1926 (
        .y(excSign),
        .a(sign),
        .b(_T_100)
    );
    wire _T_101;
    BITWISEAND #(.width(1)) bitwiseand_1927 (
        .y(_T_101),
        .a(io_signedOut),
        .b(excSign)
    );
    wire [31:0] _T_103;
    assign _T_103 = 32'h80000000;
    wire [31:0] _T_105;
    wire [31:0] _WTEMP_244;
    PAD_UNSIGNED #(.width(1), .n(32)) u_pad_1928 (
        .y(_WTEMP_244),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(32)) u_mux_1929 (
        .y(_T_105),
        .sel(_T_101),
        .a(_T_103),
        .b(_WTEMP_244)
    );
    wire _T_107;
    EQ_UNSIGNED #(.width(1)) u_eq_1930 (
        .y(_T_107),
        .a(excSign),
        .b(1'h0)
    );
    wire _T_108;
    BITWISEAND #(.width(1)) bitwiseand_1931 (
        .y(_T_108),
        .a(io_signedOut),
        .b(_T_107)
    );
    wire [30:0] _T_111;
    wire [30:0] _WTEMP_245;
    PAD_UNSIGNED #(.width(1), .n(31)) u_pad_1932 (
        .y(_WTEMP_245),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(31)) u_mux_1933 (
        .y(_T_111),
        .sel(_T_108),
        .a(31'h7FFFFFFF),
        .b(_WTEMP_245)
    );
    wire [31:0] _T_112;
    wire [31:0] _WTEMP_246;
    PAD_UNSIGNED #(.width(31), .n(32)) u_pad_1934 (
        .y(_WTEMP_246),
        .in(_T_111)
    );
    BITWISEOR #(.width(32)) bitwiseor_1935 (
        .y(_T_112),
        .a(_T_105),
        .b(_WTEMP_246)
    );
    wire _T_114;
    EQ_UNSIGNED #(.width(1)) u_eq_1936 (
        .y(_T_114),
        .a(io_signedOut),
        .b(1'h0)
    );
    wire _T_116;
    EQ_UNSIGNED #(.width(1)) u_eq_1937 (
        .y(_T_116),
        .a(excSign),
        .b(1'h0)
    );
    wire _T_117;
    BITWISEAND #(.width(1)) bitwiseand_1938 (
        .y(_T_117),
        .a(_T_114),
        .b(_T_116)
    );
    wire [31:0] _T_120;
    wire [31:0] _WTEMP_247;
    PAD_UNSIGNED #(.width(1), .n(32)) u_pad_1939 (
        .y(_WTEMP_247),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(32)) u_mux_1940 (
        .y(_T_120),
        .sel(_T_117),
        .a(32'hFFFFFFFF),
        .b(_WTEMP_247)
    );
    wire [31:0] excValue;
    BITWISEOR #(.width(32)) bitwiseor_1941 (
        .y(excValue),
        .a(_T_112),
        .b(_T_120)
    );
    wire _T_122;
    EQ_UNSIGNED #(.width(1)) u_eq_1942 (
        .y(_T_122),
        .a(invalid),
        .b(1'h0)
    );
    wire _T_123;
    BITWISEAND #(.width(1)) bitwiseand_1943 (
        .y(_T_123),
        .a(roundInexact),
        .b(_T_122)
    );
    wire _T_125;
    EQ_UNSIGNED #(.width(1)) u_eq_1944 (
        .y(_T_125),
        .a(overflow),
        .b(1'h0)
    );
    wire inexact;
    BITWISEAND #(.width(1)) bitwiseand_1945 (
        .y(inexact),
        .a(_T_123),
        .b(_T_125)
    );
    wire _T_126;
    BITWISEOR #(.width(1)) bitwiseor_1946 (
        .y(_T_126),
        .a(invalid),
        .b(overflow)
    );
    wire [31:0] _T_127;
    MUX_UNSIGNED #(.width(32)) u_mux_1947 (
        .y(_T_127),
        .sel(_T_126),
        .a(excValue),
        .b(roundedInt)
    );
    wire [1:0] _T_128;
    CAT #(.width_a(1), .width_b(1)) cat_1948 (
        .y(_T_128),
        .a(invalid),
        .b(overflow)
    );
    wire [2:0] _T_129;
    CAT #(.width_a(2), .width_b(1)) cat_1949 (
        .y(_T_129),
        .a(_T_128),
        .b(inexact)
    );
    assign io_intExceptionFlags = _T_129;
    assign io_out = _T_127;
endmodule //RecFNToIN
module RecFNToIN_1(
    input clock,
    input reset,
    input [64:0] io_in,
    input [1:0] io_roundingMode,
    input io_signedOut,
    output [63:0] io_out,
    output [2:0] io_intExceptionFlags
);
    wire sign;
    BITS #(.width(65), .high(64), .low(64)) bits_1968 (
        .y(sign),
        .in(io_in)
    );
    wire [11:0] exp;
    BITS #(.width(65), .high(63), .low(52)) bits_1969 (
        .y(exp),
        .in(io_in)
    );
    wire [51:0] fract;
    BITS #(.width(65), .high(51), .low(0)) bits_1970 (
        .y(fract),
        .in(io_in)
    );
    wire [2:0] _T_12;
    BITS #(.width(12), .high(11), .low(9)) bits_1971 (
        .y(_T_12),
        .in(exp)
    );
    wire isZero;
    wire [2:0] _WTEMP_251;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_1972 (
        .y(_WTEMP_251),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(3)) u_eq_1973 (
        .y(isZero),
        .a(_T_12),
        .b(_WTEMP_251)
    );
    wire [1:0] _T_14;
    BITS #(.width(12), .high(11), .low(10)) bits_1974 (
        .y(_T_14),
        .in(exp)
    );
    wire invalid;
    EQ_UNSIGNED #(.width(2)) u_eq_1975 (
        .y(invalid),
        .a(_T_14),
        .b(2'h3)
    );
    wire _T_16;
    BITS #(.width(12), .high(9), .low(9)) bits_1976 (
        .y(_T_16),
        .in(exp)
    );
    wire isNaN;
    BITWISEAND #(.width(1)) bitwiseand_1977 (
        .y(isNaN),
        .a(invalid),
        .b(_T_16)
    );
    wire notSpecial_magGeOne;
    BITS #(.width(12), .high(11), .low(11)) bits_1978 (
        .y(notSpecial_magGeOne),
        .in(exp)
    );
    wire [52:0] _T_17;
    CAT #(.width_a(1), .width_b(52)) cat_1979 (
        .y(_T_17),
        .a(notSpecial_magGeOne),
        .b(fract)
    );
    wire [5:0] _T_18;
    BITS #(.width(12), .high(5), .low(0)) bits_1980 (
        .y(_T_18),
        .in(exp)
    );
    wire [5:0] _T_20;
    wire [5:0] _WTEMP_252;
    PAD_UNSIGNED #(.width(1), .n(6)) u_pad_1981 (
        .y(_WTEMP_252),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(6)) u_mux_1982 (
        .y(_T_20),
        .sel(notSpecial_magGeOne),
        .a(_T_18),
        .b(_WTEMP_252)
    );
    wire [115:0] shiftedSig;
    DSHL_UNSIGNED #(.width_in(53), .width_n(6)) u_dshl_1983 (
        .y(shiftedSig),
        .in(_T_17),
        .n(_T_20)
    );
    wire [63:0] unroundedInt;
    BITS #(.width(116), .high(115), .low(52)) bits_1984 (
        .y(unroundedInt),
        .in(shiftedSig)
    );
    wire [1:0] _T_21;
    BITS #(.width(116), .high(52), .low(51)) bits_1985 (
        .y(_T_21),
        .in(shiftedSig)
    );
    wire [50:0] _T_22;
    BITS #(.width(116), .high(50), .low(0)) bits_1986 (
        .y(_T_22),
        .in(shiftedSig)
    );
    wire _T_24;
    wire [50:0] _WTEMP_253;
    PAD_UNSIGNED #(.width(1), .n(51)) u_pad_1987 (
        .y(_WTEMP_253),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(51)) u_neq_1988 (
        .y(_T_24),
        .a(_T_22),
        .b(_WTEMP_253)
    );
    wire [2:0] roundBits;
    CAT #(.width_a(2), .width_b(1)) cat_1989 (
        .y(roundBits),
        .a(_T_21),
        .b(_T_24)
    );
    wire [1:0] _T_25;
    BITS #(.width(3), .high(1), .low(0)) bits_1990 (
        .y(_T_25),
        .in(roundBits)
    );
    wire _T_27;
    wire [1:0] _WTEMP_254;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_1991 (
        .y(_WTEMP_254),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(2)) u_neq_1992 (
        .y(_T_27),
        .a(_T_25),
        .b(_WTEMP_254)
    );
    wire _T_29;
    EQ_UNSIGNED #(.width(1)) u_eq_1993 (
        .y(_T_29),
        .a(isZero),
        .b(1'h0)
    );
    wire roundInexact;
    MUX_UNSIGNED #(.width(1)) u_mux_1994 (
        .y(roundInexact),
        .sel(notSpecial_magGeOne),
        .a(_T_27),
        .b(_T_29)
    );
    wire [1:0] _T_30;
    BITS #(.width(3), .high(2), .low(1)) bits_1995 (
        .y(_T_30),
        .in(roundBits)
    );
    wire [1:0] _T_31;
    BITWISENOT #(.width(2)) bitwisenot_1996 (
        .y(_T_31),
        .in(_T_30)
    );
    wire _T_33;
    wire [1:0] _WTEMP_255;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_1997 (
        .y(_WTEMP_255),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(2)) u_eq_1998 (
        .y(_T_33),
        .a(_T_31),
        .b(_WTEMP_255)
    );
    wire [1:0] _T_34;
    BITS #(.width(3), .high(1), .low(0)) bits_1999 (
        .y(_T_34),
        .in(roundBits)
    );
    wire [1:0] _T_35;
    BITWISENOT #(.width(2)) bitwisenot_2000 (
        .y(_T_35),
        .in(_T_34)
    );
    wire _T_37;
    wire [1:0] _WTEMP_256;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2001 (
        .y(_WTEMP_256),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(2)) u_eq_2002 (
        .y(_T_37),
        .a(_T_35),
        .b(_WTEMP_256)
    );
    wire _T_38;
    BITWISEOR #(.width(1)) bitwiseor_2003 (
        .y(_T_38),
        .a(_T_33),
        .b(_T_37)
    );
    wire [10:0] _T_39;
    BITS #(.width(12), .high(10), .low(0)) bits_2004 (
        .y(_T_39),
        .in(exp)
    );
    wire [10:0] _T_40;
    BITWISENOT #(.width(11)) bitwisenot_2005 (
        .y(_T_40),
        .in(_T_39)
    );
    wire _T_42;
    wire [10:0] _WTEMP_257;
    PAD_UNSIGNED #(.width(1), .n(11)) u_pad_2006 (
        .y(_WTEMP_257),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(11)) u_eq_2007 (
        .y(_T_42),
        .a(_T_40),
        .b(_WTEMP_257)
    );
    wire [1:0] _T_43;
    BITS #(.width(3), .high(1), .low(0)) bits_2008 (
        .y(_T_43),
        .in(roundBits)
    );
    wire _T_45;
    wire [1:0] _WTEMP_258;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2009 (
        .y(_WTEMP_258),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(2)) u_neq_2010 (
        .y(_T_45),
        .a(_T_43),
        .b(_WTEMP_258)
    );
    wire _T_47;
    MUX_UNSIGNED #(.width(1)) u_mux_2011 (
        .y(_T_47),
        .sel(_T_42),
        .a(_T_45),
        .b(1'h0)
    );
    wire roundIncr_nearestEven;
    MUX_UNSIGNED #(.width(1)) u_mux_2012 (
        .y(roundIncr_nearestEven),
        .sel(notSpecial_magGeOne),
        .a(_T_38),
        .b(_T_47)
    );
    wire _T_48;
    EQ_UNSIGNED #(.width(2)) u_eq_2013 (
        .y(_T_48),
        .a(io_roundingMode),
        .b(2'h0)
    );
    wire _T_49;
    BITWISEAND #(.width(1)) bitwiseand_2014 (
        .y(_T_49),
        .a(_T_48),
        .b(roundIncr_nearestEven)
    );
    wire _T_50;
    EQ_UNSIGNED #(.width(2)) u_eq_2015 (
        .y(_T_50),
        .a(io_roundingMode),
        .b(2'h2)
    );
    wire _T_51;
    BITWISEAND #(.width(1)) bitwiseand_2016 (
        .y(_T_51),
        .a(sign),
        .b(roundInexact)
    );
    wire _T_52;
    BITWISEAND #(.width(1)) bitwiseand_2017 (
        .y(_T_52),
        .a(_T_50),
        .b(_T_51)
    );
    wire _T_53;
    BITWISEOR #(.width(1)) bitwiseor_2018 (
        .y(_T_53),
        .a(_T_49),
        .b(_T_52)
    );
    wire _T_54;
    EQ_UNSIGNED #(.width(2)) u_eq_2019 (
        .y(_T_54),
        .a(io_roundingMode),
        .b(2'h3)
    );
    wire _T_56;
    EQ_UNSIGNED #(.width(1)) u_eq_2020 (
        .y(_T_56),
        .a(sign),
        .b(1'h0)
    );
    wire _T_57;
    BITWISEAND #(.width(1)) bitwiseand_2021 (
        .y(_T_57),
        .a(_T_56),
        .b(roundInexact)
    );
    wire _T_58;
    BITWISEAND #(.width(1)) bitwiseand_2022 (
        .y(_T_58),
        .a(_T_54),
        .b(_T_57)
    );
    wire roundIncr;
    BITWISEOR #(.width(1)) bitwiseor_2023 (
        .y(roundIncr),
        .a(_T_53),
        .b(_T_58)
    );
    wire [63:0] _T_59;
    BITWISENOT #(.width(64)) bitwisenot_2024 (
        .y(_T_59),
        .in(unroundedInt)
    );
    wire [63:0] complUnroundedInt;
    MUX_UNSIGNED #(.width(64)) u_mux_2025 (
        .y(complUnroundedInt),
        .sel(sign),
        .a(_T_59),
        .b(unroundedInt)
    );
    wire _T_60;
    BITWISEXOR #(.width(1)) bitwisexor_2026 (
        .y(_T_60),
        .a(roundIncr),
        .b(sign)
    );
    wire [64:0] _T_62;
    wire [63:0] _WTEMP_259;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_2027 (
        .y(_WTEMP_259),
        .in(1'h1)
    );
    ADD_UNSIGNED #(.width(64)) u_add_2028 (
        .y(_T_62),
        .a(complUnroundedInt),
        .b(_WTEMP_259)
    );
    wire [63:0] _T_63;
    TAIL #(.width(65), .n(1)) tail_2029 (
        .y(_T_63),
        .in(_T_62)
    );
    wire [63:0] roundedInt;
    MUX_UNSIGNED #(.width(64)) u_mux_2030 (
        .y(roundedInt),
        .sel(_T_60),
        .a(_T_63),
        .b(complUnroundedInt)
    );
    wire [61:0] _T_64;
    BITS #(.width(64), .high(61), .low(0)) bits_2031 (
        .y(_T_64),
        .in(unroundedInt)
    );
    wire [61:0] _T_65;
    BITWISENOT #(.width(62)) bitwisenot_2032 (
        .y(_T_65),
        .in(_T_64)
    );
    wire _T_67;
    wire [61:0] _WTEMP_260;
    PAD_UNSIGNED #(.width(1), .n(62)) u_pad_2033 (
        .y(_WTEMP_260),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(62)) u_eq_2034 (
        .y(_T_67),
        .a(_T_65),
        .b(_WTEMP_260)
    );
    wire roundCarryBut2;
    BITWISEAND #(.width(1)) bitwiseand_2035 (
        .y(roundCarryBut2),
        .a(_T_67),
        .b(roundIncr)
    );
    wire [10:0] posExp;
    BITS #(.width(12), .high(10), .low(0)) bits_2036 (
        .y(posExp),
        .in(exp)
    );
    wire _T_69;
    wire [10:0] _WTEMP_261;
    PAD_UNSIGNED #(.width(7), .n(11)) u_pad_2037 (
        .y(_WTEMP_261),
        .in(7'h40)
    );
    GEQ_UNSIGNED #(.width(11)) u_geq_2038 (
        .y(_T_69),
        .a(posExp),
        .b(_WTEMP_261)
    );
    wire _T_71;
    wire [10:0] _WTEMP_262;
    PAD_UNSIGNED #(.width(6), .n(11)) u_pad_2039 (
        .y(_WTEMP_262),
        .in(6'h3F)
    );
    EQ_UNSIGNED #(.width(11)) u_eq_2040 (
        .y(_T_71),
        .a(posExp),
        .b(_WTEMP_262)
    );
    wire _T_73;
    EQ_UNSIGNED #(.width(1)) u_eq_2041 (
        .y(_T_73),
        .a(sign),
        .b(1'h0)
    );
    wire [62:0] _T_74;
    BITS #(.width(64), .high(62), .low(0)) bits_2042 (
        .y(_T_74),
        .in(unroundedInt)
    );
    wire _T_76;
    wire [62:0] _WTEMP_263;
    PAD_UNSIGNED #(.width(1), .n(63)) u_pad_2043 (
        .y(_WTEMP_263),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(63)) u_neq_2044 (
        .y(_T_76),
        .a(_T_74),
        .b(_WTEMP_263)
    );
    wire _T_77;
    BITWISEOR #(.width(1)) bitwiseor_2045 (
        .y(_T_77),
        .a(_T_73),
        .b(_T_76)
    );
    wire _T_78;
    BITWISEOR #(.width(1)) bitwiseor_2046 (
        .y(_T_78),
        .a(_T_77),
        .b(roundIncr)
    );
    wire _T_79;
    BITWISEAND #(.width(1)) bitwiseand_2047 (
        .y(_T_79),
        .a(_T_71),
        .b(_T_78)
    );
    wire _T_80;
    BITWISEOR #(.width(1)) bitwiseor_2048 (
        .y(_T_80),
        .a(_T_69),
        .b(_T_79)
    );
    wire _T_82;
    EQ_UNSIGNED #(.width(1)) u_eq_2049 (
        .y(_T_82),
        .a(sign),
        .b(1'h0)
    );
    wire _T_84;
    wire [10:0] _WTEMP_264;
    PAD_UNSIGNED #(.width(6), .n(11)) u_pad_2050 (
        .y(_WTEMP_264),
        .in(6'h3E)
    );
    EQ_UNSIGNED #(.width(11)) u_eq_2051 (
        .y(_T_84),
        .a(posExp),
        .b(_WTEMP_264)
    );
    wire _T_85;
    BITWISEAND #(.width(1)) bitwiseand_2052 (
        .y(_T_85),
        .a(_T_82),
        .b(_T_84)
    );
    wire _T_86;
    BITWISEAND #(.width(1)) bitwiseand_2053 (
        .y(_T_86),
        .a(_T_85),
        .b(roundCarryBut2)
    );
    wire _T_87;
    BITWISEOR #(.width(1)) bitwiseor_2054 (
        .y(_T_87),
        .a(_T_80),
        .b(_T_86)
    );
    wire overflow_signed;
    MUX_UNSIGNED #(.width(1)) u_mux_2055 (
        .y(overflow_signed),
        .sel(notSpecial_magGeOne),
        .a(_T_87),
        .b(1'h0)
    );
    wire _T_90;
    wire [10:0] _WTEMP_265;
    PAD_UNSIGNED #(.width(7), .n(11)) u_pad_2056 (
        .y(_WTEMP_265),
        .in(7'h40)
    );
    GEQ_UNSIGNED #(.width(11)) u_geq_2057 (
        .y(_T_90),
        .a(posExp),
        .b(_WTEMP_265)
    );
    wire _T_91;
    BITWISEOR #(.width(1)) bitwiseor_2058 (
        .y(_T_91),
        .a(sign),
        .b(_T_90)
    );
    wire _T_93;
    wire [10:0] _WTEMP_266;
    PAD_UNSIGNED #(.width(6), .n(11)) u_pad_2059 (
        .y(_WTEMP_266),
        .in(6'h3F)
    );
    EQ_UNSIGNED #(.width(11)) u_eq_2060 (
        .y(_T_93),
        .a(posExp),
        .b(_WTEMP_266)
    );
    wire _T_94;
    BITS #(.width(64), .high(62), .low(62)) bits_2061 (
        .y(_T_94),
        .in(unroundedInt)
    );
    wire _T_95;
    BITWISEAND #(.width(1)) bitwiseand_2062 (
        .y(_T_95),
        .a(_T_93),
        .b(_T_94)
    );
    wire _T_96;
    BITWISEAND #(.width(1)) bitwiseand_2063 (
        .y(_T_96),
        .a(_T_95),
        .b(roundCarryBut2)
    );
    wire _T_97;
    BITWISEOR #(.width(1)) bitwiseor_2064 (
        .y(_T_97),
        .a(_T_91),
        .b(_T_96)
    );
    wire _T_98;
    BITWISEAND #(.width(1)) bitwiseand_2065 (
        .y(_T_98),
        .a(sign),
        .b(roundIncr)
    );
    wire overflow_unsigned;
    MUX_UNSIGNED #(.width(1)) u_mux_2066 (
        .y(overflow_unsigned),
        .sel(notSpecial_magGeOne),
        .a(_T_97),
        .b(_T_98)
    );
    wire overflow;
    MUX_UNSIGNED #(.width(1)) u_mux_2067 (
        .y(overflow),
        .sel(io_signedOut),
        .a(overflow_signed),
        .b(overflow_unsigned)
    );
    wire _T_100;
    EQ_UNSIGNED #(.width(1)) u_eq_2068 (
        .y(_T_100),
        .a(isNaN),
        .b(1'h0)
    );
    wire excSign;
    BITWISEAND #(.width(1)) bitwiseand_2069 (
        .y(excSign),
        .a(sign),
        .b(_T_100)
    );
    wire _T_101;
    BITWISEAND #(.width(1)) bitwiseand_2070 (
        .y(_T_101),
        .a(io_signedOut),
        .b(excSign)
    );
    wire [63:0] _T_103;
    assign _T_103 = 64'h8000000000000000;
    wire [63:0] _T_105;
    wire [63:0] _WTEMP_267;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_2071 (
        .y(_WTEMP_267),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_2072 (
        .y(_T_105),
        .sel(_T_101),
        .a(_T_103),
        .b(_WTEMP_267)
    );
    wire _T_107;
    EQ_UNSIGNED #(.width(1)) u_eq_2073 (
        .y(_T_107),
        .a(excSign),
        .b(1'h0)
    );
    wire _T_108;
    BITWISEAND #(.width(1)) bitwiseand_2074 (
        .y(_T_108),
        .a(io_signedOut),
        .b(_T_107)
    );
    wire [62:0] _T_111;
    wire [62:0] _WTEMP_268;
    PAD_UNSIGNED #(.width(1), .n(63)) u_pad_2075 (
        .y(_WTEMP_268),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(63)) u_mux_2076 (
        .y(_T_111),
        .sel(_T_108),
        .a(63'h7FFFFFFFFFFFFFFF),
        .b(_WTEMP_268)
    );
    wire [63:0] _T_112;
    wire [63:0] _WTEMP_269;
    PAD_UNSIGNED #(.width(63), .n(64)) u_pad_2077 (
        .y(_WTEMP_269),
        .in(_T_111)
    );
    BITWISEOR #(.width(64)) bitwiseor_2078 (
        .y(_T_112),
        .a(_T_105),
        .b(_WTEMP_269)
    );
    wire _T_114;
    EQ_UNSIGNED #(.width(1)) u_eq_2079 (
        .y(_T_114),
        .a(io_signedOut),
        .b(1'h0)
    );
    wire _T_116;
    EQ_UNSIGNED #(.width(1)) u_eq_2080 (
        .y(_T_116),
        .a(excSign),
        .b(1'h0)
    );
    wire _T_117;
    BITWISEAND #(.width(1)) bitwiseand_2081 (
        .y(_T_117),
        .a(_T_114),
        .b(_T_116)
    );
    wire [63:0] _T_120;
    wire [63:0] _WTEMP_270;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_2082 (
        .y(_WTEMP_270),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_2083 (
        .y(_T_120),
        .sel(_T_117),
        .a(64'hFFFFFFFFFFFFFFFF),
        .b(_WTEMP_270)
    );
    wire [63:0] excValue;
    BITWISEOR #(.width(64)) bitwiseor_2084 (
        .y(excValue),
        .a(_T_112),
        .b(_T_120)
    );
    wire _T_122;
    EQ_UNSIGNED #(.width(1)) u_eq_2085 (
        .y(_T_122),
        .a(invalid),
        .b(1'h0)
    );
    wire _T_123;
    BITWISEAND #(.width(1)) bitwiseand_2086 (
        .y(_T_123),
        .a(roundInexact),
        .b(_T_122)
    );
    wire _T_125;
    EQ_UNSIGNED #(.width(1)) u_eq_2087 (
        .y(_T_125),
        .a(overflow),
        .b(1'h0)
    );
    wire inexact;
    BITWISEAND #(.width(1)) bitwiseand_2088 (
        .y(inexact),
        .a(_T_123),
        .b(_T_125)
    );
    wire _T_126;
    BITWISEOR #(.width(1)) bitwiseor_2089 (
        .y(_T_126),
        .a(invalid),
        .b(overflow)
    );
    wire [63:0] _T_127;
    MUX_UNSIGNED #(.width(64)) u_mux_2090 (
        .y(_T_127),
        .sel(_T_126),
        .a(excValue),
        .b(roundedInt)
    );
    wire [1:0] _T_128;
    CAT #(.width_a(1), .width_b(1)) cat_2091 (
        .y(_T_128),
        .a(invalid),
        .b(overflow)
    );
    wire [2:0] _T_129;
    CAT #(.width_a(2), .width_b(1)) cat_2092 (
        .y(_T_129),
        .a(_T_128),
        .b(inexact)
    );
    assign io_intExceptionFlags = _T_129;
    assign io_out = _T_127;
endmodule //RecFNToIN_1
module IntToFP(
    input clock,
    input reset,
    input io_in_valid,
    input [4:0] io_in_bits_cmd,
    input io_in_bits_ldst,
    input io_in_bits_wen,
    input io_in_bits_ren1,
    input io_in_bits_ren2,
    input io_in_bits_ren3,
    input io_in_bits_swap12,
    input io_in_bits_swap23,
    input io_in_bits_single,
    input io_in_bits_fromint,
    input io_in_bits_toint,
    input io_in_bits_fastpipe,
    input io_in_bits_fma,
    input io_in_bits_div,
    input io_in_bits_sqrt,
    input io_in_bits_wflags,
    input [2:0] io_in_bits_rm,
    input [1:0] io_in_bits_typ,
    input [64:0] io_in_bits_in1,
    input [64:0] io_in_bits_in2,
    input [64:0] io_in_bits_in3,
    output io_out_valid,
    output [64:0] io_out_bits_data,
    output [4:0] io_out_bits_exc
);
    wire __T_132__q;
    wire __T_132__d;
    DFF_POSCLK #(.width(1)) _T_132 (
        .q(__T_132__q),
        .d(__T_132__d),
        .clk(clock)
    );
    wire _WTEMP_276;
    MUX_UNSIGNED #(.width(1)) u_mux_2146 (
        .y(__T_132__d),
        .sel(reset),
        .a(1'h0),
        .b(_WTEMP_276)
    );
    wire [4:0] __T_155_cmd__q;
    wire [4:0] __T_155_cmd__d;
    DFF_POSCLK #(.width(5)) _T_155_cmd (
        .q(__T_155_cmd__q),
        .d(__T_155_cmd__d),
        .clk(clock)
    );
    wire __T_155_ldst__q;
    wire __T_155_ldst__d;
    DFF_POSCLK #(.width(1)) _T_155_ldst (
        .q(__T_155_ldst__q),
        .d(__T_155_ldst__d),
        .clk(clock)
    );
    wire __T_155_wen__q;
    wire __T_155_wen__d;
    DFF_POSCLK #(.width(1)) _T_155_wen (
        .q(__T_155_wen__q),
        .d(__T_155_wen__d),
        .clk(clock)
    );
    wire __T_155_ren1__q;
    wire __T_155_ren1__d;
    DFF_POSCLK #(.width(1)) _T_155_ren1 (
        .q(__T_155_ren1__q),
        .d(__T_155_ren1__d),
        .clk(clock)
    );
    wire __T_155_ren2__q;
    wire __T_155_ren2__d;
    DFF_POSCLK #(.width(1)) _T_155_ren2 (
        .q(__T_155_ren2__q),
        .d(__T_155_ren2__d),
        .clk(clock)
    );
    wire __T_155_ren3__q;
    wire __T_155_ren3__d;
    DFF_POSCLK #(.width(1)) _T_155_ren3 (
        .q(__T_155_ren3__q),
        .d(__T_155_ren3__d),
        .clk(clock)
    );
    wire __T_155_swap12__q;
    wire __T_155_swap12__d;
    DFF_POSCLK #(.width(1)) _T_155_swap12 (
        .q(__T_155_swap12__q),
        .d(__T_155_swap12__d),
        .clk(clock)
    );
    wire __T_155_swap23__q;
    wire __T_155_swap23__d;
    DFF_POSCLK #(.width(1)) _T_155_swap23 (
        .q(__T_155_swap23__q),
        .d(__T_155_swap23__d),
        .clk(clock)
    );
    wire __T_155_single__q;
    wire __T_155_single__d;
    DFF_POSCLK #(.width(1)) _T_155_single (
        .q(__T_155_single__q),
        .d(__T_155_single__d),
        .clk(clock)
    );
    wire __T_155_fromint__q;
    wire __T_155_fromint__d;
    DFF_POSCLK #(.width(1)) _T_155_fromint (
        .q(__T_155_fromint__q),
        .d(__T_155_fromint__d),
        .clk(clock)
    );
    wire __T_155_toint__q;
    wire __T_155_toint__d;
    DFF_POSCLK #(.width(1)) _T_155_toint (
        .q(__T_155_toint__q),
        .d(__T_155_toint__d),
        .clk(clock)
    );
    wire __T_155_fastpipe__q;
    wire __T_155_fastpipe__d;
    DFF_POSCLK #(.width(1)) _T_155_fastpipe (
        .q(__T_155_fastpipe__q),
        .d(__T_155_fastpipe__d),
        .clk(clock)
    );
    wire __T_155_fma__q;
    wire __T_155_fma__d;
    DFF_POSCLK #(.width(1)) _T_155_fma (
        .q(__T_155_fma__q),
        .d(__T_155_fma__d),
        .clk(clock)
    );
    wire __T_155_div__q;
    wire __T_155_div__d;
    DFF_POSCLK #(.width(1)) _T_155_div (
        .q(__T_155_div__q),
        .d(__T_155_div__d),
        .clk(clock)
    );
    wire __T_155_sqrt__q;
    wire __T_155_sqrt__d;
    DFF_POSCLK #(.width(1)) _T_155_sqrt (
        .q(__T_155_sqrt__q),
        .d(__T_155_sqrt__d),
        .clk(clock)
    );
    wire __T_155_wflags__q;
    wire __T_155_wflags__d;
    DFF_POSCLK #(.width(1)) _T_155_wflags (
        .q(__T_155_wflags__q),
        .d(__T_155_wflags__d),
        .clk(clock)
    );
    wire [2:0] __T_155_rm__q;
    wire [2:0] __T_155_rm__d;
    DFF_POSCLK #(.width(3)) _T_155_rm (
        .q(__T_155_rm__q),
        .d(__T_155_rm__d),
        .clk(clock)
    );
    wire [1:0] __T_155_typ__q;
    wire [1:0] __T_155_typ__d;
    DFF_POSCLK #(.width(2)) _T_155_typ (
        .q(__T_155_typ__q),
        .d(__T_155_typ__d),
        .clk(clock)
    );
    wire [64:0] __T_155_in1__q;
    wire [64:0] __T_155_in1__d;
    DFF_POSCLK #(.width(65)) _T_155_in1 (
        .q(__T_155_in1__q),
        .d(__T_155_in1__d),
        .clk(clock)
    );
    wire [64:0] __T_155_in2__q;
    wire [64:0] __T_155_in2__d;
    DFF_POSCLK #(.width(65)) _T_155_in2 (
        .q(__T_155_in2__q),
        .d(__T_155_in2__d),
        .clk(clock)
    );
    wire [64:0] __T_155_in3__q;
    wire [64:0] __T_155_in3__d;
    DFF_POSCLK #(.width(65)) _T_155_in3 (
        .q(__T_155_in3__q),
        .d(__T_155_in3__d),
        .clk(clock)
    );
    wire in_valid;
    wire [4:0] in_bits_cmd;
    wire in_bits_ldst;
    wire in_bits_wen;
    wire in_bits_ren1;
    wire in_bits_ren2;
    wire in_bits_ren3;
    wire in_bits_swap12;
    wire in_bits_swap23;
    wire in_bits_single;
    wire in_bits_fromint;
    wire in_bits_toint;
    wire in_bits_fastpipe;
    wire in_bits_fma;
    wire in_bits_div;
    wire in_bits_sqrt;
    wire in_bits_wflags;
    wire [2:0] in_bits_rm;
    wire [1:0] in_bits_typ;
    wire [64:0] in_bits_in1;
    wire [64:0] in_bits_in2;
    wire [64:0] in_bits_in3;
    wire [64:0] mux_data;
    wire [4:0] mux_exc;
    wire _T_276;
    BITS #(.width(65), .high(31), .low(31)) bits_2147 (
        .y(_T_276),
        .in(in_bits_in1)
    );
    wire [7:0] _T_277;
    BITS #(.width(65), .high(30), .low(23)) bits_2148 (
        .y(_T_277),
        .in(in_bits_in1)
    );
    wire [22:0] _T_278;
    BITS #(.width(65), .high(22), .low(0)) bits_2149 (
        .y(_T_278),
        .in(in_bits_in1)
    );
    wire _T_280;
    wire [7:0] _WTEMP_277;
    PAD_UNSIGNED #(.width(1), .n(8)) u_pad_2150 (
        .y(_WTEMP_277),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(8)) u_eq_2151 (
        .y(_T_280),
        .a(_T_277),
        .b(_WTEMP_277)
    );
    wire _T_282;
    wire [22:0] _WTEMP_278;
    PAD_UNSIGNED #(.width(1), .n(23)) u_pad_2152 (
        .y(_WTEMP_278),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(23)) u_eq_2153 (
        .y(_T_282),
        .a(_T_278),
        .b(_WTEMP_278)
    );
    wire _T_283;
    BITWISEAND #(.width(1)) bitwiseand_2154 (
        .y(_T_283),
        .a(_T_280),
        .b(_T_282)
    );
    wire [31:0] _T_284;
    SHL_UNSIGNED #(.width(23), .n(9)) u_shl_2155 (
        .y(_T_284),
        .in(_T_278)
    );
    wire [15:0] _T_285;
    BITS #(.width(32), .high(31), .low(16)) bits_2156 (
        .y(_T_285),
        .in(_T_284)
    );
    wire [15:0] _T_286;
    BITS #(.width(32), .high(15), .low(0)) bits_2157 (
        .y(_T_286),
        .in(_T_284)
    );
    wire _T_288;
    wire [15:0] _WTEMP_279;
    PAD_UNSIGNED #(.width(1), .n(16)) u_pad_2158 (
        .y(_WTEMP_279),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(16)) u_neq_2159 (
        .y(_T_288),
        .a(_T_285),
        .b(_WTEMP_279)
    );
    wire [7:0] _T_289;
    BITS #(.width(16), .high(15), .low(8)) bits_2160 (
        .y(_T_289),
        .in(_T_285)
    );
    wire [7:0] _T_290;
    BITS #(.width(16), .high(7), .low(0)) bits_2161 (
        .y(_T_290),
        .in(_T_285)
    );
    wire _T_292;
    wire [7:0] _WTEMP_280;
    PAD_UNSIGNED #(.width(1), .n(8)) u_pad_2162 (
        .y(_WTEMP_280),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(8)) u_neq_2163 (
        .y(_T_292),
        .a(_T_289),
        .b(_WTEMP_280)
    );
    wire [3:0] _T_293;
    BITS #(.width(8), .high(7), .low(4)) bits_2164 (
        .y(_T_293),
        .in(_T_289)
    );
    wire [3:0] _T_294;
    BITS #(.width(8), .high(3), .low(0)) bits_2165 (
        .y(_T_294),
        .in(_T_289)
    );
    wire _T_296;
    wire [3:0] _WTEMP_281;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_2166 (
        .y(_WTEMP_281),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_2167 (
        .y(_T_296),
        .a(_T_293),
        .b(_WTEMP_281)
    );
    wire _T_297;
    BITS #(.width(4), .high(3), .low(3)) bits_2168 (
        .y(_T_297),
        .in(_T_293)
    );
    wire _T_299;
    BITS #(.width(4), .high(2), .low(2)) bits_2169 (
        .y(_T_299),
        .in(_T_293)
    );
    wire _T_301;
    BITS #(.width(4), .high(1), .low(1)) bits_2170 (
        .y(_T_301),
        .in(_T_293)
    );
    wire [1:0] _T_302;
    wire [1:0] _WTEMP_282;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2171 (
        .y(_WTEMP_282),
        .in(_T_301)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_2172 (
        .y(_T_302),
        .sel(_T_299),
        .a(2'h2),
        .b(_WTEMP_282)
    );
    wire [1:0] _T_303;
    MUX_UNSIGNED #(.width(2)) u_mux_2173 (
        .y(_T_303),
        .sel(_T_297),
        .a(2'h3),
        .b(_T_302)
    );
    wire _T_304;
    BITS #(.width(4), .high(3), .low(3)) bits_2174 (
        .y(_T_304),
        .in(_T_294)
    );
    wire _T_306;
    BITS #(.width(4), .high(2), .low(2)) bits_2175 (
        .y(_T_306),
        .in(_T_294)
    );
    wire _T_308;
    BITS #(.width(4), .high(1), .low(1)) bits_2176 (
        .y(_T_308),
        .in(_T_294)
    );
    wire [1:0] _T_309;
    wire [1:0] _WTEMP_283;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2177 (
        .y(_WTEMP_283),
        .in(_T_308)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_2178 (
        .y(_T_309),
        .sel(_T_306),
        .a(2'h2),
        .b(_WTEMP_283)
    );
    wire [1:0] _T_310;
    MUX_UNSIGNED #(.width(2)) u_mux_2179 (
        .y(_T_310),
        .sel(_T_304),
        .a(2'h3),
        .b(_T_309)
    );
    wire [1:0] _T_311;
    MUX_UNSIGNED #(.width(2)) u_mux_2180 (
        .y(_T_311),
        .sel(_T_296),
        .a(_T_303),
        .b(_T_310)
    );
    wire [2:0] _T_312;
    CAT #(.width_a(1), .width_b(2)) cat_2181 (
        .y(_T_312),
        .a(_T_296),
        .b(_T_311)
    );
    wire [3:0] _T_313;
    BITS #(.width(8), .high(7), .low(4)) bits_2182 (
        .y(_T_313),
        .in(_T_290)
    );
    wire [3:0] _T_314;
    BITS #(.width(8), .high(3), .low(0)) bits_2183 (
        .y(_T_314),
        .in(_T_290)
    );
    wire _T_316;
    wire [3:0] _WTEMP_284;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_2184 (
        .y(_WTEMP_284),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_2185 (
        .y(_T_316),
        .a(_T_313),
        .b(_WTEMP_284)
    );
    wire _T_317;
    BITS #(.width(4), .high(3), .low(3)) bits_2186 (
        .y(_T_317),
        .in(_T_313)
    );
    wire _T_319;
    BITS #(.width(4), .high(2), .low(2)) bits_2187 (
        .y(_T_319),
        .in(_T_313)
    );
    wire _T_321;
    BITS #(.width(4), .high(1), .low(1)) bits_2188 (
        .y(_T_321),
        .in(_T_313)
    );
    wire [1:0] _T_322;
    wire [1:0] _WTEMP_285;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2189 (
        .y(_WTEMP_285),
        .in(_T_321)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_2190 (
        .y(_T_322),
        .sel(_T_319),
        .a(2'h2),
        .b(_WTEMP_285)
    );
    wire [1:0] _T_323;
    MUX_UNSIGNED #(.width(2)) u_mux_2191 (
        .y(_T_323),
        .sel(_T_317),
        .a(2'h3),
        .b(_T_322)
    );
    wire _T_324;
    BITS #(.width(4), .high(3), .low(3)) bits_2192 (
        .y(_T_324),
        .in(_T_314)
    );
    wire _T_326;
    BITS #(.width(4), .high(2), .low(2)) bits_2193 (
        .y(_T_326),
        .in(_T_314)
    );
    wire _T_328;
    BITS #(.width(4), .high(1), .low(1)) bits_2194 (
        .y(_T_328),
        .in(_T_314)
    );
    wire [1:0] _T_329;
    wire [1:0] _WTEMP_286;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2195 (
        .y(_WTEMP_286),
        .in(_T_328)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_2196 (
        .y(_T_329),
        .sel(_T_326),
        .a(2'h2),
        .b(_WTEMP_286)
    );
    wire [1:0] _T_330;
    MUX_UNSIGNED #(.width(2)) u_mux_2197 (
        .y(_T_330),
        .sel(_T_324),
        .a(2'h3),
        .b(_T_329)
    );
    wire [1:0] _T_331;
    MUX_UNSIGNED #(.width(2)) u_mux_2198 (
        .y(_T_331),
        .sel(_T_316),
        .a(_T_323),
        .b(_T_330)
    );
    wire [2:0] _T_332;
    CAT #(.width_a(1), .width_b(2)) cat_2199 (
        .y(_T_332),
        .a(_T_316),
        .b(_T_331)
    );
    wire [2:0] _T_333;
    MUX_UNSIGNED #(.width(3)) u_mux_2200 (
        .y(_T_333),
        .sel(_T_292),
        .a(_T_312),
        .b(_T_332)
    );
    wire [3:0] _T_334;
    CAT #(.width_a(1), .width_b(3)) cat_2201 (
        .y(_T_334),
        .a(_T_292),
        .b(_T_333)
    );
    wire [7:0] _T_335;
    BITS #(.width(16), .high(15), .low(8)) bits_2202 (
        .y(_T_335),
        .in(_T_286)
    );
    wire [7:0] _T_336;
    BITS #(.width(16), .high(7), .low(0)) bits_2203 (
        .y(_T_336),
        .in(_T_286)
    );
    wire _T_338;
    wire [7:0] _WTEMP_287;
    PAD_UNSIGNED #(.width(1), .n(8)) u_pad_2204 (
        .y(_WTEMP_287),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(8)) u_neq_2205 (
        .y(_T_338),
        .a(_T_335),
        .b(_WTEMP_287)
    );
    wire [3:0] _T_339;
    BITS #(.width(8), .high(7), .low(4)) bits_2206 (
        .y(_T_339),
        .in(_T_335)
    );
    wire [3:0] _T_340;
    BITS #(.width(8), .high(3), .low(0)) bits_2207 (
        .y(_T_340),
        .in(_T_335)
    );
    wire _T_342;
    wire [3:0] _WTEMP_288;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_2208 (
        .y(_WTEMP_288),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_2209 (
        .y(_T_342),
        .a(_T_339),
        .b(_WTEMP_288)
    );
    wire _T_343;
    BITS #(.width(4), .high(3), .low(3)) bits_2210 (
        .y(_T_343),
        .in(_T_339)
    );
    wire _T_345;
    BITS #(.width(4), .high(2), .low(2)) bits_2211 (
        .y(_T_345),
        .in(_T_339)
    );
    wire _T_347;
    BITS #(.width(4), .high(1), .low(1)) bits_2212 (
        .y(_T_347),
        .in(_T_339)
    );
    wire [1:0] _T_348;
    wire [1:0] _WTEMP_289;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2213 (
        .y(_WTEMP_289),
        .in(_T_347)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_2214 (
        .y(_T_348),
        .sel(_T_345),
        .a(2'h2),
        .b(_WTEMP_289)
    );
    wire [1:0] _T_349;
    MUX_UNSIGNED #(.width(2)) u_mux_2215 (
        .y(_T_349),
        .sel(_T_343),
        .a(2'h3),
        .b(_T_348)
    );
    wire _T_350;
    BITS #(.width(4), .high(3), .low(3)) bits_2216 (
        .y(_T_350),
        .in(_T_340)
    );
    wire _T_352;
    BITS #(.width(4), .high(2), .low(2)) bits_2217 (
        .y(_T_352),
        .in(_T_340)
    );
    wire _T_354;
    BITS #(.width(4), .high(1), .low(1)) bits_2218 (
        .y(_T_354),
        .in(_T_340)
    );
    wire [1:0] _T_355;
    wire [1:0] _WTEMP_290;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2219 (
        .y(_WTEMP_290),
        .in(_T_354)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_2220 (
        .y(_T_355),
        .sel(_T_352),
        .a(2'h2),
        .b(_WTEMP_290)
    );
    wire [1:0] _T_356;
    MUX_UNSIGNED #(.width(2)) u_mux_2221 (
        .y(_T_356),
        .sel(_T_350),
        .a(2'h3),
        .b(_T_355)
    );
    wire [1:0] _T_357;
    MUX_UNSIGNED #(.width(2)) u_mux_2222 (
        .y(_T_357),
        .sel(_T_342),
        .a(_T_349),
        .b(_T_356)
    );
    wire [2:0] _T_358;
    CAT #(.width_a(1), .width_b(2)) cat_2223 (
        .y(_T_358),
        .a(_T_342),
        .b(_T_357)
    );
    wire [3:0] _T_359;
    BITS #(.width(8), .high(7), .low(4)) bits_2224 (
        .y(_T_359),
        .in(_T_336)
    );
    wire [3:0] _T_360;
    BITS #(.width(8), .high(3), .low(0)) bits_2225 (
        .y(_T_360),
        .in(_T_336)
    );
    wire _T_362;
    wire [3:0] _WTEMP_291;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_2226 (
        .y(_WTEMP_291),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_2227 (
        .y(_T_362),
        .a(_T_359),
        .b(_WTEMP_291)
    );
    wire _T_363;
    BITS #(.width(4), .high(3), .low(3)) bits_2228 (
        .y(_T_363),
        .in(_T_359)
    );
    wire _T_365;
    BITS #(.width(4), .high(2), .low(2)) bits_2229 (
        .y(_T_365),
        .in(_T_359)
    );
    wire _T_367;
    BITS #(.width(4), .high(1), .low(1)) bits_2230 (
        .y(_T_367),
        .in(_T_359)
    );
    wire [1:0] _T_368;
    wire [1:0] _WTEMP_292;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2231 (
        .y(_WTEMP_292),
        .in(_T_367)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_2232 (
        .y(_T_368),
        .sel(_T_365),
        .a(2'h2),
        .b(_WTEMP_292)
    );
    wire [1:0] _T_369;
    MUX_UNSIGNED #(.width(2)) u_mux_2233 (
        .y(_T_369),
        .sel(_T_363),
        .a(2'h3),
        .b(_T_368)
    );
    wire _T_370;
    BITS #(.width(4), .high(3), .low(3)) bits_2234 (
        .y(_T_370),
        .in(_T_360)
    );
    wire _T_372;
    BITS #(.width(4), .high(2), .low(2)) bits_2235 (
        .y(_T_372),
        .in(_T_360)
    );
    wire _T_374;
    BITS #(.width(4), .high(1), .low(1)) bits_2236 (
        .y(_T_374),
        .in(_T_360)
    );
    wire [1:0] _T_375;
    wire [1:0] _WTEMP_293;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2237 (
        .y(_WTEMP_293),
        .in(_T_374)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_2238 (
        .y(_T_375),
        .sel(_T_372),
        .a(2'h2),
        .b(_WTEMP_293)
    );
    wire [1:0] _T_376;
    MUX_UNSIGNED #(.width(2)) u_mux_2239 (
        .y(_T_376),
        .sel(_T_370),
        .a(2'h3),
        .b(_T_375)
    );
    wire [1:0] _T_377;
    MUX_UNSIGNED #(.width(2)) u_mux_2240 (
        .y(_T_377),
        .sel(_T_362),
        .a(_T_369),
        .b(_T_376)
    );
    wire [2:0] _T_378;
    CAT #(.width_a(1), .width_b(2)) cat_2241 (
        .y(_T_378),
        .a(_T_362),
        .b(_T_377)
    );
    wire [2:0] _T_379;
    MUX_UNSIGNED #(.width(3)) u_mux_2242 (
        .y(_T_379),
        .sel(_T_338),
        .a(_T_358),
        .b(_T_378)
    );
    wire [3:0] _T_380;
    CAT #(.width_a(1), .width_b(3)) cat_2243 (
        .y(_T_380),
        .a(_T_338),
        .b(_T_379)
    );
    wire [3:0] _T_381;
    MUX_UNSIGNED #(.width(4)) u_mux_2244 (
        .y(_T_381),
        .sel(_T_288),
        .a(_T_334),
        .b(_T_380)
    );
    wire [4:0] _T_382;
    CAT #(.width_a(1), .width_b(4)) cat_2245 (
        .y(_T_382),
        .a(_T_288),
        .b(_T_381)
    );
    wire [4:0] _T_383;
    BITWISENOT #(.width(5)) bitwisenot_2246 (
        .y(_T_383),
        .in(_T_382)
    );
    wire [53:0] _T_384;
    DSHL_UNSIGNED #(.width_in(23), .width_n(5)) u_dshl_2247 (
        .y(_T_384),
        .in(_T_278),
        .n(_T_383)
    );
    wire [21:0] _T_385;
    BITS #(.width(54), .high(21), .low(0)) bits_2248 (
        .y(_T_385),
        .in(_T_384)
    );
    wire [22:0] _T_387;
    CAT #(.width_a(22), .width_b(1)) cat_2249 (
        .y(_T_387),
        .a(_T_385),
        .b(1'h0)
    );
    wire [8:0] _T_392;
    assign _T_392 = 9'h1FF;
    wire [8:0] _T_393;
    wire [8:0] _WTEMP_294;
    PAD_UNSIGNED #(.width(5), .n(9)) u_pad_2250 (
        .y(_WTEMP_294),
        .in(_T_383)
    );
    BITWISEXOR #(.width(9)) bitwisexor_2251 (
        .y(_T_393),
        .a(_WTEMP_294),
        .b(_T_392)
    );
    wire [8:0] _T_394;
    wire [8:0] _WTEMP_295;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_2252 (
        .y(_WTEMP_295),
        .in(_T_277)
    );
    MUX_UNSIGNED #(.width(9)) u_mux_2253 (
        .y(_T_394),
        .sel(_T_280),
        .a(_T_393),
        .b(_WTEMP_295)
    );
    wire [1:0] _T_398;
    wire [1:0] _WTEMP_296;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2254 (
        .y(_WTEMP_296),
        .in(1'h1)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_2255 (
        .y(_T_398),
        .sel(_T_280),
        .a(2'h2),
        .b(_WTEMP_296)
    );
    wire [7:0] _T_399;
    wire [7:0] _WTEMP_297;
    PAD_UNSIGNED #(.width(2), .n(8)) u_pad_2256 (
        .y(_WTEMP_297),
        .in(_T_398)
    );
    BITWISEOR #(.width(8)) bitwiseor_2257 (
        .y(_T_399),
        .a(8'h80),
        .b(_WTEMP_297)
    );
    wire [9:0] _T_400;
    wire [8:0] _WTEMP_298;
    PAD_UNSIGNED #(.width(8), .n(9)) u_pad_2258 (
        .y(_WTEMP_298),
        .in(_T_399)
    );
    ADD_UNSIGNED #(.width(9)) u_add_2259 (
        .y(_T_400),
        .a(_T_394),
        .b(_WTEMP_298)
    );
    wire [8:0] _T_401;
    TAIL #(.width(10), .n(1)) tail_2260 (
        .y(_T_401),
        .in(_T_400)
    );
    wire [1:0] _T_402;
    BITS #(.width(9), .high(8), .low(7)) bits_2261 (
        .y(_T_402),
        .in(_T_401)
    );
    wire _T_404;
    EQ_UNSIGNED #(.width(2)) u_eq_2262 (
        .y(_T_404),
        .a(_T_402),
        .b(2'h3)
    );
    wire _T_406;
    EQ_UNSIGNED #(.width(1)) u_eq_2263 (
        .y(_T_406),
        .a(_T_282),
        .b(1'h0)
    );
    wire _T_407;
    BITWISEAND #(.width(1)) bitwiseand_2264 (
        .y(_T_407),
        .a(_T_404),
        .b(_T_406)
    );
    wire _T_408;
    BITS #(.width(1), .high(0), .low(0)) bits_2265 (
        .y(_T_408),
        .in(_T_283)
    );
    wire [2:0] _T_411;
    MUX_UNSIGNED #(.width(3)) u_mux_2266 (
        .y(_T_411),
        .sel(_T_408),
        .a(3'h7),
        .b(3'h0)
    );
    wire [8:0] _T_412;
    SHL_UNSIGNED #(.width(3), .n(6)) u_shl_2267 (
        .y(_T_412),
        .in(_T_411)
    );
    wire [8:0] _T_413;
    BITWISENOT #(.width(9)) bitwisenot_2268 (
        .y(_T_413),
        .in(_T_412)
    );
    wire [8:0] _T_414;
    BITWISEAND #(.width(9)) bitwiseand_2269 (
        .y(_T_414),
        .a(_T_401),
        .b(_T_413)
    );
    wire [6:0] _T_415;
    SHL_UNSIGNED #(.width(1), .n(6)) u_shl_2270 (
        .y(_T_415),
        .in(_T_407)
    );
    wire [8:0] _T_416;
    wire [8:0] _WTEMP_299;
    PAD_UNSIGNED #(.width(7), .n(9)) u_pad_2271 (
        .y(_WTEMP_299),
        .in(_T_415)
    );
    BITWISEOR #(.width(9)) bitwiseor_2272 (
        .y(_T_416),
        .a(_T_414),
        .b(_WTEMP_299)
    );
    wire [22:0] _T_417;
    MUX_UNSIGNED #(.width(23)) u_mux_2273 (
        .y(_T_417),
        .sel(_T_280),
        .a(_T_387),
        .b(_T_278)
    );
    wire [9:0] _T_418;
    CAT #(.width_a(1), .width_b(9)) cat_2274 (
        .y(_T_418),
        .a(_T_276),
        .b(_T_416)
    );
    wire [32:0] _T_419;
    CAT #(.width_a(10), .width_b(23)) cat_2275 (
        .y(_T_419),
        .a(_T_418),
        .b(_T_417)
    );
    wire _T_421;
    EQ_UNSIGNED #(.width(1)) u_eq_2276 (
        .y(_T_421),
        .a(in_bits_single),
        .b(1'h0)
    );
    wire _T_422;
    BITS #(.width(65), .high(63), .low(63)) bits_2277 (
        .y(_T_422),
        .in(in_bits_in1)
    );
    wire [10:0] _T_423;
    BITS #(.width(65), .high(62), .low(52)) bits_2278 (
        .y(_T_423),
        .in(in_bits_in1)
    );
    wire [51:0] _T_424;
    BITS #(.width(65), .high(51), .low(0)) bits_2279 (
        .y(_T_424),
        .in(in_bits_in1)
    );
    wire _T_426;
    wire [10:0] _WTEMP_300;
    PAD_UNSIGNED #(.width(1), .n(11)) u_pad_2280 (
        .y(_WTEMP_300),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(11)) u_eq_2281 (
        .y(_T_426),
        .a(_T_423),
        .b(_WTEMP_300)
    );
    wire _T_428;
    wire [51:0] _WTEMP_301;
    PAD_UNSIGNED #(.width(1), .n(52)) u_pad_2282 (
        .y(_WTEMP_301),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(52)) u_eq_2283 (
        .y(_T_428),
        .a(_T_424),
        .b(_WTEMP_301)
    );
    wire _T_429;
    BITWISEAND #(.width(1)) bitwiseand_2284 (
        .y(_T_429),
        .a(_T_426),
        .b(_T_428)
    );
    wire [63:0] _T_430;
    SHL_UNSIGNED #(.width(52), .n(12)) u_shl_2285 (
        .y(_T_430),
        .in(_T_424)
    );
    wire [31:0] _T_431;
    BITS #(.width(64), .high(63), .low(32)) bits_2286 (
        .y(_T_431),
        .in(_T_430)
    );
    wire [31:0] _T_432;
    BITS #(.width(64), .high(31), .low(0)) bits_2287 (
        .y(_T_432),
        .in(_T_430)
    );
    wire _T_434;
    wire [31:0] _WTEMP_302;
    PAD_UNSIGNED #(.width(1), .n(32)) u_pad_2288 (
        .y(_WTEMP_302),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(32)) u_neq_2289 (
        .y(_T_434),
        .a(_T_431),
        .b(_WTEMP_302)
    );
    wire [15:0] _T_435;
    BITS #(.width(32), .high(31), .low(16)) bits_2290 (
        .y(_T_435),
        .in(_T_431)
    );
    wire [15:0] _T_436;
    BITS #(.width(32), .high(15), .low(0)) bits_2291 (
        .y(_T_436),
        .in(_T_431)
    );
    wire _T_438;
    wire [15:0] _WTEMP_303;
    PAD_UNSIGNED #(.width(1), .n(16)) u_pad_2292 (
        .y(_WTEMP_303),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(16)) u_neq_2293 (
        .y(_T_438),
        .a(_T_435),
        .b(_WTEMP_303)
    );
    wire [7:0] _T_439;
    BITS #(.width(16), .high(15), .low(8)) bits_2294 (
        .y(_T_439),
        .in(_T_435)
    );
    wire [7:0] _T_440;
    BITS #(.width(16), .high(7), .low(0)) bits_2295 (
        .y(_T_440),
        .in(_T_435)
    );
    wire _T_442;
    wire [7:0] _WTEMP_304;
    PAD_UNSIGNED #(.width(1), .n(8)) u_pad_2296 (
        .y(_WTEMP_304),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(8)) u_neq_2297 (
        .y(_T_442),
        .a(_T_439),
        .b(_WTEMP_304)
    );
    wire [3:0] _T_443;
    BITS #(.width(8), .high(7), .low(4)) bits_2298 (
        .y(_T_443),
        .in(_T_439)
    );
    wire [3:0] _T_444;
    BITS #(.width(8), .high(3), .low(0)) bits_2299 (
        .y(_T_444),
        .in(_T_439)
    );
    wire _T_446;
    wire [3:0] _WTEMP_305;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_2300 (
        .y(_WTEMP_305),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_2301 (
        .y(_T_446),
        .a(_T_443),
        .b(_WTEMP_305)
    );
    wire _T_447;
    BITS #(.width(4), .high(3), .low(3)) bits_2302 (
        .y(_T_447),
        .in(_T_443)
    );
    wire _T_449;
    BITS #(.width(4), .high(2), .low(2)) bits_2303 (
        .y(_T_449),
        .in(_T_443)
    );
    wire _T_451;
    BITS #(.width(4), .high(1), .low(1)) bits_2304 (
        .y(_T_451),
        .in(_T_443)
    );
    wire [1:0] _T_452;
    wire [1:0] _WTEMP_306;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2305 (
        .y(_WTEMP_306),
        .in(_T_451)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_2306 (
        .y(_T_452),
        .sel(_T_449),
        .a(2'h2),
        .b(_WTEMP_306)
    );
    wire [1:0] _T_453;
    MUX_UNSIGNED #(.width(2)) u_mux_2307 (
        .y(_T_453),
        .sel(_T_447),
        .a(2'h3),
        .b(_T_452)
    );
    wire _T_454;
    BITS #(.width(4), .high(3), .low(3)) bits_2308 (
        .y(_T_454),
        .in(_T_444)
    );
    wire _T_456;
    BITS #(.width(4), .high(2), .low(2)) bits_2309 (
        .y(_T_456),
        .in(_T_444)
    );
    wire _T_458;
    BITS #(.width(4), .high(1), .low(1)) bits_2310 (
        .y(_T_458),
        .in(_T_444)
    );
    wire [1:0] _T_459;
    wire [1:0] _WTEMP_307;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2311 (
        .y(_WTEMP_307),
        .in(_T_458)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_2312 (
        .y(_T_459),
        .sel(_T_456),
        .a(2'h2),
        .b(_WTEMP_307)
    );
    wire [1:0] _T_460;
    MUX_UNSIGNED #(.width(2)) u_mux_2313 (
        .y(_T_460),
        .sel(_T_454),
        .a(2'h3),
        .b(_T_459)
    );
    wire [1:0] _T_461;
    MUX_UNSIGNED #(.width(2)) u_mux_2314 (
        .y(_T_461),
        .sel(_T_446),
        .a(_T_453),
        .b(_T_460)
    );
    wire [2:0] _T_462;
    CAT #(.width_a(1), .width_b(2)) cat_2315 (
        .y(_T_462),
        .a(_T_446),
        .b(_T_461)
    );
    wire [3:0] _T_463;
    BITS #(.width(8), .high(7), .low(4)) bits_2316 (
        .y(_T_463),
        .in(_T_440)
    );
    wire [3:0] _T_464;
    BITS #(.width(8), .high(3), .low(0)) bits_2317 (
        .y(_T_464),
        .in(_T_440)
    );
    wire _T_466;
    wire [3:0] _WTEMP_308;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_2318 (
        .y(_WTEMP_308),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_2319 (
        .y(_T_466),
        .a(_T_463),
        .b(_WTEMP_308)
    );
    wire _T_467;
    BITS #(.width(4), .high(3), .low(3)) bits_2320 (
        .y(_T_467),
        .in(_T_463)
    );
    wire _T_469;
    BITS #(.width(4), .high(2), .low(2)) bits_2321 (
        .y(_T_469),
        .in(_T_463)
    );
    wire _T_471;
    BITS #(.width(4), .high(1), .low(1)) bits_2322 (
        .y(_T_471),
        .in(_T_463)
    );
    wire [1:0] _T_472;
    wire [1:0] _WTEMP_309;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2323 (
        .y(_WTEMP_309),
        .in(_T_471)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_2324 (
        .y(_T_472),
        .sel(_T_469),
        .a(2'h2),
        .b(_WTEMP_309)
    );
    wire [1:0] _T_473;
    MUX_UNSIGNED #(.width(2)) u_mux_2325 (
        .y(_T_473),
        .sel(_T_467),
        .a(2'h3),
        .b(_T_472)
    );
    wire _T_474;
    BITS #(.width(4), .high(3), .low(3)) bits_2326 (
        .y(_T_474),
        .in(_T_464)
    );
    wire _T_476;
    BITS #(.width(4), .high(2), .low(2)) bits_2327 (
        .y(_T_476),
        .in(_T_464)
    );
    wire _T_478;
    BITS #(.width(4), .high(1), .low(1)) bits_2328 (
        .y(_T_478),
        .in(_T_464)
    );
    wire [1:0] _T_479;
    wire [1:0] _WTEMP_310;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2329 (
        .y(_WTEMP_310),
        .in(_T_478)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_2330 (
        .y(_T_479),
        .sel(_T_476),
        .a(2'h2),
        .b(_WTEMP_310)
    );
    wire [1:0] _T_480;
    MUX_UNSIGNED #(.width(2)) u_mux_2331 (
        .y(_T_480),
        .sel(_T_474),
        .a(2'h3),
        .b(_T_479)
    );
    wire [1:0] _T_481;
    MUX_UNSIGNED #(.width(2)) u_mux_2332 (
        .y(_T_481),
        .sel(_T_466),
        .a(_T_473),
        .b(_T_480)
    );
    wire [2:0] _T_482;
    CAT #(.width_a(1), .width_b(2)) cat_2333 (
        .y(_T_482),
        .a(_T_466),
        .b(_T_481)
    );
    wire [2:0] _T_483;
    MUX_UNSIGNED #(.width(3)) u_mux_2334 (
        .y(_T_483),
        .sel(_T_442),
        .a(_T_462),
        .b(_T_482)
    );
    wire [3:0] _T_484;
    CAT #(.width_a(1), .width_b(3)) cat_2335 (
        .y(_T_484),
        .a(_T_442),
        .b(_T_483)
    );
    wire [7:0] _T_485;
    BITS #(.width(16), .high(15), .low(8)) bits_2336 (
        .y(_T_485),
        .in(_T_436)
    );
    wire [7:0] _T_486;
    BITS #(.width(16), .high(7), .low(0)) bits_2337 (
        .y(_T_486),
        .in(_T_436)
    );
    wire _T_488;
    wire [7:0] _WTEMP_311;
    PAD_UNSIGNED #(.width(1), .n(8)) u_pad_2338 (
        .y(_WTEMP_311),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(8)) u_neq_2339 (
        .y(_T_488),
        .a(_T_485),
        .b(_WTEMP_311)
    );
    wire [3:0] _T_489;
    BITS #(.width(8), .high(7), .low(4)) bits_2340 (
        .y(_T_489),
        .in(_T_485)
    );
    wire [3:0] _T_490;
    BITS #(.width(8), .high(3), .low(0)) bits_2341 (
        .y(_T_490),
        .in(_T_485)
    );
    wire _T_492;
    wire [3:0] _WTEMP_312;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_2342 (
        .y(_WTEMP_312),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_2343 (
        .y(_T_492),
        .a(_T_489),
        .b(_WTEMP_312)
    );
    wire _T_493;
    BITS #(.width(4), .high(3), .low(3)) bits_2344 (
        .y(_T_493),
        .in(_T_489)
    );
    wire _T_495;
    BITS #(.width(4), .high(2), .low(2)) bits_2345 (
        .y(_T_495),
        .in(_T_489)
    );
    wire _T_497;
    BITS #(.width(4), .high(1), .low(1)) bits_2346 (
        .y(_T_497),
        .in(_T_489)
    );
    wire [1:0] _T_498;
    wire [1:0] _WTEMP_313;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2347 (
        .y(_WTEMP_313),
        .in(_T_497)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_2348 (
        .y(_T_498),
        .sel(_T_495),
        .a(2'h2),
        .b(_WTEMP_313)
    );
    wire [1:0] _T_499;
    MUX_UNSIGNED #(.width(2)) u_mux_2349 (
        .y(_T_499),
        .sel(_T_493),
        .a(2'h3),
        .b(_T_498)
    );
    wire _T_500;
    BITS #(.width(4), .high(3), .low(3)) bits_2350 (
        .y(_T_500),
        .in(_T_490)
    );
    wire _T_502;
    BITS #(.width(4), .high(2), .low(2)) bits_2351 (
        .y(_T_502),
        .in(_T_490)
    );
    wire _T_504;
    BITS #(.width(4), .high(1), .low(1)) bits_2352 (
        .y(_T_504),
        .in(_T_490)
    );
    wire [1:0] _T_505;
    wire [1:0] _WTEMP_314;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2353 (
        .y(_WTEMP_314),
        .in(_T_504)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_2354 (
        .y(_T_505),
        .sel(_T_502),
        .a(2'h2),
        .b(_WTEMP_314)
    );
    wire [1:0] _T_506;
    MUX_UNSIGNED #(.width(2)) u_mux_2355 (
        .y(_T_506),
        .sel(_T_500),
        .a(2'h3),
        .b(_T_505)
    );
    wire [1:0] _T_507;
    MUX_UNSIGNED #(.width(2)) u_mux_2356 (
        .y(_T_507),
        .sel(_T_492),
        .a(_T_499),
        .b(_T_506)
    );
    wire [2:0] _T_508;
    CAT #(.width_a(1), .width_b(2)) cat_2357 (
        .y(_T_508),
        .a(_T_492),
        .b(_T_507)
    );
    wire [3:0] _T_509;
    BITS #(.width(8), .high(7), .low(4)) bits_2358 (
        .y(_T_509),
        .in(_T_486)
    );
    wire [3:0] _T_510;
    BITS #(.width(8), .high(3), .low(0)) bits_2359 (
        .y(_T_510),
        .in(_T_486)
    );
    wire _T_512;
    wire [3:0] _WTEMP_315;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_2360 (
        .y(_WTEMP_315),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_2361 (
        .y(_T_512),
        .a(_T_509),
        .b(_WTEMP_315)
    );
    wire _T_513;
    BITS #(.width(4), .high(3), .low(3)) bits_2362 (
        .y(_T_513),
        .in(_T_509)
    );
    wire _T_515;
    BITS #(.width(4), .high(2), .low(2)) bits_2363 (
        .y(_T_515),
        .in(_T_509)
    );
    wire _T_517;
    BITS #(.width(4), .high(1), .low(1)) bits_2364 (
        .y(_T_517),
        .in(_T_509)
    );
    wire [1:0] _T_518;
    wire [1:0] _WTEMP_316;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2365 (
        .y(_WTEMP_316),
        .in(_T_517)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_2366 (
        .y(_T_518),
        .sel(_T_515),
        .a(2'h2),
        .b(_WTEMP_316)
    );
    wire [1:0] _T_519;
    MUX_UNSIGNED #(.width(2)) u_mux_2367 (
        .y(_T_519),
        .sel(_T_513),
        .a(2'h3),
        .b(_T_518)
    );
    wire _T_520;
    BITS #(.width(4), .high(3), .low(3)) bits_2368 (
        .y(_T_520),
        .in(_T_510)
    );
    wire _T_522;
    BITS #(.width(4), .high(2), .low(2)) bits_2369 (
        .y(_T_522),
        .in(_T_510)
    );
    wire _T_524;
    BITS #(.width(4), .high(1), .low(1)) bits_2370 (
        .y(_T_524),
        .in(_T_510)
    );
    wire [1:0] _T_525;
    wire [1:0] _WTEMP_317;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2371 (
        .y(_WTEMP_317),
        .in(_T_524)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_2372 (
        .y(_T_525),
        .sel(_T_522),
        .a(2'h2),
        .b(_WTEMP_317)
    );
    wire [1:0] _T_526;
    MUX_UNSIGNED #(.width(2)) u_mux_2373 (
        .y(_T_526),
        .sel(_T_520),
        .a(2'h3),
        .b(_T_525)
    );
    wire [1:0] _T_527;
    MUX_UNSIGNED #(.width(2)) u_mux_2374 (
        .y(_T_527),
        .sel(_T_512),
        .a(_T_519),
        .b(_T_526)
    );
    wire [2:0] _T_528;
    CAT #(.width_a(1), .width_b(2)) cat_2375 (
        .y(_T_528),
        .a(_T_512),
        .b(_T_527)
    );
    wire [2:0] _T_529;
    MUX_UNSIGNED #(.width(3)) u_mux_2376 (
        .y(_T_529),
        .sel(_T_488),
        .a(_T_508),
        .b(_T_528)
    );
    wire [3:0] _T_530;
    CAT #(.width_a(1), .width_b(3)) cat_2377 (
        .y(_T_530),
        .a(_T_488),
        .b(_T_529)
    );
    wire [3:0] _T_531;
    MUX_UNSIGNED #(.width(4)) u_mux_2378 (
        .y(_T_531),
        .sel(_T_438),
        .a(_T_484),
        .b(_T_530)
    );
    wire [4:0] _T_532;
    CAT #(.width_a(1), .width_b(4)) cat_2379 (
        .y(_T_532),
        .a(_T_438),
        .b(_T_531)
    );
    wire [15:0] _T_533;
    BITS #(.width(32), .high(31), .low(16)) bits_2380 (
        .y(_T_533),
        .in(_T_432)
    );
    wire [15:0] _T_534;
    BITS #(.width(32), .high(15), .low(0)) bits_2381 (
        .y(_T_534),
        .in(_T_432)
    );
    wire _T_536;
    wire [15:0] _WTEMP_318;
    PAD_UNSIGNED #(.width(1), .n(16)) u_pad_2382 (
        .y(_WTEMP_318),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(16)) u_neq_2383 (
        .y(_T_536),
        .a(_T_533),
        .b(_WTEMP_318)
    );
    wire [7:0] _T_537;
    BITS #(.width(16), .high(15), .low(8)) bits_2384 (
        .y(_T_537),
        .in(_T_533)
    );
    wire [7:0] _T_538;
    BITS #(.width(16), .high(7), .low(0)) bits_2385 (
        .y(_T_538),
        .in(_T_533)
    );
    wire _T_540;
    wire [7:0] _WTEMP_319;
    PAD_UNSIGNED #(.width(1), .n(8)) u_pad_2386 (
        .y(_WTEMP_319),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(8)) u_neq_2387 (
        .y(_T_540),
        .a(_T_537),
        .b(_WTEMP_319)
    );
    wire [3:0] _T_541;
    BITS #(.width(8), .high(7), .low(4)) bits_2388 (
        .y(_T_541),
        .in(_T_537)
    );
    wire [3:0] _T_542;
    BITS #(.width(8), .high(3), .low(0)) bits_2389 (
        .y(_T_542),
        .in(_T_537)
    );
    wire _T_544;
    wire [3:0] _WTEMP_320;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_2390 (
        .y(_WTEMP_320),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_2391 (
        .y(_T_544),
        .a(_T_541),
        .b(_WTEMP_320)
    );
    wire _T_545;
    BITS #(.width(4), .high(3), .low(3)) bits_2392 (
        .y(_T_545),
        .in(_T_541)
    );
    wire _T_547;
    BITS #(.width(4), .high(2), .low(2)) bits_2393 (
        .y(_T_547),
        .in(_T_541)
    );
    wire _T_549;
    BITS #(.width(4), .high(1), .low(1)) bits_2394 (
        .y(_T_549),
        .in(_T_541)
    );
    wire [1:0] _T_550;
    wire [1:0] _WTEMP_321;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2395 (
        .y(_WTEMP_321),
        .in(_T_549)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_2396 (
        .y(_T_550),
        .sel(_T_547),
        .a(2'h2),
        .b(_WTEMP_321)
    );
    wire [1:0] _T_551;
    MUX_UNSIGNED #(.width(2)) u_mux_2397 (
        .y(_T_551),
        .sel(_T_545),
        .a(2'h3),
        .b(_T_550)
    );
    wire _T_552;
    BITS #(.width(4), .high(3), .low(3)) bits_2398 (
        .y(_T_552),
        .in(_T_542)
    );
    wire _T_554;
    BITS #(.width(4), .high(2), .low(2)) bits_2399 (
        .y(_T_554),
        .in(_T_542)
    );
    wire _T_556;
    BITS #(.width(4), .high(1), .low(1)) bits_2400 (
        .y(_T_556),
        .in(_T_542)
    );
    wire [1:0] _T_557;
    wire [1:0] _WTEMP_322;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2401 (
        .y(_WTEMP_322),
        .in(_T_556)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_2402 (
        .y(_T_557),
        .sel(_T_554),
        .a(2'h2),
        .b(_WTEMP_322)
    );
    wire [1:0] _T_558;
    MUX_UNSIGNED #(.width(2)) u_mux_2403 (
        .y(_T_558),
        .sel(_T_552),
        .a(2'h3),
        .b(_T_557)
    );
    wire [1:0] _T_559;
    MUX_UNSIGNED #(.width(2)) u_mux_2404 (
        .y(_T_559),
        .sel(_T_544),
        .a(_T_551),
        .b(_T_558)
    );
    wire [2:0] _T_560;
    CAT #(.width_a(1), .width_b(2)) cat_2405 (
        .y(_T_560),
        .a(_T_544),
        .b(_T_559)
    );
    wire [3:0] _T_561;
    BITS #(.width(8), .high(7), .low(4)) bits_2406 (
        .y(_T_561),
        .in(_T_538)
    );
    wire [3:0] _T_562;
    BITS #(.width(8), .high(3), .low(0)) bits_2407 (
        .y(_T_562),
        .in(_T_538)
    );
    wire _T_564;
    wire [3:0] _WTEMP_323;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_2408 (
        .y(_WTEMP_323),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_2409 (
        .y(_T_564),
        .a(_T_561),
        .b(_WTEMP_323)
    );
    wire _T_565;
    BITS #(.width(4), .high(3), .low(3)) bits_2410 (
        .y(_T_565),
        .in(_T_561)
    );
    wire _T_567;
    BITS #(.width(4), .high(2), .low(2)) bits_2411 (
        .y(_T_567),
        .in(_T_561)
    );
    wire _T_569;
    BITS #(.width(4), .high(1), .low(1)) bits_2412 (
        .y(_T_569),
        .in(_T_561)
    );
    wire [1:0] _T_570;
    wire [1:0] _WTEMP_324;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2413 (
        .y(_WTEMP_324),
        .in(_T_569)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_2414 (
        .y(_T_570),
        .sel(_T_567),
        .a(2'h2),
        .b(_WTEMP_324)
    );
    wire [1:0] _T_571;
    MUX_UNSIGNED #(.width(2)) u_mux_2415 (
        .y(_T_571),
        .sel(_T_565),
        .a(2'h3),
        .b(_T_570)
    );
    wire _T_572;
    BITS #(.width(4), .high(3), .low(3)) bits_2416 (
        .y(_T_572),
        .in(_T_562)
    );
    wire _T_574;
    BITS #(.width(4), .high(2), .low(2)) bits_2417 (
        .y(_T_574),
        .in(_T_562)
    );
    wire _T_576;
    BITS #(.width(4), .high(1), .low(1)) bits_2418 (
        .y(_T_576),
        .in(_T_562)
    );
    wire [1:0] _T_577;
    wire [1:0] _WTEMP_325;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2419 (
        .y(_WTEMP_325),
        .in(_T_576)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_2420 (
        .y(_T_577),
        .sel(_T_574),
        .a(2'h2),
        .b(_WTEMP_325)
    );
    wire [1:0] _T_578;
    MUX_UNSIGNED #(.width(2)) u_mux_2421 (
        .y(_T_578),
        .sel(_T_572),
        .a(2'h3),
        .b(_T_577)
    );
    wire [1:0] _T_579;
    MUX_UNSIGNED #(.width(2)) u_mux_2422 (
        .y(_T_579),
        .sel(_T_564),
        .a(_T_571),
        .b(_T_578)
    );
    wire [2:0] _T_580;
    CAT #(.width_a(1), .width_b(2)) cat_2423 (
        .y(_T_580),
        .a(_T_564),
        .b(_T_579)
    );
    wire [2:0] _T_581;
    MUX_UNSIGNED #(.width(3)) u_mux_2424 (
        .y(_T_581),
        .sel(_T_540),
        .a(_T_560),
        .b(_T_580)
    );
    wire [3:0] _T_582;
    CAT #(.width_a(1), .width_b(3)) cat_2425 (
        .y(_T_582),
        .a(_T_540),
        .b(_T_581)
    );
    wire [7:0] _T_583;
    BITS #(.width(16), .high(15), .low(8)) bits_2426 (
        .y(_T_583),
        .in(_T_534)
    );
    wire [7:0] _T_584;
    BITS #(.width(16), .high(7), .low(0)) bits_2427 (
        .y(_T_584),
        .in(_T_534)
    );
    wire _T_586;
    wire [7:0] _WTEMP_326;
    PAD_UNSIGNED #(.width(1), .n(8)) u_pad_2428 (
        .y(_WTEMP_326),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(8)) u_neq_2429 (
        .y(_T_586),
        .a(_T_583),
        .b(_WTEMP_326)
    );
    wire [3:0] _T_587;
    BITS #(.width(8), .high(7), .low(4)) bits_2430 (
        .y(_T_587),
        .in(_T_583)
    );
    wire [3:0] _T_588;
    BITS #(.width(8), .high(3), .low(0)) bits_2431 (
        .y(_T_588),
        .in(_T_583)
    );
    wire _T_590;
    wire [3:0] _WTEMP_327;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_2432 (
        .y(_WTEMP_327),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_2433 (
        .y(_T_590),
        .a(_T_587),
        .b(_WTEMP_327)
    );
    wire _T_591;
    BITS #(.width(4), .high(3), .low(3)) bits_2434 (
        .y(_T_591),
        .in(_T_587)
    );
    wire _T_593;
    BITS #(.width(4), .high(2), .low(2)) bits_2435 (
        .y(_T_593),
        .in(_T_587)
    );
    wire _T_595;
    BITS #(.width(4), .high(1), .low(1)) bits_2436 (
        .y(_T_595),
        .in(_T_587)
    );
    wire [1:0] _T_596;
    wire [1:0] _WTEMP_328;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2437 (
        .y(_WTEMP_328),
        .in(_T_595)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_2438 (
        .y(_T_596),
        .sel(_T_593),
        .a(2'h2),
        .b(_WTEMP_328)
    );
    wire [1:0] _T_597;
    MUX_UNSIGNED #(.width(2)) u_mux_2439 (
        .y(_T_597),
        .sel(_T_591),
        .a(2'h3),
        .b(_T_596)
    );
    wire _T_598;
    BITS #(.width(4), .high(3), .low(3)) bits_2440 (
        .y(_T_598),
        .in(_T_588)
    );
    wire _T_600;
    BITS #(.width(4), .high(2), .low(2)) bits_2441 (
        .y(_T_600),
        .in(_T_588)
    );
    wire _T_602;
    BITS #(.width(4), .high(1), .low(1)) bits_2442 (
        .y(_T_602),
        .in(_T_588)
    );
    wire [1:0] _T_603;
    wire [1:0] _WTEMP_329;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2443 (
        .y(_WTEMP_329),
        .in(_T_602)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_2444 (
        .y(_T_603),
        .sel(_T_600),
        .a(2'h2),
        .b(_WTEMP_329)
    );
    wire [1:0] _T_604;
    MUX_UNSIGNED #(.width(2)) u_mux_2445 (
        .y(_T_604),
        .sel(_T_598),
        .a(2'h3),
        .b(_T_603)
    );
    wire [1:0] _T_605;
    MUX_UNSIGNED #(.width(2)) u_mux_2446 (
        .y(_T_605),
        .sel(_T_590),
        .a(_T_597),
        .b(_T_604)
    );
    wire [2:0] _T_606;
    CAT #(.width_a(1), .width_b(2)) cat_2447 (
        .y(_T_606),
        .a(_T_590),
        .b(_T_605)
    );
    wire [3:0] _T_607;
    BITS #(.width(8), .high(7), .low(4)) bits_2448 (
        .y(_T_607),
        .in(_T_584)
    );
    wire [3:0] _T_608;
    BITS #(.width(8), .high(3), .low(0)) bits_2449 (
        .y(_T_608),
        .in(_T_584)
    );
    wire _T_610;
    wire [3:0] _WTEMP_330;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_2450 (
        .y(_WTEMP_330),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_2451 (
        .y(_T_610),
        .a(_T_607),
        .b(_WTEMP_330)
    );
    wire _T_611;
    BITS #(.width(4), .high(3), .low(3)) bits_2452 (
        .y(_T_611),
        .in(_T_607)
    );
    wire _T_613;
    BITS #(.width(4), .high(2), .low(2)) bits_2453 (
        .y(_T_613),
        .in(_T_607)
    );
    wire _T_615;
    BITS #(.width(4), .high(1), .low(1)) bits_2454 (
        .y(_T_615),
        .in(_T_607)
    );
    wire [1:0] _T_616;
    wire [1:0] _WTEMP_331;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2455 (
        .y(_WTEMP_331),
        .in(_T_615)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_2456 (
        .y(_T_616),
        .sel(_T_613),
        .a(2'h2),
        .b(_WTEMP_331)
    );
    wire [1:0] _T_617;
    MUX_UNSIGNED #(.width(2)) u_mux_2457 (
        .y(_T_617),
        .sel(_T_611),
        .a(2'h3),
        .b(_T_616)
    );
    wire _T_618;
    BITS #(.width(4), .high(3), .low(3)) bits_2458 (
        .y(_T_618),
        .in(_T_608)
    );
    wire _T_620;
    BITS #(.width(4), .high(2), .low(2)) bits_2459 (
        .y(_T_620),
        .in(_T_608)
    );
    wire _T_622;
    BITS #(.width(4), .high(1), .low(1)) bits_2460 (
        .y(_T_622),
        .in(_T_608)
    );
    wire [1:0] _T_623;
    wire [1:0] _WTEMP_332;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2461 (
        .y(_WTEMP_332),
        .in(_T_622)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_2462 (
        .y(_T_623),
        .sel(_T_620),
        .a(2'h2),
        .b(_WTEMP_332)
    );
    wire [1:0] _T_624;
    MUX_UNSIGNED #(.width(2)) u_mux_2463 (
        .y(_T_624),
        .sel(_T_618),
        .a(2'h3),
        .b(_T_623)
    );
    wire [1:0] _T_625;
    MUX_UNSIGNED #(.width(2)) u_mux_2464 (
        .y(_T_625),
        .sel(_T_610),
        .a(_T_617),
        .b(_T_624)
    );
    wire [2:0] _T_626;
    CAT #(.width_a(1), .width_b(2)) cat_2465 (
        .y(_T_626),
        .a(_T_610),
        .b(_T_625)
    );
    wire [2:0] _T_627;
    MUX_UNSIGNED #(.width(3)) u_mux_2466 (
        .y(_T_627),
        .sel(_T_586),
        .a(_T_606),
        .b(_T_626)
    );
    wire [3:0] _T_628;
    CAT #(.width_a(1), .width_b(3)) cat_2467 (
        .y(_T_628),
        .a(_T_586),
        .b(_T_627)
    );
    wire [3:0] _T_629;
    MUX_UNSIGNED #(.width(4)) u_mux_2468 (
        .y(_T_629),
        .sel(_T_536),
        .a(_T_582),
        .b(_T_628)
    );
    wire [4:0] _T_630;
    CAT #(.width_a(1), .width_b(4)) cat_2469 (
        .y(_T_630),
        .a(_T_536),
        .b(_T_629)
    );
    wire [4:0] _T_631;
    MUX_UNSIGNED #(.width(5)) u_mux_2470 (
        .y(_T_631),
        .sel(_T_434),
        .a(_T_532),
        .b(_T_630)
    );
    wire [5:0] _T_632;
    CAT #(.width_a(1), .width_b(5)) cat_2471 (
        .y(_T_632),
        .a(_T_434),
        .b(_T_631)
    );
    wire [5:0] _T_633;
    BITWISENOT #(.width(6)) bitwisenot_2472 (
        .y(_T_633),
        .in(_T_632)
    );
    wire [114:0] _T_634;
    DSHL_UNSIGNED #(.width_in(52), .width_n(6)) u_dshl_2473 (
        .y(_T_634),
        .in(_T_424),
        .n(_T_633)
    );
    wire [50:0] _T_635;
    BITS #(.width(115), .high(50), .low(0)) bits_2474 (
        .y(_T_635),
        .in(_T_634)
    );
    wire [51:0] _T_637;
    CAT #(.width_a(51), .width_b(1)) cat_2475 (
        .y(_T_637),
        .a(_T_635),
        .b(1'h0)
    );
    wire [11:0] _T_642;
    assign _T_642 = 12'hFFF;
    wire [11:0] _T_643;
    wire [11:0] _WTEMP_333;
    PAD_UNSIGNED #(.width(6), .n(12)) u_pad_2476 (
        .y(_WTEMP_333),
        .in(_T_633)
    );
    BITWISEXOR #(.width(12)) bitwisexor_2477 (
        .y(_T_643),
        .a(_WTEMP_333),
        .b(_T_642)
    );
    wire [11:0] _T_644;
    wire [11:0] _WTEMP_334;
    PAD_UNSIGNED #(.width(11), .n(12)) u_pad_2478 (
        .y(_WTEMP_334),
        .in(_T_423)
    );
    MUX_UNSIGNED #(.width(12)) u_mux_2479 (
        .y(_T_644),
        .sel(_T_426),
        .a(_T_643),
        .b(_WTEMP_334)
    );
    wire [1:0] _T_648;
    wire [1:0] _WTEMP_335;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2480 (
        .y(_WTEMP_335),
        .in(1'h1)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_2481 (
        .y(_T_648),
        .sel(_T_426),
        .a(2'h2),
        .b(_WTEMP_335)
    );
    wire [10:0] _T_649;
    wire [10:0] _WTEMP_336;
    PAD_UNSIGNED #(.width(2), .n(11)) u_pad_2482 (
        .y(_WTEMP_336),
        .in(_T_648)
    );
    BITWISEOR #(.width(11)) bitwiseor_2483 (
        .y(_T_649),
        .a(11'h400),
        .b(_WTEMP_336)
    );
    wire [12:0] _T_650;
    wire [11:0] _WTEMP_337;
    PAD_UNSIGNED #(.width(11), .n(12)) u_pad_2484 (
        .y(_WTEMP_337),
        .in(_T_649)
    );
    ADD_UNSIGNED #(.width(12)) u_add_2485 (
        .y(_T_650),
        .a(_T_644),
        .b(_WTEMP_337)
    );
    wire [11:0] _T_651;
    TAIL #(.width(13), .n(1)) tail_2486 (
        .y(_T_651),
        .in(_T_650)
    );
    wire [1:0] _T_652;
    BITS #(.width(12), .high(11), .low(10)) bits_2487 (
        .y(_T_652),
        .in(_T_651)
    );
    wire _T_654;
    EQ_UNSIGNED #(.width(2)) u_eq_2488 (
        .y(_T_654),
        .a(_T_652),
        .b(2'h3)
    );
    wire _T_656;
    EQ_UNSIGNED #(.width(1)) u_eq_2489 (
        .y(_T_656),
        .a(_T_428),
        .b(1'h0)
    );
    wire _T_657;
    BITWISEAND #(.width(1)) bitwiseand_2490 (
        .y(_T_657),
        .a(_T_654),
        .b(_T_656)
    );
    wire _T_658;
    BITS #(.width(1), .high(0), .low(0)) bits_2491 (
        .y(_T_658),
        .in(_T_429)
    );
    wire [2:0] _T_661;
    MUX_UNSIGNED #(.width(3)) u_mux_2492 (
        .y(_T_661),
        .sel(_T_658),
        .a(3'h7),
        .b(3'h0)
    );
    wire [11:0] _T_662;
    SHL_UNSIGNED #(.width(3), .n(9)) u_shl_2493 (
        .y(_T_662),
        .in(_T_661)
    );
    wire [11:0] _T_663;
    BITWISENOT #(.width(12)) bitwisenot_2494 (
        .y(_T_663),
        .in(_T_662)
    );
    wire [11:0] _T_664;
    BITWISEAND #(.width(12)) bitwiseand_2495 (
        .y(_T_664),
        .a(_T_651),
        .b(_T_663)
    );
    wire [9:0] _T_665;
    SHL_UNSIGNED #(.width(1), .n(9)) u_shl_2496 (
        .y(_T_665),
        .in(_T_657)
    );
    wire [11:0] _T_666;
    wire [11:0] _WTEMP_338;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_2497 (
        .y(_WTEMP_338),
        .in(_T_665)
    );
    BITWISEOR #(.width(12)) bitwiseor_2498 (
        .y(_T_666),
        .a(_T_664),
        .b(_WTEMP_338)
    );
    wire [51:0] _T_667;
    MUX_UNSIGNED #(.width(52)) u_mux_2499 (
        .y(_T_667),
        .sel(_T_426),
        .a(_T_637),
        .b(_T_424)
    );
    wire [12:0] _T_668;
    CAT #(.width_a(1), .width_b(12)) cat_2500 (
        .y(_T_668),
        .a(_T_422),
        .b(_T_666)
    );
    wire [64:0] _T_669;
    CAT #(.width_a(13), .width_b(52)) cat_2501 (
        .y(_T_669),
        .a(_T_668),
        .b(_T_667)
    );
    wire [64:0] _T_670;
    ASSINT #(.width(65)) assint_2502 (
        .y(_T_670),
        .in(in_bits_in1)
    );
    wire [64:0] _T_671;
    wire [31:0] _T_672;
    BITS #(.width(65), .high(31), .low(0)) bits_2503 (
        .y(_T_672),
        .in(in_bits_in1)
    );
    wire _T_673;
    BITS #(.width(2), .high(1), .low(1)) bits_2504 (
        .y(_T_673),
        .in(in_bits_typ)
    );
    wire _T_675;
    EQ_UNSIGNED #(.width(1)) u_eq_2505 (
        .y(_T_675),
        .a(_T_673),
        .b(1'h0)
    );
    wire _T_676;
    BITS #(.width(2), .high(0), .low(0)) bits_2506 (
        .y(_T_676),
        .in(in_bits_typ)
    );
    wire [32:0] _T_677;
    CVT_UNSIGNED #(.width(32)) u_cvt_2507 (
        .y(_T_677),
        .in(_T_672)
    );
    wire [31:0] _T_678;
    ASSINT #(.width(32)) assint_2508 (
        .y(_T_678),
        .in(_T_672)
    );
    wire [32:0] _T_679;
    wire [32:0] _WTEMP_339;
    PAD_SIGNED #(.width(32), .n(33)) s_pad_2509 (
        .y(_WTEMP_339),
        .in(_T_678)
    );
    MUX_SIGNED #(.width(33)) s_mux_2510 (
        .y(_T_679),
        .sel(_T_676),
        .a(_T_677),
        .b(_WTEMP_339)
    );
    wire [64:0] intValue;
    ASUINT #(.width(65)) asuint_2511 (
        .y(intValue),
        .in(_T_671)
    );
    wire [4:0] _T_682;
    wire [4:0] _WTEMP_340;
    PAD_UNSIGNED #(.width(3), .n(5)) u_pad_2512 (
        .y(_WTEMP_340),
        .in(3'h4)
    );
    BITWISEAND #(.width(5)) bitwiseand_2513 (
        .y(_T_682),
        .a(in_bits_cmd),
        .b(_WTEMP_340)
    );
    wire _T_683;
    wire [4:0] _WTEMP_341;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_2514 (
        .y(_WTEMP_341),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(5)) u_eq_2515 (
        .y(_T_683),
        .a(_WTEMP_341),
        .b(_T_682)
    );
    wire _INToRecFN__clock;
    wire _INToRecFN__reset;
    wire _INToRecFN__io_signedIn;
    wire [63:0] _INToRecFN__io_in;
    wire [1:0] _INToRecFN__io_roundingMode;
    wire [32:0] _INToRecFN__io_out;
    wire [4:0] _INToRecFN__io_exceptionFlags;
    INToRecFN INToRecFN (
        .clock(_INToRecFN__clock),
        .reset(_INToRecFN__reset),
        .io_signedIn(_INToRecFN__io_signedIn),
        .io_in(_INToRecFN__io_in),
        .io_roundingMode(_INToRecFN__io_roundingMode),
        .io_out(_INToRecFN__io_out),
        .io_exceptionFlags(_INToRecFN__io_exceptionFlags)
    );
    wire _T_684;
    BITS #(.width(2), .high(0), .low(0)) bits_2763 (
        .y(_T_684),
        .in(in_bits_typ)
    );
    wire _T_685;
    BITWISENOT #(.width(1)) bitwisenot_2764 (
        .y(_T_685),
        .in(_T_684)
    );
    wire _INToRecFN_1__clock;
    wire _INToRecFN_1__reset;
    wire _INToRecFN_1__io_signedIn;
    wire [63:0] _INToRecFN_1__io_in;
    wire [1:0] _INToRecFN_1__io_roundingMode;
    wire [64:0] _INToRecFN_1__io_out;
    wire [4:0] _INToRecFN_1__io_exceptionFlags;
    INToRecFN_1 INToRecFN_1 (
        .clock(_INToRecFN_1__clock),
        .reset(_INToRecFN_1__reset),
        .io_signedIn(_INToRecFN_1__io_signedIn),
        .io_in(_INToRecFN_1__io_in),
        .io_roundingMode(_INToRecFN_1__io_roundingMode),
        .io_out(_INToRecFN_1__io_out),
        .io_exceptionFlags(_INToRecFN_1__io_exceptionFlags)
    );
    wire _T_686;
    BITS #(.width(2), .high(0), .low(0)) bits_3012 (
        .y(_T_686),
        .in(in_bits_typ)
    );
    wire _T_687;
    BITWISENOT #(.width(1)) bitwisenot_3013 (
        .y(_T_687),
        .in(_T_686)
    );
    wire [31:0] _T_688;
    SHR_UNSIGNED #(.width(65), .n(33)) u_shr_3014 (
        .y(_T_688),
        .in(_INToRecFN_1__io_out)
    );
    wire [64:0] _T_689;
    CAT #(.width_a(32), .width_b(33)) cat_3015 (
        .y(_T_689),
        .a(_T_688),
        .b(_INToRecFN__io_out)
    );
    wire _T_691;
    EQ_UNSIGNED #(.width(1)) u_eq_3016 (
        .y(_T_691),
        .a(in_bits_single),
        .b(1'h0)
    );
    wire [64:0] _node_27;
    MUX_UNSIGNED #(.width(65)) u_mux_3017 (
        .y(_node_27),
        .sel(_T_691),
        .a(_INToRecFN_1__io_out),
        .b(_T_689)
    );
    wire [64:0] _node_28;
    wire [64:0] _WTEMP_418;
    PAD_UNSIGNED #(.width(33), .n(65)) u_pad_3018 (
        .y(_WTEMP_418),
        .in(_T_419)
    );
    MUX_UNSIGNED #(.width(65)) u_mux_3019 (
        .y(_node_28),
        .sel(_T_421),
        .a(_T_669),
        .b(_WTEMP_418)
    );
    wire [4:0] _node_29;
    MUX_UNSIGNED #(.width(5)) u_mux_3020 (
        .y(_node_29),
        .sel(_T_691),
        .a(_INToRecFN_1__io_exceptionFlags),
        .b(_INToRecFN__io_exceptionFlags)
    );
    wire __T_694__q;
    wire __T_694__d;
    DFF_POSCLK #(.width(1)) _T_694 (
        .q(__T_694__q),
        .d(__T_694__d),
        .clk(clock)
    );
    wire _WTEMP_419;
    MUX_UNSIGNED #(.width(1)) u_mux_3021 (
        .y(__T_694__d),
        .sel(reset),
        .a(1'h0),
        .b(_WTEMP_419)
    );
    wire [64:0] __T_698_data__q;
    wire [64:0] __T_698_data__d;
    DFF_POSCLK #(.width(65)) _T_698_data (
        .q(__T_698_data__q),
        .d(__T_698_data__d),
        .clk(clock)
    );
    wire [4:0] __T_698_exc__q;
    wire [4:0] __T_698_exc__d;
    DFF_POSCLK #(.width(5)) _T_698_exc (
        .q(__T_698_exc__q),
        .d(__T_698_exc__d),
        .clk(clock)
    );
    wire _T_710_valid;
    wire [64:0] _T_710_bits_data;
    wire [4:0] _T_710_bits_exc;
    assign _INToRecFN__clock = clock;
    BITS #(.width(65), .high(63), .low(0)) bits_3022 (
        .y(_INToRecFN__io_in),
        .in(intValue)
    );
    BITS #(.width(3), .high(1), .low(0)) bits_3023 (
        .y(_INToRecFN__io_roundingMode),
        .in(in_bits_rm)
    );
    assign _INToRecFN__io_signedIn = _T_685;
    assign _INToRecFN__reset = reset;
    assign _INToRecFN_1__clock = clock;
    BITS #(.width(65), .high(63), .low(0)) bits_3024 (
        .y(_INToRecFN_1__io_in),
        .in(intValue)
    );
    BITS #(.width(3), .high(1), .low(0)) bits_3025 (
        .y(_INToRecFN_1__io_roundingMode),
        .in(in_bits_rm)
    );
    assign _INToRecFN_1__io_signedIn = _T_687;
    assign _INToRecFN_1__reset = reset;
    assign _WTEMP_276 = io_in_valid;
    MUX_UNSIGNED #(.width(5)) u_mux_3026 (
        .y(__T_155_cmd__d),
        .sel(io_in_valid),
        .a(io_in_bits_cmd),
        .b(__T_155_cmd__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_3027 (
        .y(__T_155_div__d),
        .sel(io_in_valid),
        .a(io_in_bits_div),
        .b(__T_155_div__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_3028 (
        .y(__T_155_fastpipe__d),
        .sel(io_in_valid),
        .a(io_in_bits_fastpipe),
        .b(__T_155_fastpipe__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_3029 (
        .y(__T_155_fma__d),
        .sel(io_in_valid),
        .a(io_in_bits_fma),
        .b(__T_155_fma__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_3030 (
        .y(__T_155_fromint__d),
        .sel(io_in_valid),
        .a(io_in_bits_fromint),
        .b(__T_155_fromint__q)
    );
    MUX_UNSIGNED #(.width(65)) u_mux_3031 (
        .y(__T_155_in1__d),
        .sel(io_in_valid),
        .a(io_in_bits_in1),
        .b(__T_155_in1__q)
    );
    MUX_UNSIGNED #(.width(65)) u_mux_3032 (
        .y(__T_155_in2__d),
        .sel(io_in_valid),
        .a(io_in_bits_in2),
        .b(__T_155_in2__q)
    );
    MUX_UNSIGNED #(.width(65)) u_mux_3033 (
        .y(__T_155_in3__d),
        .sel(io_in_valid),
        .a(io_in_bits_in3),
        .b(__T_155_in3__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_3034 (
        .y(__T_155_ldst__d),
        .sel(io_in_valid),
        .a(io_in_bits_ldst),
        .b(__T_155_ldst__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_3035 (
        .y(__T_155_ren1__d),
        .sel(io_in_valid),
        .a(io_in_bits_ren1),
        .b(__T_155_ren1__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_3036 (
        .y(__T_155_ren2__d),
        .sel(io_in_valid),
        .a(io_in_bits_ren2),
        .b(__T_155_ren2__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_3037 (
        .y(__T_155_ren3__d),
        .sel(io_in_valid),
        .a(io_in_bits_ren3),
        .b(__T_155_ren3__q)
    );
    MUX_UNSIGNED #(.width(3)) u_mux_3038 (
        .y(__T_155_rm__d),
        .sel(io_in_valid),
        .a(io_in_bits_rm),
        .b(__T_155_rm__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_3039 (
        .y(__T_155_single__d),
        .sel(io_in_valid),
        .a(io_in_bits_single),
        .b(__T_155_single__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_3040 (
        .y(__T_155_sqrt__d),
        .sel(io_in_valid),
        .a(io_in_bits_sqrt),
        .b(__T_155_sqrt__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_3041 (
        .y(__T_155_swap12__d),
        .sel(io_in_valid),
        .a(io_in_bits_swap12),
        .b(__T_155_swap12__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_3042 (
        .y(__T_155_swap23__d),
        .sel(io_in_valid),
        .a(io_in_bits_swap23),
        .b(__T_155_swap23__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_3043 (
        .y(__T_155_toint__d),
        .sel(io_in_valid),
        .a(io_in_bits_toint),
        .b(__T_155_toint__q)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_3044 (
        .y(__T_155_typ__d),
        .sel(io_in_valid),
        .a(io_in_bits_typ),
        .b(__T_155_typ__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_3045 (
        .y(__T_155_wen__d),
        .sel(io_in_valid),
        .a(io_in_bits_wen),
        .b(__T_155_wen__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_3046 (
        .y(__T_155_wflags__d),
        .sel(io_in_valid),
        .a(io_in_bits_wflags),
        .b(__T_155_wflags__q)
    );
    wire [64:0] _WTEMP_420;
    PAD_SIGNED #(.width(33), .n(65)) s_pad_3047 (
        .y(_WTEMP_420),
        .in(_T_679)
    );
    MUX_SIGNED #(.width(65)) s_mux_3048 (
        .y(_T_671),
        .sel(_T_675),
        .a(_WTEMP_420),
        .b(_T_670)
    );
    assign _WTEMP_419 = in_valid;
    MUX_UNSIGNED #(.width(65)) u_mux_3049 (
        .y(__T_698_data__d),
        .sel(in_valid),
        .a(mux_data),
        .b(__T_698_data__q)
    );
    MUX_UNSIGNED #(.width(5)) u_mux_3050 (
        .y(__T_698_exc__d),
        .sel(in_valid),
        .a(mux_exc),
        .b(__T_698_exc__q)
    );
    assign _T_710_bits_data = __T_698_data__q;
    assign _T_710_bits_exc = __T_698_exc__q;
    assign _T_710_valid = __T_694__q;
    assign in_bits_cmd = __T_155_cmd__q;
    assign in_bits_div = __T_155_div__q;
    assign in_bits_fastpipe = __T_155_fastpipe__q;
    assign in_bits_fma = __T_155_fma__q;
    assign in_bits_fromint = __T_155_fromint__q;
    assign in_bits_in1 = __T_155_in1__q;
    assign in_bits_in2 = __T_155_in2__q;
    assign in_bits_in3 = __T_155_in3__q;
    assign in_bits_ldst = __T_155_ldst__q;
    assign in_bits_ren1 = __T_155_ren1__q;
    assign in_bits_ren2 = __T_155_ren2__q;
    assign in_bits_ren3 = __T_155_ren3__q;
    assign in_bits_rm = __T_155_rm__q;
    assign in_bits_single = __T_155_single__q;
    assign in_bits_sqrt = __T_155_sqrt__q;
    assign in_bits_swap12 = __T_155_swap12__q;
    assign in_bits_swap23 = __T_155_swap23__q;
    assign in_bits_toint = __T_155_toint__q;
    assign in_bits_typ = __T_155_typ__q;
    assign in_bits_wen = __T_155_wen__q;
    assign in_bits_wflags = __T_155_wflags__q;
    assign in_valid = __T_132__q;
    assign io_out_bits_data = _T_710_bits_data;
    assign io_out_bits_exc = _T_710_bits_exc;
    assign io_out_valid = _T_710_valid;
    MUX_UNSIGNED #(.width(65)) u_mux_3051 (
        .y(mux_data),
        .sel(_T_683),
        .a(_node_27),
        .b(_node_28)
    );
    wire [4:0] _WTEMP_421;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_3052 (
        .y(_WTEMP_421),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(5)) u_mux_3053 (
        .y(mux_exc),
        .sel(_T_683),
        .a(_node_29),
        .b(_WTEMP_421)
    );
endmodule //IntToFP
module PAD_SIGNED(y, in);
    parameter width = 4;
    parameter n = 4;
    output [(n > width ? n : width)-1:0] y;
    input [width-1:0] in;
    assign y = n > width ? {{(n - width){in[width-1]}}, in} : in;
endmodule // PAD_SIGNED
module MUX_SIGNED(y, sel, a, b);
    parameter width = 4;
    output [width-1:0] y;
    input sel;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = sel ? $signed(a) : $signed(b);
endmodule // MUX_SIGNED
module INToRecFN(
    input clock,
    input reset,
    input io_signedIn,
    input [63:0] io_in,
    input [1:0] io_roundingMode,
    output [32:0] io_out,
    output [4:0] io_exceptionFlags
);
    wire _T_12;
    BITS #(.width(64), .high(63), .low(63)) bits_2516 (
        .y(_T_12),
        .in(io_in)
    );
    wire sign;
    BITWISEAND #(.width(1)) bitwiseand_2517 (
        .y(sign),
        .a(io_signedIn),
        .b(_T_12)
    );
    wire [64:0] _T_14;
    wire [63:0] _WTEMP_342;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_2518 (
        .y(_WTEMP_342),
        .in(1'h0)
    );
    SUB_UNSIGNED #(.width(64)) u_sub_2519 (
        .y(_T_14),
        .a(_WTEMP_342),
        .b(io_in)
    );
    wire [64:0] _T_15;
    ASUINT #(.width(65)) asuint_2520 (
        .y(_T_15),
        .in(_T_14)
    );
    wire [63:0] _T_16;
    TAIL #(.width(65), .n(1)) tail_2521 (
        .y(_T_16),
        .in(_T_15)
    );
    wire [63:0] absIn;
    MUX_UNSIGNED #(.width(64)) u_mux_2522 (
        .y(absIn),
        .sel(sign),
        .a(_T_16),
        .b(io_in)
    );
    wire [63:0] _T_17;
    SHL_UNSIGNED #(.width(64), .n(0)) u_shl_2523 (
        .y(_T_17),
        .in(absIn)
    );
    wire [31:0] _T_18;
    BITS #(.width(64), .high(63), .low(32)) bits_2524 (
        .y(_T_18),
        .in(_T_17)
    );
    wire [31:0] _T_19;
    BITS #(.width(64), .high(31), .low(0)) bits_2525 (
        .y(_T_19),
        .in(_T_17)
    );
    wire _T_21;
    wire [31:0] _WTEMP_343;
    PAD_UNSIGNED #(.width(1), .n(32)) u_pad_2526 (
        .y(_WTEMP_343),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(32)) u_neq_2527 (
        .y(_T_21),
        .a(_T_18),
        .b(_WTEMP_343)
    );
    wire [15:0] _T_22;
    BITS #(.width(32), .high(31), .low(16)) bits_2528 (
        .y(_T_22),
        .in(_T_18)
    );
    wire [15:0] _T_23;
    BITS #(.width(32), .high(15), .low(0)) bits_2529 (
        .y(_T_23),
        .in(_T_18)
    );
    wire _T_25;
    wire [15:0] _WTEMP_344;
    PAD_UNSIGNED #(.width(1), .n(16)) u_pad_2530 (
        .y(_WTEMP_344),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(16)) u_neq_2531 (
        .y(_T_25),
        .a(_T_22),
        .b(_WTEMP_344)
    );
    wire [7:0] _T_26;
    BITS #(.width(16), .high(15), .low(8)) bits_2532 (
        .y(_T_26),
        .in(_T_22)
    );
    wire [7:0] _T_27;
    BITS #(.width(16), .high(7), .low(0)) bits_2533 (
        .y(_T_27),
        .in(_T_22)
    );
    wire _T_29;
    wire [7:0] _WTEMP_345;
    PAD_UNSIGNED #(.width(1), .n(8)) u_pad_2534 (
        .y(_WTEMP_345),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(8)) u_neq_2535 (
        .y(_T_29),
        .a(_T_26),
        .b(_WTEMP_345)
    );
    wire [3:0] _T_30;
    BITS #(.width(8), .high(7), .low(4)) bits_2536 (
        .y(_T_30),
        .in(_T_26)
    );
    wire [3:0] _T_31;
    BITS #(.width(8), .high(3), .low(0)) bits_2537 (
        .y(_T_31),
        .in(_T_26)
    );
    wire _T_33;
    wire [3:0] _WTEMP_346;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_2538 (
        .y(_WTEMP_346),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_2539 (
        .y(_T_33),
        .a(_T_30),
        .b(_WTEMP_346)
    );
    wire _T_34;
    BITS #(.width(4), .high(3), .low(3)) bits_2540 (
        .y(_T_34),
        .in(_T_30)
    );
    wire _T_36;
    BITS #(.width(4), .high(2), .low(2)) bits_2541 (
        .y(_T_36),
        .in(_T_30)
    );
    wire _T_38;
    BITS #(.width(4), .high(1), .low(1)) bits_2542 (
        .y(_T_38),
        .in(_T_30)
    );
    wire [1:0] _T_39;
    wire [1:0] _WTEMP_347;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2543 (
        .y(_WTEMP_347),
        .in(_T_38)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_2544 (
        .y(_T_39),
        .sel(_T_36),
        .a(2'h2),
        .b(_WTEMP_347)
    );
    wire [1:0] _T_40;
    MUX_UNSIGNED #(.width(2)) u_mux_2545 (
        .y(_T_40),
        .sel(_T_34),
        .a(2'h3),
        .b(_T_39)
    );
    wire _T_41;
    BITS #(.width(4), .high(3), .low(3)) bits_2546 (
        .y(_T_41),
        .in(_T_31)
    );
    wire _T_43;
    BITS #(.width(4), .high(2), .low(2)) bits_2547 (
        .y(_T_43),
        .in(_T_31)
    );
    wire _T_45;
    BITS #(.width(4), .high(1), .low(1)) bits_2548 (
        .y(_T_45),
        .in(_T_31)
    );
    wire [1:0] _T_46;
    wire [1:0] _WTEMP_348;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2549 (
        .y(_WTEMP_348),
        .in(_T_45)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_2550 (
        .y(_T_46),
        .sel(_T_43),
        .a(2'h2),
        .b(_WTEMP_348)
    );
    wire [1:0] _T_47;
    MUX_UNSIGNED #(.width(2)) u_mux_2551 (
        .y(_T_47),
        .sel(_T_41),
        .a(2'h3),
        .b(_T_46)
    );
    wire [1:0] _T_48;
    MUX_UNSIGNED #(.width(2)) u_mux_2552 (
        .y(_T_48),
        .sel(_T_33),
        .a(_T_40),
        .b(_T_47)
    );
    wire [2:0] _T_49;
    CAT #(.width_a(1), .width_b(2)) cat_2553 (
        .y(_T_49),
        .a(_T_33),
        .b(_T_48)
    );
    wire [3:0] _T_50;
    BITS #(.width(8), .high(7), .low(4)) bits_2554 (
        .y(_T_50),
        .in(_T_27)
    );
    wire [3:0] _T_51;
    BITS #(.width(8), .high(3), .low(0)) bits_2555 (
        .y(_T_51),
        .in(_T_27)
    );
    wire _T_53;
    wire [3:0] _WTEMP_349;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_2556 (
        .y(_WTEMP_349),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_2557 (
        .y(_T_53),
        .a(_T_50),
        .b(_WTEMP_349)
    );
    wire _T_54;
    BITS #(.width(4), .high(3), .low(3)) bits_2558 (
        .y(_T_54),
        .in(_T_50)
    );
    wire _T_56;
    BITS #(.width(4), .high(2), .low(2)) bits_2559 (
        .y(_T_56),
        .in(_T_50)
    );
    wire _T_58;
    BITS #(.width(4), .high(1), .low(1)) bits_2560 (
        .y(_T_58),
        .in(_T_50)
    );
    wire [1:0] _T_59;
    wire [1:0] _WTEMP_350;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2561 (
        .y(_WTEMP_350),
        .in(_T_58)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_2562 (
        .y(_T_59),
        .sel(_T_56),
        .a(2'h2),
        .b(_WTEMP_350)
    );
    wire [1:0] _T_60;
    MUX_UNSIGNED #(.width(2)) u_mux_2563 (
        .y(_T_60),
        .sel(_T_54),
        .a(2'h3),
        .b(_T_59)
    );
    wire _T_61;
    BITS #(.width(4), .high(3), .low(3)) bits_2564 (
        .y(_T_61),
        .in(_T_51)
    );
    wire _T_63;
    BITS #(.width(4), .high(2), .low(2)) bits_2565 (
        .y(_T_63),
        .in(_T_51)
    );
    wire _T_65;
    BITS #(.width(4), .high(1), .low(1)) bits_2566 (
        .y(_T_65),
        .in(_T_51)
    );
    wire [1:0] _T_66;
    wire [1:0] _WTEMP_351;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2567 (
        .y(_WTEMP_351),
        .in(_T_65)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_2568 (
        .y(_T_66),
        .sel(_T_63),
        .a(2'h2),
        .b(_WTEMP_351)
    );
    wire [1:0] _T_67;
    MUX_UNSIGNED #(.width(2)) u_mux_2569 (
        .y(_T_67),
        .sel(_T_61),
        .a(2'h3),
        .b(_T_66)
    );
    wire [1:0] _T_68;
    MUX_UNSIGNED #(.width(2)) u_mux_2570 (
        .y(_T_68),
        .sel(_T_53),
        .a(_T_60),
        .b(_T_67)
    );
    wire [2:0] _T_69;
    CAT #(.width_a(1), .width_b(2)) cat_2571 (
        .y(_T_69),
        .a(_T_53),
        .b(_T_68)
    );
    wire [2:0] _T_70;
    MUX_UNSIGNED #(.width(3)) u_mux_2572 (
        .y(_T_70),
        .sel(_T_29),
        .a(_T_49),
        .b(_T_69)
    );
    wire [3:0] _T_71;
    CAT #(.width_a(1), .width_b(3)) cat_2573 (
        .y(_T_71),
        .a(_T_29),
        .b(_T_70)
    );
    wire [7:0] _T_72;
    BITS #(.width(16), .high(15), .low(8)) bits_2574 (
        .y(_T_72),
        .in(_T_23)
    );
    wire [7:0] _T_73;
    BITS #(.width(16), .high(7), .low(0)) bits_2575 (
        .y(_T_73),
        .in(_T_23)
    );
    wire _T_75;
    wire [7:0] _WTEMP_352;
    PAD_UNSIGNED #(.width(1), .n(8)) u_pad_2576 (
        .y(_WTEMP_352),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(8)) u_neq_2577 (
        .y(_T_75),
        .a(_T_72),
        .b(_WTEMP_352)
    );
    wire [3:0] _T_76;
    BITS #(.width(8), .high(7), .low(4)) bits_2578 (
        .y(_T_76),
        .in(_T_72)
    );
    wire [3:0] _T_77;
    BITS #(.width(8), .high(3), .low(0)) bits_2579 (
        .y(_T_77),
        .in(_T_72)
    );
    wire _T_79;
    wire [3:0] _WTEMP_353;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_2580 (
        .y(_WTEMP_353),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_2581 (
        .y(_T_79),
        .a(_T_76),
        .b(_WTEMP_353)
    );
    wire _T_80;
    BITS #(.width(4), .high(3), .low(3)) bits_2582 (
        .y(_T_80),
        .in(_T_76)
    );
    wire _T_82;
    BITS #(.width(4), .high(2), .low(2)) bits_2583 (
        .y(_T_82),
        .in(_T_76)
    );
    wire _T_84;
    BITS #(.width(4), .high(1), .low(1)) bits_2584 (
        .y(_T_84),
        .in(_T_76)
    );
    wire [1:0] _T_85;
    wire [1:0] _WTEMP_354;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2585 (
        .y(_WTEMP_354),
        .in(_T_84)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_2586 (
        .y(_T_85),
        .sel(_T_82),
        .a(2'h2),
        .b(_WTEMP_354)
    );
    wire [1:0] _T_86;
    MUX_UNSIGNED #(.width(2)) u_mux_2587 (
        .y(_T_86),
        .sel(_T_80),
        .a(2'h3),
        .b(_T_85)
    );
    wire _T_87;
    BITS #(.width(4), .high(3), .low(3)) bits_2588 (
        .y(_T_87),
        .in(_T_77)
    );
    wire _T_89;
    BITS #(.width(4), .high(2), .low(2)) bits_2589 (
        .y(_T_89),
        .in(_T_77)
    );
    wire _T_91;
    BITS #(.width(4), .high(1), .low(1)) bits_2590 (
        .y(_T_91),
        .in(_T_77)
    );
    wire [1:0] _T_92;
    wire [1:0] _WTEMP_355;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2591 (
        .y(_WTEMP_355),
        .in(_T_91)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_2592 (
        .y(_T_92),
        .sel(_T_89),
        .a(2'h2),
        .b(_WTEMP_355)
    );
    wire [1:0] _T_93;
    MUX_UNSIGNED #(.width(2)) u_mux_2593 (
        .y(_T_93),
        .sel(_T_87),
        .a(2'h3),
        .b(_T_92)
    );
    wire [1:0] _T_94;
    MUX_UNSIGNED #(.width(2)) u_mux_2594 (
        .y(_T_94),
        .sel(_T_79),
        .a(_T_86),
        .b(_T_93)
    );
    wire [2:0] _T_95;
    CAT #(.width_a(1), .width_b(2)) cat_2595 (
        .y(_T_95),
        .a(_T_79),
        .b(_T_94)
    );
    wire [3:0] _T_96;
    BITS #(.width(8), .high(7), .low(4)) bits_2596 (
        .y(_T_96),
        .in(_T_73)
    );
    wire [3:0] _T_97;
    BITS #(.width(8), .high(3), .low(0)) bits_2597 (
        .y(_T_97),
        .in(_T_73)
    );
    wire _T_99;
    wire [3:0] _WTEMP_356;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_2598 (
        .y(_WTEMP_356),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_2599 (
        .y(_T_99),
        .a(_T_96),
        .b(_WTEMP_356)
    );
    wire _T_100;
    BITS #(.width(4), .high(3), .low(3)) bits_2600 (
        .y(_T_100),
        .in(_T_96)
    );
    wire _T_102;
    BITS #(.width(4), .high(2), .low(2)) bits_2601 (
        .y(_T_102),
        .in(_T_96)
    );
    wire _T_104;
    BITS #(.width(4), .high(1), .low(1)) bits_2602 (
        .y(_T_104),
        .in(_T_96)
    );
    wire [1:0] _T_105;
    wire [1:0] _WTEMP_357;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2603 (
        .y(_WTEMP_357),
        .in(_T_104)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_2604 (
        .y(_T_105),
        .sel(_T_102),
        .a(2'h2),
        .b(_WTEMP_357)
    );
    wire [1:0] _T_106;
    MUX_UNSIGNED #(.width(2)) u_mux_2605 (
        .y(_T_106),
        .sel(_T_100),
        .a(2'h3),
        .b(_T_105)
    );
    wire _T_107;
    BITS #(.width(4), .high(3), .low(3)) bits_2606 (
        .y(_T_107),
        .in(_T_97)
    );
    wire _T_109;
    BITS #(.width(4), .high(2), .low(2)) bits_2607 (
        .y(_T_109),
        .in(_T_97)
    );
    wire _T_111;
    BITS #(.width(4), .high(1), .low(1)) bits_2608 (
        .y(_T_111),
        .in(_T_97)
    );
    wire [1:0] _T_112;
    wire [1:0] _WTEMP_358;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2609 (
        .y(_WTEMP_358),
        .in(_T_111)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_2610 (
        .y(_T_112),
        .sel(_T_109),
        .a(2'h2),
        .b(_WTEMP_358)
    );
    wire [1:0] _T_113;
    MUX_UNSIGNED #(.width(2)) u_mux_2611 (
        .y(_T_113),
        .sel(_T_107),
        .a(2'h3),
        .b(_T_112)
    );
    wire [1:0] _T_114;
    MUX_UNSIGNED #(.width(2)) u_mux_2612 (
        .y(_T_114),
        .sel(_T_99),
        .a(_T_106),
        .b(_T_113)
    );
    wire [2:0] _T_115;
    CAT #(.width_a(1), .width_b(2)) cat_2613 (
        .y(_T_115),
        .a(_T_99),
        .b(_T_114)
    );
    wire [2:0] _T_116;
    MUX_UNSIGNED #(.width(3)) u_mux_2614 (
        .y(_T_116),
        .sel(_T_75),
        .a(_T_95),
        .b(_T_115)
    );
    wire [3:0] _T_117;
    CAT #(.width_a(1), .width_b(3)) cat_2615 (
        .y(_T_117),
        .a(_T_75),
        .b(_T_116)
    );
    wire [3:0] _T_118;
    MUX_UNSIGNED #(.width(4)) u_mux_2616 (
        .y(_T_118),
        .sel(_T_25),
        .a(_T_71),
        .b(_T_117)
    );
    wire [4:0] _T_119;
    CAT #(.width_a(1), .width_b(4)) cat_2617 (
        .y(_T_119),
        .a(_T_25),
        .b(_T_118)
    );
    wire [15:0] _T_120;
    BITS #(.width(32), .high(31), .low(16)) bits_2618 (
        .y(_T_120),
        .in(_T_19)
    );
    wire [15:0] _T_121;
    BITS #(.width(32), .high(15), .low(0)) bits_2619 (
        .y(_T_121),
        .in(_T_19)
    );
    wire _T_123;
    wire [15:0] _WTEMP_359;
    PAD_UNSIGNED #(.width(1), .n(16)) u_pad_2620 (
        .y(_WTEMP_359),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(16)) u_neq_2621 (
        .y(_T_123),
        .a(_T_120),
        .b(_WTEMP_359)
    );
    wire [7:0] _T_124;
    BITS #(.width(16), .high(15), .low(8)) bits_2622 (
        .y(_T_124),
        .in(_T_120)
    );
    wire [7:0] _T_125;
    BITS #(.width(16), .high(7), .low(0)) bits_2623 (
        .y(_T_125),
        .in(_T_120)
    );
    wire _T_127;
    wire [7:0] _WTEMP_360;
    PAD_UNSIGNED #(.width(1), .n(8)) u_pad_2624 (
        .y(_WTEMP_360),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(8)) u_neq_2625 (
        .y(_T_127),
        .a(_T_124),
        .b(_WTEMP_360)
    );
    wire [3:0] _T_128;
    BITS #(.width(8), .high(7), .low(4)) bits_2626 (
        .y(_T_128),
        .in(_T_124)
    );
    wire [3:0] _T_129;
    BITS #(.width(8), .high(3), .low(0)) bits_2627 (
        .y(_T_129),
        .in(_T_124)
    );
    wire _T_131;
    wire [3:0] _WTEMP_361;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_2628 (
        .y(_WTEMP_361),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_2629 (
        .y(_T_131),
        .a(_T_128),
        .b(_WTEMP_361)
    );
    wire _T_132;
    BITS #(.width(4), .high(3), .low(3)) bits_2630 (
        .y(_T_132),
        .in(_T_128)
    );
    wire _T_134;
    BITS #(.width(4), .high(2), .low(2)) bits_2631 (
        .y(_T_134),
        .in(_T_128)
    );
    wire _T_136;
    BITS #(.width(4), .high(1), .low(1)) bits_2632 (
        .y(_T_136),
        .in(_T_128)
    );
    wire [1:0] _T_137;
    wire [1:0] _WTEMP_362;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2633 (
        .y(_WTEMP_362),
        .in(_T_136)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_2634 (
        .y(_T_137),
        .sel(_T_134),
        .a(2'h2),
        .b(_WTEMP_362)
    );
    wire [1:0] _T_138;
    MUX_UNSIGNED #(.width(2)) u_mux_2635 (
        .y(_T_138),
        .sel(_T_132),
        .a(2'h3),
        .b(_T_137)
    );
    wire _T_139;
    BITS #(.width(4), .high(3), .low(3)) bits_2636 (
        .y(_T_139),
        .in(_T_129)
    );
    wire _T_141;
    BITS #(.width(4), .high(2), .low(2)) bits_2637 (
        .y(_T_141),
        .in(_T_129)
    );
    wire _T_143;
    BITS #(.width(4), .high(1), .low(1)) bits_2638 (
        .y(_T_143),
        .in(_T_129)
    );
    wire [1:0] _T_144;
    wire [1:0] _WTEMP_363;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2639 (
        .y(_WTEMP_363),
        .in(_T_143)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_2640 (
        .y(_T_144),
        .sel(_T_141),
        .a(2'h2),
        .b(_WTEMP_363)
    );
    wire [1:0] _T_145;
    MUX_UNSIGNED #(.width(2)) u_mux_2641 (
        .y(_T_145),
        .sel(_T_139),
        .a(2'h3),
        .b(_T_144)
    );
    wire [1:0] _T_146;
    MUX_UNSIGNED #(.width(2)) u_mux_2642 (
        .y(_T_146),
        .sel(_T_131),
        .a(_T_138),
        .b(_T_145)
    );
    wire [2:0] _T_147;
    CAT #(.width_a(1), .width_b(2)) cat_2643 (
        .y(_T_147),
        .a(_T_131),
        .b(_T_146)
    );
    wire [3:0] _T_148;
    BITS #(.width(8), .high(7), .low(4)) bits_2644 (
        .y(_T_148),
        .in(_T_125)
    );
    wire [3:0] _T_149;
    BITS #(.width(8), .high(3), .low(0)) bits_2645 (
        .y(_T_149),
        .in(_T_125)
    );
    wire _T_151;
    wire [3:0] _WTEMP_364;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_2646 (
        .y(_WTEMP_364),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_2647 (
        .y(_T_151),
        .a(_T_148),
        .b(_WTEMP_364)
    );
    wire _T_152;
    BITS #(.width(4), .high(3), .low(3)) bits_2648 (
        .y(_T_152),
        .in(_T_148)
    );
    wire _T_154;
    BITS #(.width(4), .high(2), .low(2)) bits_2649 (
        .y(_T_154),
        .in(_T_148)
    );
    wire _T_156;
    BITS #(.width(4), .high(1), .low(1)) bits_2650 (
        .y(_T_156),
        .in(_T_148)
    );
    wire [1:0] _T_157;
    wire [1:0] _WTEMP_365;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2651 (
        .y(_WTEMP_365),
        .in(_T_156)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_2652 (
        .y(_T_157),
        .sel(_T_154),
        .a(2'h2),
        .b(_WTEMP_365)
    );
    wire [1:0] _T_158;
    MUX_UNSIGNED #(.width(2)) u_mux_2653 (
        .y(_T_158),
        .sel(_T_152),
        .a(2'h3),
        .b(_T_157)
    );
    wire _T_159;
    BITS #(.width(4), .high(3), .low(3)) bits_2654 (
        .y(_T_159),
        .in(_T_149)
    );
    wire _T_161;
    BITS #(.width(4), .high(2), .low(2)) bits_2655 (
        .y(_T_161),
        .in(_T_149)
    );
    wire _T_163;
    BITS #(.width(4), .high(1), .low(1)) bits_2656 (
        .y(_T_163),
        .in(_T_149)
    );
    wire [1:0] _T_164;
    wire [1:0] _WTEMP_366;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2657 (
        .y(_WTEMP_366),
        .in(_T_163)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_2658 (
        .y(_T_164),
        .sel(_T_161),
        .a(2'h2),
        .b(_WTEMP_366)
    );
    wire [1:0] _T_165;
    MUX_UNSIGNED #(.width(2)) u_mux_2659 (
        .y(_T_165),
        .sel(_T_159),
        .a(2'h3),
        .b(_T_164)
    );
    wire [1:0] _T_166;
    MUX_UNSIGNED #(.width(2)) u_mux_2660 (
        .y(_T_166),
        .sel(_T_151),
        .a(_T_158),
        .b(_T_165)
    );
    wire [2:0] _T_167;
    CAT #(.width_a(1), .width_b(2)) cat_2661 (
        .y(_T_167),
        .a(_T_151),
        .b(_T_166)
    );
    wire [2:0] _T_168;
    MUX_UNSIGNED #(.width(3)) u_mux_2662 (
        .y(_T_168),
        .sel(_T_127),
        .a(_T_147),
        .b(_T_167)
    );
    wire [3:0] _T_169;
    CAT #(.width_a(1), .width_b(3)) cat_2663 (
        .y(_T_169),
        .a(_T_127),
        .b(_T_168)
    );
    wire [7:0] _T_170;
    BITS #(.width(16), .high(15), .low(8)) bits_2664 (
        .y(_T_170),
        .in(_T_121)
    );
    wire [7:0] _T_171;
    BITS #(.width(16), .high(7), .low(0)) bits_2665 (
        .y(_T_171),
        .in(_T_121)
    );
    wire _T_173;
    wire [7:0] _WTEMP_367;
    PAD_UNSIGNED #(.width(1), .n(8)) u_pad_2666 (
        .y(_WTEMP_367),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(8)) u_neq_2667 (
        .y(_T_173),
        .a(_T_170),
        .b(_WTEMP_367)
    );
    wire [3:0] _T_174;
    BITS #(.width(8), .high(7), .low(4)) bits_2668 (
        .y(_T_174),
        .in(_T_170)
    );
    wire [3:0] _T_175;
    BITS #(.width(8), .high(3), .low(0)) bits_2669 (
        .y(_T_175),
        .in(_T_170)
    );
    wire _T_177;
    wire [3:0] _WTEMP_368;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_2670 (
        .y(_WTEMP_368),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_2671 (
        .y(_T_177),
        .a(_T_174),
        .b(_WTEMP_368)
    );
    wire _T_178;
    BITS #(.width(4), .high(3), .low(3)) bits_2672 (
        .y(_T_178),
        .in(_T_174)
    );
    wire _T_180;
    BITS #(.width(4), .high(2), .low(2)) bits_2673 (
        .y(_T_180),
        .in(_T_174)
    );
    wire _T_182;
    BITS #(.width(4), .high(1), .low(1)) bits_2674 (
        .y(_T_182),
        .in(_T_174)
    );
    wire [1:0] _T_183;
    wire [1:0] _WTEMP_369;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2675 (
        .y(_WTEMP_369),
        .in(_T_182)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_2676 (
        .y(_T_183),
        .sel(_T_180),
        .a(2'h2),
        .b(_WTEMP_369)
    );
    wire [1:0] _T_184;
    MUX_UNSIGNED #(.width(2)) u_mux_2677 (
        .y(_T_184),
        .sel(_T_178),
        .a(2'h3),
        .b(_T_183)
    );
    wire _T_185;
    BITS #(.width(4), .high(3), .low(3)) bits_2678 (
        .y(_T_185),
        .in(_T_175)
    );
    wire _T_187;
    BITS #(.width(4), .high(2), .low(2)) bits_2679 (
        .y(_T_187),
        .in(_T_175)
    );
    wire _T_189;
    BITS #(.width(4), .high(1), .low(1)) bits_2680 (
        .y(_T_189),
        .in(_T_175)
    );
    wire [1:0] _T_190;
    wire [1:0] _WTEMP_370;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2681 (
        .y(_WTEMP_370),
        .in(_T_189)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_2682 (
        .y(_T_190),
        .sel(_T_187),
        .a(2'h2),
        .b(_WTEMP_370)
    );
    wire [1:0] _T_191;
    MUX_UNSIGNED #(.width(2)) u_mux_2683 (
        .y(_T_191),
        .sel(_T_185),
        .a(2'h3),
        .b(_T_190)
    );
    wire [1:0] _T_192;
    MUX_UNSIGNED #(.width(2)) u_mux_2684 (
        .y(_T_192),
        .sel(_T_177),
        .a(_T_184),
        .b(_T_191)
    );
    wire [2:0] _T_193;
    CAT #(.width_a(1), .width_b(2)) cat_2685 (
        .y(_T_193),
        .a(_T_177),
        .b(_T_192)
    );
    wire [3:0] _T_194;
    BITS #(.width(8), .high(7), .low(4)) bits_2686 (
        .y(_T_194),
        .in(_T_171)
    );
    wire [3:0] _T_195;
    BITS #(.width(8), .high(3), .low(0)) bits_2687 (
        .y(_T_195),
        .in(_T_171)
    );
    wire _T_197;
    wire [3:0] _WTEMP_371;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_2688 (
        .y(_WTEMP_371),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_2689 (
        .y(_T_197),
        .a(_T_194),
        .b(_WTEMP_371)
    );
    wire _T_198;
    BITS #(.width(4), .high(3), .low(3)) bits_2690 (
        .y(_T_198),
        .in(_T_194)
    );
    wire _T_200;
    BITS #(.width(4), .high(2), .low(2)) bits_2691 (
        .y(_T_200),
        .in(_T_194)
    );
    wire _T_202;
    BITS #(.width(4), .high(1), .low(1)) bits_2692 (
        .y(_T_202),
        .in(_T_194)
    );
    wire [1:0] _T_203;
    wire [1:0] _WTEMP_372;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2693 (
        .y(_WTEMP_372),
        .in(_T_202)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_2694 (
        .y(_T_203),
        .sel(_T_200),
        .a(2'h2),
        .b(_WTEMP_372)
    );
    wire [1:0] _T_204;
    MUX_UNSIGNED #(.width(2)) u_mux_2695 (
        .y(_T_204),
        .sel(_T_198),
        .a(2'h3),
        .b(_T_203)
    );
    wire _T_205;
    BITS #(.width(4), .high(3), .low(3)) bits_2696 (
        .y(_T_205),
        .in(_T_195)
    );
    wire _T_207;
    BITS #(.width(4), .high(2), .low(2)) bits_2697 (
        .y(_T_207),
        .in(_T_195)
    );
    wire _T_209;
    BITS #(.width(4), .high(1), .low(1)) bits_2698 (
        .y(_T_209),
        .in(_T_195)
    );
    wire [1:0] _T_210;
    wire [1:0] _WTEMP_373;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2699 (
        .y(_WTEMP_373),
        .in(_T_209)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_2700 (
        .y(_T_210),
        .sel(_T_207),
        .a(2'h2),
        .b(_WTEMP_373)
    );
    wire [1:0] _T_211;
    MUX_UNSIGNED #(.width(2)) u_mux_2701 (
        .y(_T_211),
        .sel(_T_205),
        .a(2'h3),
        .b(_T_210)
    );
    wire [1:0] _T_212;
    MUX_UNSIGNED #(.width(2)) u_mux_2702 (
        .y(_T_212),
        .sel(_T_197),
        .a(_T_204),
        .b(_T_211)
    );
    wire [2:0] _T_213;
    CAT #(.width_a(1), .width_b(2)) cat_2703 (
        .y(_T_213),
        .a(_T_197),
        .b(_T_212)
    );
    wire [2:0] _T_214;
    MUX_UNSIGNED #(.width(3)) u_mux_2704 (
        .y(_T_214),
        .sel(_T_173),
        .a(_T_193),
        .b(_T_213)
    );
    wire [3:0] _T_215;
    CAT #(.width_a(1), .width_b(3)) cat_2705 (
        .y(_T_215),
        .a(_T_173),
        .b(_T_214)
    );
    wire [3:0] _T_216;
    MUX_UNSIGNED #(.width(4)) u_mux_2706 (
        .y(_T_216),
        .sel(_T_123),
        .a(_T_169),
        .b(_T_215)
    );
    wire [4:0] _T_217;
    CAT #(.width_a(1), .width_b(4)) cat_2707 (
        .y(_T_217),
        .a(_T_123),
        .b(_T_216)
    );
    wire [4:0] _T_218;
    MUX_UNSIGNED #(.width(5)) u_mux_2708 (
        .y(_T_218),
        .sel(_T_21),
        .a(_T_119),
        .b(_T_217)
    );
    wire [5:0] _T_219;
    CAT #(.width_a(1), .width_b(5)) cat_2709 (
        .y(_T_219),
        .a(_T_21),
        .b(_T_218)
    );
    wire [5:0] normCount;
    BITWISENOT #(.width(6)) bitwisenot_2710 (
        .y(normCount),
        .in(_T_219)
    );
    wire [126:0] _T_220;
    DSHL_UNSIGNED #(.width_in(64), .width_n(6)) u_dshl_2711 (
        .y(_T_220),
        .in(absIn),
        .n(normCount)
    );
    wire [63:0] normAbsIn;
    BITS #(.width(127), .high(63), .low(0)) bits_2712 (
        .y(normAbsIn),
        .in(_T_220)
    );
    wire [1:0] _T_222;
    BITS #(.width(64), .high(40), .low(39)) bits_2713 (
        .y(_T_222),
        .in(normAbsIn)
    );
    wire [38:0] _T_223;
    BITS #(.width(64), .high(38), .low(0)) bits_2714 (
        .y(_T_223),
        .in(normAbsIn)
    );
    wire _T_225;
    wire [38:0] _WTEMP_374;
    PAD_UNSIGNED #(.width(1), .n(39)) u_pad_2715 (
        .y(_WTEMP_374),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(39)) u_neq_2716 (
        .y(_T_225),
        .a(_T_223),
        .b(_WTEMP_374)
    );
    wire [2:0] roundBits;
    CAT #(.width_a(2), .width_b(1)) cat_2717 (
        .y(roundBits),
        .a(_T_222),
        .b(_T_225)
    );
    wire [1:0] _T_226;
    BITS #(.width(3), .high(1), .low(0)) bits_2718 (
        .y(_T_226),
        .in(roundBits)
    );
    wire roundInexact;
    wire [1:0] _WTEMP_375;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2719 (
        .y(_WTEMP_375),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(2)) u_neq_2720 (
        .y(roundInexact),
        .a(_T_226),
        .b(_WTEMP_375)
    );
    wire _T_228;
    EQ_UNSIGNED #(.width(2)) u_eq_2721 (
        .y(_T_228),
        .a(io_roundingMode),
        .b(2'h0)
    );
    wire [1:0] _T_229;
    BITS #(.width(3), .high(2), .low(1)) bits_2722 (
        .y(_T_229),
        .in(roundBits)
    );
    wire [1:0] _T_230;
    BITWISENOT #(.width(2)) bitwisenot_2723 (
        .y(_T_230),
        .in(_T_229)
    );
    wire _T_232;
    wire [1:0] _WTEMP_376;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2724 (
        .y(_WTEMP_376),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(2)) u_eq_2725 (
        .y(_T_232),
        .a(_T_230),
        .b(_WTEMP_376)
    );
    wire [1:0] _T_233;
    BITS #(.width(3), .high(1), .low(0)) bits_2726 (
        .y(_T_233),
        .in(roundBits)
    );
    wire [1:0] _T_234;
    BITWISENOT #(.width(2)) bitwisenot_2727 (
        .y(_T_234),
        .in(_T_233)
    );
    wire _T_236;
    wire [1:0] _WTEMP_377;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2728 (
        .y(_WTEMP_377),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(2)) u_eq_2729 (
        .y(_T_236),
        .a(_T_234),
        .b(_WTEMP_377)
    );
    wire _T_237;
    BITWISEOR #(.width(1)) bitwiseor_2730 (
        .y(_T_237),
        .a(_T_232),
        .b(_T_236)
    );
    wire _T_239;
    MUX_UNSIGNED #(.width(1)) u_mux_2731 (
        .y(_T_239),
        .sel(_T_228),
        .a(_T_237),
        .b(1'h0)
    );
    wire _T_240;
    EQ_UNSIGNED #(.width(2)) u_eq_2732 (
        .y(_T_240),
        .a(io_roundingMode),
        .b(2'h2)
    );
    wire _T_241;
    BITWISEAND #(.width(1)) bitwiseand_2733 (
        .y(_T_241),
        .a(sign),
        .b(roundInexact)
    );
    wire _T_243;
    MUX_UNSIGNED #(.width(1)) u_mux_2734 (
        .y(_T_243),
        .sel(_T_240),
        .a(_T_241),
        .b(1'h0)
    );
    wire _T_244;
    BITWISEOR #(.width(1)) bitwiseor_2735 (
        .y(_T_244),
        .a(_T_239),
        .b(_T_243)
    );
    wire _T_245;
    EQ_UNSIGNED #(.width(2)) u_eq_2736 (
        .y(_T_245),
        .a(io_roundingMode),
        .b(2'h3)
    );
    wire _T_247;
    EQ_UNSIGNED #(.width(1)) u_eq_2737 (
        .y(_T_247),
        .a(sign),
        .b(1'h0)
    );
    wire _T_248;
    BITWISEAND #(.width(1)) bitwiseand_2738 (
        .y(_T_248),
        .a(_T_247),
        .b(roundInexact)
    );
    wire _T_250;
    MUX_UNSIGNED #(.width(1)) u_mux_2739 (
        .y(_T_250),
        .sel(_T_245),
        .a(_T_248),
        .b(1'h0)
    );
    wire round;
    BITWISEOR #(.width(1)) bitwiseor_2740 (
        .y(round),
        .a(_T_244),
        .b(_T_250)
    );
    wire [23:0] _T_252;
    BITS #(.width(64), .high(63), .low(40)) bits_2741 (
        .y(_T_252),
        .in(normAbsIn)
    );
    wire [24:0] unroundedNorm;
    CAT #(.width_a(1), .width_b(24)) cat_2742 (
        .y(unroundedNorm),
        .a(1'h0),
        .b(_T_252)
    );
    wire [25:0] _T_255;
    wire [24:0] _WTEMP_378;
    PAD_UNSIGNED #(.width(1), .n(25)) u_pad_2743 (
        .y(_WTEMP_378),
        .in(1'h1)
    );
    ADD_UNSIGNED #(.width(25)) u_add_2744 (
        .y(_T_255),
        .a(unroundedNorm),
        .b(_WTEMP_378)
    );
    wire [24:0] _T_256;
    TAIL #(.width(26), .n(1)) tail_2745 (
        .y(_T_256),
        .in(_T_255)
    );
    wire [24:0] roundedNorm;
    MUX_UNSIGNED #(.width(25)) u_mux_2746 (
        .y(roundedNorm),
        .sel(round),
        .a(_T_256),
        .b(unroundedNorm)
    );
    wire [5:0] _T_257;
    BITWISENOT #(.width(6)) bitwisenot_2747 (
        .y(_T_257),
        .in(normCount)
    );
    wire [6:0] unroundedExp;
    CAT #(.width_a(1), .width_b(6)) cat_2748 (
        .y(unroundedExp),
        .a(1'h0),
        .b(_T_257)
    );
    wire [7:0] _T_260;
    CAT #(.width_a(1), .width_b(7)) cat_2749 (
        .y(_T_260),
        .a(1'h0),
        .b(unroundedExp)
    );
    wire _T_261;
    BITS #(.width(25), .high(24), .low(24)) bits_2750 (
        .y(_T_261),
        .in(roundedNorm)
    );
    wire [8:0] _T_262;
    wire [7:0] _WTEMP_379;
    PAD_UNSIGNED #(.width(1), .n(8)) u_pad_2751 (
        .y(_WTEMP_379),
        .in(_T_261)
    );
    ADD_UNSIGNED #(.width(8)) u_add_2752 (
        .y(_T_262),
        .a(_T_260),
        .b(_WTEMP_379)
    );
    wire [7:0] roundedExp;
    TAIL #(.width(9), .n(1)) tail_2753 (
        .y(roundedExp),
        .in(_T_262)
    );
    wire _T_263;
    BITS #(.width(64), .high(63), .low(63)) bits_2754 (
        .y(_T_263),
        .in(normAbsIn)
    );
    wire [7:0] _T_265;
    BITS #(.width(8), .high(7), .low(0)) bits_2755 (
        .y(_T_265),
        .in(roundedExp)
    );
    wire [7:0] _T_266;
    assign _T_266 = _T_265;
    wire [8:0] expOut;
    CAT #(.width_a(1), .width_b(8)) cat_2756 (
        .y(expOut),
        .a(_T_263),
        .b(_T_266)
    );
    wire overflow;
    assign overflow = 1'h0;
    wire inexact;
    BITWISEOR #(.width(1)) bitwiseor_2757 (
        .y(inexact),
        .a(roundInexact),
        .b(overflow)
    );
    wire [22:0] _T_267;
    BITS #(.width(25), .high(22), .low(0)) bits_2758 (
        .y(_T_267),
        .in(roundedNorm)
    );
    wire [9:0] _T_268;
    CAT #(.width_a(1), .width_b(9)) cat_2759 (
        .y(_T_268),
        .a(sign),
        .b(expOut)
    );
    wire [32:0] _T_269;
    CAT #(.width_a(10), .width_b(23)) cat_2760 (
        .y(_T_269),
        .a(_T_268),
        .b(_T_267)
    );
    wire [1:0] _T_272;
    CAT #(.width_a(1), .width_b(1)) cat_2761 (
        .y(_T_272),
        .a(1'h0),
        .b(inexact)
    );
    wire [2:0] _T_273;
    assign _T_273 = 3'h0;
    wire [4:0] _T_274;
    CAT #(.width_a(3), .width_b(2)) cat_2762 (
        .y(_T_274),
        .a(_T_273),
        .b(_T_272)
    );
    assign io_exceptionFlags = _T_274;
    assign io_out = _T_269;
endmodule //INToRecFN
module INToRecFN_1(
    input clock,
    input reset,
    input io_signedIn,
    input [63:0] io_in,
    input [1:0] io_roundingMode,
    output [64:0] io_out,
    output [4:0] io_exceptionFlags
);
    wire _T_12;
    BITS #(.width(64), .high(63), .low(63)) bits_2765 (
        .y(_T_12),
        .in(io_in)
    );
    wire sign;
    BITWISEAND #(.width(1)) bitwiseand_2766 (
        .y(sign),
        .a(io_signedIn),
        .b(_T_12)
    );
    wire [64:0] _T_14;
    wire [63:0] _WTEMP_380;
    PAD_UNSIGNED #(.width(1), .n(64)) u_pad_2767 (
        .y(_WTEMP_380),
        .in(1'h0)
    );
    SUB_UNSIGNED #(.width(64)) u_sub_2768 (
        .y(_T_14),
        .a(_WTEMP_380),
        .b(io_in)
    );
    wire [64:0] _T_15;
    ASUINT #(.width(65)) asuint_2769 (
        .y(_T_15),
        .in(_T_14)
    );
    wire [63:0] _T_16;
    TAIL #(.width(65), .n(1)) tail_2770 (
        .y(_T_16),
        .in(_T_15)
    );
    wire [63:0] absIn;
    MUX_UNSIGNED #(.width(64)) u_mux_2771 (
        .y(absIn),
        .sel(sign),
        .a(_T_16),
        .b(io_in)
    );
    wire [63:0] _T_17;
    SHL_UNSIGNED #(.width(64), .n(0)) u_shl_2772 (
        .y(_T_17),
        .in(absIn)
    );
    wire [31:0] _T_18;
    BITS #(.width(64), .high(63), .low(32)) bits_2773 (
        .y(_T_18),
        .in(_T_17)
    );
    wire [31:0] _T_19;
    BITS #(.width(64), .high(31), .low(0)) bits_2774 (
        .y(_T_19),
        .in(_T_17)
    );
    wire _T_21;
    wire [31:0] _WTEMP_381;
    PAD_UNSIGNED #(.width(1), .n(32)) u_pad_2775 (
        .y(_WTEMP_381),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(32)) u_neq_2776 (
        .y(_T_21),
        .a(_T_18),
        .b(_WTEMP_381)
    );
    wire [15:0] _T_22;
    BITS #(.width(32), .high(31), .low(16)) bits_2777 (
        .y(_T_22),
        .in(_T_18)
    );
    wire [15:0] _T_23;
    BITS #(.width(32), .high(15), .low(0)) bits_2778 (
        .y(_T_23),
        .in(_T_18)
    );
    wire _T_25;
    wire [15:0] _WTEMP_382;
    PAD_UNSIGNED #(.width(1), .n(16)) u_pad_2779 (
        .y(_WTEMP_382),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(16)) u_neq_2780 (
        .y(_T_25),
        .a(_T_22),
        .b(_WTEMP_382)
    );
    wire [7:0] _T_26;
    BITS #(.width(16), .high(15), .low(8)) bits_2781 (
        .y(_T_26),
        .in(_T_22)
    );
    wire [7:0] _T_27;
    BITS #(.width(16), .high(7), .low(0)) bits_2782 (
        .y(_T_27),
        .in(_T_22)
    );
    wire _T_29;
    wire [7:0] _WTEMP_383;
    PAD_UNSIGNED #(.width(1), .n(8)) u_pad_2783 (
        .y(_WTEMP_383),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(8)) u_neq_2784 (
        .y(_T_29),
        .a(_T_26),
        .b(_WTEMP_383)
    );
    wire [3:0] _T_30;
    BITS #(.width(8), .high(7), .low(4)) bits_2785 (
        .y(_T_30),
        .in(_T_26)
    );
    wire [3:0] _T_31;
    BITS #(.width(8), .high(3), .low(0)) bits_2786 (
        .y(_T_31),
        .in(_T_26)
    );
    wire _T_33;
    wire [3:0] _WTEMP_384;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_2787 (
        .y(_WTEMP_384),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_2788 (
        .y(_T_33),
        .a(_T_30),
        .b(_WTEMP_384)
    );
    wire _T_34;
    BITS #(.width(4), .high(3), .low(3)) bits_2789 (
        .y(_T_34),
        .in(_T_30)
    );
    wire _T_36;
    BITS #(.width(4), .high(2), .low(2)) bits_2790 (
        .y(_T_36),
        .in(_T_30)
    );
    wire _T_38;
    BITS #(.width(4), .high(1), .low(1)) bits_2791 (
        .y(_T_38),
        .in(_T_30)
    );
    wire [1:0] _T_39;
    wire [1:0] _WTEMP_385;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2792 (
        .y(_WTEMP_385),
        .in(_T_38)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_2793 (
        .y(_T_39),
        .sel(_T_36),
        .a(2'h2),
        .b(_WTEMP_385)
    );
    wire [1:0] _T_40;
    MUX_UNSIGNED #(.width(2)) u_mux_2794 (
        .y(_T_40),
        .sel(_T_34),
        .a(2'h3),
        .b(_T_39)
    );
    wire _T_41;
    BITS #(.width(4), .high(3), .low(3)) bits_2795 (
        .y(_T_41),
        .in(_T_31)
    );
    wire _T_43;
    BITS #(.width(4), .high(2), .low(2)) bits_2796 (
        .y(_T_43),
        .in(_T_31)
    );
    wire _T_45;
    BITS #(.width(4), .high(1), .low(1)) bits_2797 (
        .y(_T_45),
        .in(_T_31)
    );
    wire [1:0] _T_46;
    wire [1:0] _WTEMP_386;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2798 (
        .y(_WTEMP_386),
        .in(_T_45)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_2799 (
        .y(_T_46),
        .sel(_T_43),
        .a(2'h2),
        .b(_WTEMP_386)
    );
    wire [1:0] _T_47;
    MUX_UNSIGNED #(.width(2)) u_mux_2800 (
        .y(_T_47),
        .sel(_T_41),
        .a(2'h3),
        .b(_T_46)
    );
    wire [1:0] _T_48;
    MUX_UNSIGNED #(.width(2)) u_mux_2801 (
        .y(_T_48),
        .sel(_T_33),
        .a(_T_40),
        .b(_T_47)
    );
    wire [2:0] _T_49;
    CAT #(.width_a(1), .width_b(2)) cat_2802 (
        .y(_T_49),
        .a(_T_33),
        .b(_T_48)
    );
    wire [3:0] _T_50;
    BITS #(.width(8), .high(7), .low(4)) bits_2803 (
        .y(_T_50),
        .in(_T_27)
    );
    wire [3:0] _T_51;
    BITS #(.width(8), .high(3), .low(0)) bits_2804 (
        .y(_T_51),
        .in(_T_27)
    );
    wire _T_53;
    wire [3:0] _WTEMP_387;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_2805 (
        .y(_WTEMP_387),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_2806 (
        .y(_T_53),
        .a(_T_50),
        .b(_WTEMP_387)
    );
    wire _T_54;
    BITS #(.width(4), .high(3), .low(3)) bits_2807 (
        .y(_T_54),
        .in(_T_50)
    );
    wire _T_56;
    BITS #(.width(4), .high(2), .low(2)) bits_2808 (
        .y(_T_56),
        .in(_T_50)
    );
    wire _T_58;
    BITS #(.width(4), .high(1), .low(1)) bits_2809 (
        .y(_T_58),
        .in(_T_50)
    );
    wire [1:0] _T_59;
    wire [1:0] _WTEMP_388;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2810 (
        .y(_WTEMP_388),
        .in(_T_58)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_2811 (
        .y(_T_59),
        .sel(_T_56),
        .a(2'h2),
        .b(_WTEMP_388)
    );
    wire [1:0] _T_60;
    MUX_UNSIGNED #(.width(2)) u_mux_2812 (
        .y(_T_60),
        .sel(_T_54),
        .a(2'h3),
        .b(_T_59)
    );
    wire _T_61;
    BITS #(.width(4), .high(3), .low(3)) bits_2813 (
        .y(_T_61),
        .in(_T_51)
    );
    wire _T_63;
    BITS #(.width(4), .high(2), .low(2)) bits_2814 (
        .y(_T_63),
        .in(_T_51)
    );
    wire _T_65;
    BITS #(.width(4), .high(1), .low(1)) bits_2815 (
        .y(_T_65),
        .in(_T_51)
    );
    wire [1:0] _T_66;
    wire [1:0] _WTEMP_389;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2816 (
        .y(_WTEMP_389),
        .in(_T_65)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_2817 (
        .y(_T_66),
        .sel(_T_63),
        .a(2'h2),
        .b(_WTEMP_389)
    );
    wire [1:0] _T_67;
    MUX_UNSIGNED #(.width(2)) u_mux_2818 (
        .y(_T_67),
        .sel(_T_61),
        .a(2'h3),
        .b(_T_66)
    );
    wire [1:0] _T_68;
    MUX_UNSIGNED #(.width(2)) u_mux_2819 (
        .y(_T_68),
        .sel(_T_53),
        .a(_T_60),
        .b(_T_67)
    );
    wire [2:0] _T_69;
    CAT #(.width_a(1), .width_b(2)) cat_2820 (
        .y(_T_69),
        .a(_T_53),
        .b(_T_68)
    );
    wire [2:0] _T_70;
    MUX_UNSIGNED #(.width(3)) u_mux_2821 (
        .y(_T_70),
        .sel(_T_29),
        .a(_T_49),
        .b(_T_69)
    );
    wire [3:0] _T_71;
    CAT #(.width_a(1), .width_b(3)) cat_2822 (
        .y(_T_71),
        .a(_T_29),
        .b(_T_70)
    );
    wire [7:0] _T_72;
    BITS #(.width(16), .high(15), .low(8)) bits_2823 (
        .y(_T_72),
        .in(_T_23)
    );
    wire [7:0] _T_73;
    BITS #(.width(16), .high(7), .low(0)) bits_2824 (
        .y(_T_73),
        .in(_T_23)
    );
    wire _T_75;
    wire [7:0] _WTEMP_390;
    PAD_UNSIGNED #(.width(1), .n(8)) u_pad_2825 (
        .y(_WTEMP_390),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(8)) u_neq_2826 (
        .y(_T_75),
        .a(_T_72),
        .b(_WTEMP_390)
    );
    wire [3:0] _T_76;
    BITS #(.width(8), .high(7), .low(4)) bits_2827 (
        .y(_T_76),
        .in(_T_72)
    );
    wire [3:0] _T_77;
    BITS #(.width(8), .high(3), .low(0)) bits_2828 (
        .y(_T_77),
        .in(_T_72)
    );
    wire _T_79;
    wire [3:0] _WTEMP_391;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_2829 (
        .y(_WTEMP_391),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_2830 (
        .y(_T_79),
        .a(_T_76),
        .b(_WTEMP_391)
    );
    wire _T_80;
    BITS #(.width(4), .high(3), .low(3)) bits_2831 (
        .y(_T_80),
        .in(_T_76)
    );
    wire _T_82;
    BITS #(.width(4), .high(2), .low(2)) bits_2832 (
        .y(_T_82),
        .in(_T_76)
    );
    wire _T_84;
    BITS #(.width(4), .high(1), .low(1)) bits_2833 (
        .y(_T_84),
        .in(_T_76)
    );
    wire [1:0] _T_85;
    wire [1:0] _WTEMP_392;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2834 (
        .y(_WTEMP_392),
        .in(_T_84)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_2835 (
        .y(_T_85),
        .sel(_T_82),
        .a(2'h2),
        .b(_WTEMP_392)
    );
    wire [1:0] _T_86;
    MUX_UNSIGNED #(.width(2)) u_mux_2836 (
        .y(_T_86),
        .sel(_T_80),
        .a(2'h3),
        .b(_T_85)
    );
    wire _T_87;
    BITS #(.width(4), .high(3), .low(3)) bits_2837 (
        .y(_T_87),
        .in(_T_77)
    );
    wire _T_89;
    BITS #(.width(4), .high(2), .low(2)) bits_2838 (
        .y(_T_89),
        .in(_T_77)
    );
    wire _T_91;
    BITS #(.width(4), .high(1), .low(1)) bits_2839 (
        .y(_T_91),
        .in(_T_77)
    );
    wire [1:0] _T_92;
    wire [1:0] _WTEMP_393;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2840 (
        .y(_WTEMP_393),
        .in(_T_91)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_2841 (
        .y(_T_92),
        .sel(_T_89),
        .a(2'h2),
        .b(_WTEMP_393)
    );
    wire [1:0] _T_93;
    MUX_UNSIGNED #(.width(2)) u_mux_2842 (
        .y(_T_93),
        .sel(_T_87),
        .a(2'h3),
        .b(_T_92)
    );
    wire [1:0] _T_94;
    MUX_UNSIGNED #(.width(2)) u_mux_2843 (
        .y(_T_94),
        .sel(_T_79),
        .a(_T_86),
        .b(_T_93)
    );
    wire [2:0] _T_95;
    CAT #(.width_a(1), .width_b(2)) cat_2844 (
        .y(_T_95),
        .a(_T_79),
        .b(_T_94)
    );
    wire [3:0] _T_96;
    BITS #(.width(8), .high(7), .low(4)) bits_2845 (
        .y(_T_96),
        .in(_T_73)
    );
    wire [3:0] _T_97;
    BITS #(.width(8), .high(3), .low(0)) bits_2846 (
        .y(_T_97),
        .in(_T_73)
    );
    wire _T_99;
    wire [3:0] _WTEMP_394;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_2847 (
        .y(_WTEMP_394),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_2848 (
        .y(_T_99),
        .a(_T_96),
        .b(_WTEMP_394)
    );
    wire _T_100;
    BITS #(.width(4), .high(3), .low(3)) bits_2849 (
        .y(_T_100),
        .in(_T_96)
    );
    wire _T_102;
    BITS #(.width(4), .high(2), .low(2)) bits_2850 (
        .y(_T_102),
        .in(_T_96)
    );
    wire _T_104;
    BITS #(.width(4), .high(1), .low(1)) bits_2851 (
        .y(_T_104),
        .in(_T_96)
    );
    wire [1:0] _T_105;
    wire [1:0] _WTEMP_395;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2852 (
        .y(_WTEMP_395),
        .in(_T_104)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_2853 (
        .y(_T_105),
        .sel(_T_102),
        .a(2'h2),
        .b(_WTEMP_395)
    );
    wire [1:0] _T_106;
    MUX_UNSIGNED #(.width(2)) u_mux_2854 (
        .y(_T_106),
        .sel(_T_100),
        .a(2'h3),
        .b(_T_105)
    );
    wire _T_107;
    BITS #(.width(4), .high(3), .low(3)) bits_2855 (
        .y(_T_107),
        .in(_T_97)
    );
    wire _T_109;
    BITS #(.width(4), .high(2), .low(2)) bits_2856 (
        .y(_T_109),
        .in(_T_97)
    );
    wire _T_111;
    BITS #(.width(4), .high(1), .low(1)) bits_2857 (
        .y(_T_111),
        .in(_T_97)
    );
    wire [1:0] _T_112;
    wire [1:0] _WTEMP_396;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2858 (
        .y(_WTEMP_396),
        .in(_T_111)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_2859 (
        .y(_T_112),
        .sel(_T_109),
        .a(2'h2),
        .b(_WTEMP_396)
    );
    wire [1:0] _T_113;
    MUX_UNSIGNED #(.width(2)) u_mux_2860 (
        .y(_T_113),
        .sel(_T_107),
        .a(2'h3),
        .b(_T_112)
    );
    wire [1:0] _T_114;
    MUX_UNSIGNED #(.width(2)) u_mux_2861 (
        .y(_T_114),
        .sel(_T_99),
        .a(_T_106),
        .b(_T_113)
    );
    wire [2:0] _T_115;
    CAT #(.width_a(1), .width_b(2)) cat_2862 (
        .y(_T_115),
        .a(_T_99),
        .b(_T_114)
    );
    wire [2:0] _T_116;
    MUX_UNSIGNED #(.width(3)) u_mux_2863 (
        .y(_T_116),
        .sel(_T_75),
        .a(_T_95),
        .b(_T_115)
    );
    wire [3:0] _T_117;
    CAT #(.width_a(1), .width_b(3)) cat_2864 (
        .y(_T_117),
        .a(_T_75),
        .b(_T_116)
    );
    wire [3:0] _T_118;
    MUX_UNSIGNED #(.width(4)) u_mux_2865 (
        .y(_T_118),
        .sel(_T_25),
        .a(_T_71),
        .b(_T_117)
    );
    wire [4:0] _T_119;
    CAT #(.width_a(1), .width_b(4)) cat_2866 (
        .y(_T_119),
        .a(_T_25),
        .b(_T_118)
    );
    wire [15:0] _T_120;
    BITS #(.width(32), .high(31), .low(16)) bits_2867 (
        .y(_T_120),
        .in(_T_19)
    );
    wire [15:0] _T_121;
    BITS #(.width(32), .high(15), .low(0)) bits_2868 (
        .y(_T_121),
        .in(_T_19)
    );
    wire _T_123;
    wire [15:0] _WTEMP_397;
    PAD_UNSIGNED #(.width(1), .n(16)) u_pad_2869 (
        .y(_WTEMP_397),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(16)) u_neq_2870 (
        .y(_T_123),
        .a(_T_120),
        .b(_WTEMP_397)
    );
    wire [7:0] _T_124;
    BITS #(.width(16), .high(15), .low(8)) bits_2871 (
        .y(_T_124),
        .in(_T_120)
    );
    wire [7:0] _T_125;
    BITS #(.width(16), .high(7), .low(0)) bits_2872 (
        .y(_T_125),
        .in(_T_120)
    );
    wire _T_127;
    wire [7:0] _WTEMP_398;
    PAD_UNSIGNED #(.width(1), .n(8)) u_pad_2873 (
        .y(_WTEMP_398),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(8)) u_neq_2874 (
        .y(_T_127),
        .a(_T_124),
        .b(_WTEMP_398)
    );
    wire [3:0] _T_128;
    BITS #(.width(8), .high(7), .low(4)) bits_2875 (
        .y(_T_128),
        .in(_T_124)
    );
    wire [3:0] _T_129;
    BITS #(.width(8), .high(3), .low(0)) bits_2876 (
        .y(_T_129),
        .in(_T_124)
    );
    wire _T_131;
    wire [3:0] _WTEMP_399;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_2877 (
        .y(_WTEMP_399),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_2878 (
        .y(_T_131),
        .a(_T_128),
        .b(_WTEMP_399)
    );
    wire _T_132;
    BITS #(.width(4), .high(3), .low(3)) bits_2879 (
        .y(_T_132),
        .in(_T_128)
    );
    wire _T_134;
    BITS #(.width(4), .high(2), .low(2)) bits_2880 (
        .y(_T_134),
        .in(_T_128)
    );
    wire _T_136;
    BITS #(.width(4), .high(1), .low(1)) bits_2881 (
        .y(_T_136),
        .in(_T_128)
    );
    wire [1:0] _T_137;
    wire [1:0] _WTEMP_400;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2882 (
        .y(_WTEMP_400),
        .in(_T_136)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_2883 (
        .y(_T_137),
        .sel(_T_134),
        .a(2'h2),
        .b(_WTEMP_400)
    );
    wire [1:0] _T_138;
    MUX_UNSIGNED #(.width(2)) u_mux_2884 (
        .y(_T_138),
        .sel(_T_132),
        .a(2'h3),
        .b(_T_137)
    );
    wire _T_139;
    BITS #(.width(4), .high(3), .low(3)) bits_2885 (
        .y(_T_139),
        .in(_T_129)
    );
    wire _T_141;
    BITS #(.width(4), .high(2), .low(2)) bits_2886 (
        .y(_T_141),
        .in(_T_129)
    );
    wire _T_143;
    BITS #(.width(4), .high(1), .low(1)) bits_2887 (
        .y(_T_143),
        .in(_T_129)
    );
    wire [1:0] _T_144;
    wire [1:0] _WTEMP_401;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2888 (
        .y(_WTEMP_401),
        .in(_T_143)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_2889 (
        .y(_T_144),
        .sel(_T_141),
        .a(2'h2),
        .b(_WTEMP_401)
    );
    wire [1:0] _T_145;
    MUX_UNSIGNED #(.width(2)) u_mux_2890 (
        .y(_T_145),
        .sel(_T_139),
        .a(2'h3),
        .b(_T_144)
    );
    wire [1:0] _T_146;
    MUX_UNSIGNED #(.width(2)) u_mux_2891 (
        .y(_T_146),
        .sel(_T_131),
        .a(_T_138),
        .b(_T_145)
    );
    wire [2:0] _T_147;
    CAT #(.width_a(1), .width_b(2)) cat_2892 (
        .y(_T_147),
        .a(_T_131),
        .b(_T_146)
    );
    wire [3:0] _T_148;
    BITS #(.width(8), .high(7), .low(4)) bits_2893 (
        .y(_T_148),
        .in(_T_125)
    );
    wire [3:0] _T_149;
    BITS #(.width(8), .high(3), .low(0)) bits_2894 (
        .y(_T_149),
        .in(_T_125)
    );
    wire _T_151;
    wire [3:0] _WTEMP_402;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_2895 (
        .y(_WTEMP_402),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_2896 (
        .y(_T_151),
        .a(_T_148),
        .b(_WTEMP_402)
    );
    wire _T_152;
    BITS #(.width(4), .high(3), .low(3)) bits_2897 (
        .y(_T_152),
        .in(_T_148)
    );
    wire _T_154;
    BITS #(.width(4), .high(2), .low(2)) bits_2898 (
        .y(_T_154),
        .in(_T_148)
    );
    wire _T_156;
    BITS #(.width(4), .high(1), .low(1)) bits_2899 (
        .y(_T_156),
        .in(_T_148)
    );
    wire [1:0] _T_157;
    wire [1:0] _WTEMP_403;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2900 (
        .y(_WTEMP_403),
        .in(_T_156)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_2901 (
        .y(_T_157),
        .sel(_T_154),
        .a(2'h2),
        .b(_WTEMP_403)
    );
    wire [1:0] _T_158;
    MUX_UNSIGNED #(.width(2)) u_mux_2902 (
        .y(_T_158),
        .sel(_T_152),
        .a(2'h3),
        .b(_T_157)
    );
    wire _T_159;
    BITS #(.width(4), .high(3), .low(3)) bits_2903 (
        .y(_T_159),
        .in(_T_149)
    );
    wire _T_161;
    BITS #(.width(4), .high(2), .low(2)) bits_2904 (
        .y(_T_161),
        .in(_T_149)
    );
    wire _T_163;
    BITS #(.width(4), .high(1), .low(1)) bits_2905 (
        .y(_T_163),
        .in(_T_149)
    );
    wire [1:0] _T_164;
    wire [1:0] _WTEMP_404;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2906 (
        .y(_WTEMP_404),
        .in(_T_163)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_2907 (
        .y(_T_164),
        .sel(_T_161),
        .a(2'h2),
        .b(_WTEMP_404)
    );
    wire [1:0] _T_165;
    MUX_UNSIGNED #(.width(2)) u_mux_2908 (
        .y(_T_165),
        .sel(_T_159),
        .a(2'h3),
        .b(_T_164)
    );
    wire [1:0] _T_166;
    MUX_UNSIGNED #(.width(2)) u_mux_2909 (
        .y(_T_166),
        .sel(_T_151),
        .a(_T_158),
        .b(_T_165)
    );
    wire [2:0] _T_167;
    CAT #(.width_a(1), .width_b(2)) cat_2910 (
        .y(_T_167),
        .a(_T_151),
        .b(_T_166)
    );
    wire [2:0] _T_168;
    MUX_UNSIGNED #(.width(3)) u_mux_2911 (
        .y(_T_168),
        .sel(_T_127),
        .a(_T_147),
        .b(_T_167)
    );
    wire [3:0] _T_169;
    CAT #(.width_a(1), .width_b(3)) cat_2912 (
        .y(_T_169),
        .a(_T_127),
        .b(_T_168)
    );
    wire [7:0] _T_170;
    BITS #(.width(16), .high(15), .low(8)) bits_2913 (
        .y(_T_170),
        .in(_T_121)
    );
    wire [7:0] _T_171;
    BITS #(.width(16), .high(7), .low(0)) bits_2914 (
        .y(_T_171),
        .in(_T_121)
    );
    wire _T_173;
    wire [7:0] _WTEMP_405;
    PAD_UNSIGNED #(.width(1), .n(8)) u_pad_2915 (
        .y(_WTEMP_405),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(8)) u_neq_2916 (
        .y(_T_173),
        .a(_T_170),
        .b(_WTEMP_405)
    );
    wire [3:0] _T_174;
    BITS #(.width(8), .high(7), .low(4)) bits_2917 (
        .y(_T_174),
        .in(_T_170)
    );
    wire [3:0] _T_175;
    BITS #(.width(8), .high(3), .low(0)) bits_2918 (
        .y(_T_175),
        .in(_T_170)
    );
    wire _T_177;
    wire [3:0] _WTEMP_406;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_2919 (
        .y(_WTEMP_406),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_2920 (
        .y(_T_177),
        .a(_T_174),
        .b(_WTEMP_406)
    );
    wire _T_178;
    BITS #(.width(4), .high(3), .low(3)) bits_2921 (
        .y(_T_178),
        .in(_T_174)
    );
    wire _T_180;
    BITS #(.width(4), .high(2), .low(2)) bits_2922 (
        .y(_T_180),
        .in(_T_174)
    );
    wire _T_182;
    BITS #(.width(4), .high(1), .low(1)) bits_2923 (
        .y(_T_182),
        .in(_T_174)
    );
    wire [1:0] _T_183;
    wire [1:0] _WTEMP_407;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2924 (
        .y(_WTEMP_407),
        .in(_T_182)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_2925 (
        .y(_T_183),
        .sel(_T_180),
        .a(2'h2),
        .b(_WTEMP_407)
    );
    wire [1:0] _T_184;
    MUX_UNSIGNED #(.width(2)) u_mux_2926 (
        .y(_T_184),
        .sel(_T_178),
        .a(2'h3),
        .b(_T_183)
    );
    wire _T_185;
    BITS #(.width(4), .high(3), .low(3)) bits_2927 (
        .y(_T_185),
        .in(_T_175)
    );
    wire _T_187;
    BITS #(.width(4), .high(2), .low(2)) bits_2928 (
        .y(_T_187),
        .in(_T_175)
    );
    wire _T_189;
    BITS #(.width(4), .high(1), .low(1)) bits_2929 (
        .y(_T_189),
        .in(_T_175)
    );
    wire [1:0] _T_190;
    wire [1:0] _WTEMP_408;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2930 (
        .y(_WTEMP_408),
        .in(_T_189)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_2931 (
        .y(_T_190),
        .sel(_T_187),
        .a(2'h2),
        .b(_WTEMP_408)
    );
    wire [1:0] _T_191;
    MUX_UNSIGNED #(.width(2)) u_mux_2932 (
        .y(_T_191),
        .sel(_T_185),
        .a(2'h3),
        .b(_T_190)
    );
    wire [1:0] _T_192;
    MUX_UNSIGNED #(.width(2)) u_mux_2933 (
        .y(_T_192),
        .sel(_T_177),
        .a(_T_184),
        .b(_T_191)
    );
    wire [2:0] _T_193;
    CAT #(.width_a(1), .width_b(2)) cat_2934 (
        .y(_T_193),
        .a(_T_177),
        .b(_T_192)
    );
    wire [3:0] _T_194;
    BITS #(.width(8), .high(7), .low(4)) bits_2935 (
        .y(_T_194),
        .in(_T_171)
    );
    wire [3:0] _T_195;
    BITS #(.width(8), .high(3), .low(0)) bits_2936 (
        .y(_T_195),
        .in(_T_171)
    );
    wire _T_197;
    wire [3:0] _WTEMP_409;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_2937 (
        .y(_WTEMP_409),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_2938 (
        .y(_T_197),
        .a(_T_194),
        .b(_WTEMP_409)
    );
    wire _T_198;
    BITS #(.width(4), .high(3), .low(3)) bits_2939 (
        .y(_T_198),
        .in(_T_194)
    );
    wire _T_200;
    BITS #(.width(4), .high(2), .low(2)) bits_2940 (
        .y(_T_200),
        .in(_T_194)
    );
    wire _T_202;
    BITS #(.width(4), .high(1), .low(1)) bits_2941 (
        .y(_T_202),
        .in(_T_194)
    );
    wire [1:0] _T_203;
    wire [1:0] _WTEMP_410;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2942 (
        .y(_WTEMP_410),
        .in(_T_202)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_2943 (
        .y(_T_203),
        .sel(_T_200),
        .a(2'h2),
        .b(_WTEMP_410)
    );
    wire [1:0] _T_204;
    MUX_UNSIGNED #(.width(2)) u_mux_2944 (
        .y(_T_204),
        .sel(_T_198),
        .a(2'h3),
        .b(_T_203)
    );
    wire _T_205;
    BITS #(.width(4), .high(3), .low(3)) bits_2945 (
        .y(_T_205),
        .in(_T_195)
    );
    wire _T_207;
    BITS #(.width(4), .high(2), .low(2)) bits_2946 (
        .y(_T_207),
        .in(_T_195)
    );
    wire _T_209;
    BITS #(.width(4), .high(1), .low(1)) bits_2947 (
        .y(_T_209),
        .in(_T_195)
    );
    wire [1:0] _T_210;
    wire [1:0] _WTEMP_411;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2948 (
        .y(_WTEMP_411),
        .in(_T_209)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_2949 (
        .y(_T_210),
        .sel(_T_207),
        .a(2'h2),
        .b(_WTEMP_411)
    );
    wire [1:0] _T_211;
    MUX_UNSIGNED #(.width(2)) u_mux_2950 (
        .y(_T_211),
        .sel(_T_205),
        .a(2'h3),
        .b(_T_210)
    );
    wire [1:0] _T_212;
    MUX_UNSIGNED #(.width(2)) u_mux_2951 (
        .y(_T_212),
        .sel(_T_197),
        .a(_T_204),
        .b(_T_211)
    );
    wire [2:0] _T_213;
    CAT #(.width_a(1), .width_b(2)) cat_2952 (
        .y(_T_213),
        .a(_T_197),
        .b(_T_212)
    );
    wire [2:0] _T_214;
    MUX_UNSIGNED #(.width(3)) u_mux_2953 (
        .y(_T_214),
        .sel(_T_173),
        .a(_T_193),
        .b(_T_213)
    );
    wire [3:0] _T_215;
    CAT #(.width_a(1), .width_b(3)) cat_2954 (
        .y(_T_215),
        .a(_T_173),
        .b(_T_214)
    );
    wire [3:0] _T_216;
    MUX_UNSIGNED #(.width(4)) u_mux_2955 (
        .y(_T_216),
        .sel(_T_123),
        .a(_T_169),
        .b(_T_215)
    );
    wire [4:0] _T_217;
    CAT #(.width_a(1), .width_b(4)) cat_2956 (
        .y(_T_217),
        .a(_T_123),
        .b(_T_216)
    );
    wire [4:0] _T_218;
    MUX_UNSIGNED #(.width(5)) u_mux_2957 (
        .y(_T_218),
        .sel(_T_21),
        .a(_T_119),
        .b(_T_217)
    );
    wire [5:0] _T_219;
    CAT #(.width_a(1), .width_b(5)) cat_2958 (
        .y(_T_219),
        .a(_T_21),
        .b(_T_218)
    );
    wire [5:0] normCount;
    BITWISENOT #(.width(6)) bitwisenot_2959 (
        .y(normCount),
        .in(_T_219)
    );
    wire [126:0] _T_220;
    DSHL_UNSIGNED #(.width_in(64), .width_n(6)) u_dshl_2960 (
        .y(_T_220),
        .in(absIn),
        .n(normCount)
    );
    wire [63:0] normAbsIn;
    BITS #(.width(127), .high(63), .low(0)) bits_2961 (
        .y(normAbsIn),
        .in(_T_220)
    );
    wire [1:0] _T_222;
    BITS #(.width(64), .high(11), .low(10)) bits_2962 (
        .y(_T_222),
        .in(normAbsIn)
    );
    wire [9:0] _T_223;
    BITS #(.width(64), .high(9), .low(0)) bits_2963 (
        .y(_T_223),
        .in(normAbsIn)
    );
    wire _T_225;
    wire [9:0] _WTEMP_412;
    PAD_UNSIGNED #(.width(1), .n(10)) u_pad_2964 (
        .y(_WTEMP_412),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(10)) u_neq_2965 (
        .y(_T_225),
        .a(_T_223),
        .b(_WTEMP_412)
    );
    wire [2:0] roundBits;
    CAT #(.width_a(2), .width_b(1)) cat_2966 (
        .y(roundBits),
        .a(_T_222),
        .b(_T_225)
    );
    wire [1:0] _T_226;
    BITS #(.width(3), .high(1), .low(0)) bits_2967 (
        .y(_T_226),
        .in(roundBits)
    );
    wire roundInexact;
    wire [1:0] _WTEMP_413;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2968 (
        .y(_WTEMP_413),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(2)) u_neq_2969 (
        .y(roundInexact),
        .a(_T_226),
        .b(_WTEMP_413)
    );
    wire _T_228;
    EQ_UNSIGNED #(.width(2)) u_eq_2970 (
        .y(_T_228),
        .a(io_roundingMode),
        .b(2'h0)
    );
    wire [1:0] _T_229;
    BITS #(.width(3), .high(2), .low(1)) bits_2971 (
        .y(_T_229),
        .in(roundBits)
    );
    wire [1:0] _T_230;
    BITWISENOT #(.width(2)) bitwisenot_2972 (
        .y(_T_230),
        .in(_T_229)
    );
    wire _T_232;
    wire [1:0] _WTEMP_414;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2973 (
        .y(_WTEMP_414),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(2)) u_eq_2974 (
        .y(_T_232),
        .a(_T_230),
        .b(_WTEMP_414)
    );
    wire [1:0] _T_233;
    BITS #(.width(3), .high(1), .low(0)) bits_2975 (
        .y(_T_233),
        .in(roundBits)
    );
    wire [1:0] _T_234;
    BITWISENOT #(.width(2)) bitwisenot_2976 (
        .y(_T_234),
        .in(_T_233)
    );
    wire _T_236;
    wire [1:0] _WTEMP_415;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_2977 (
        .y(_WTEMP_415),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(2)) u_eq_2978 (
        .y(_T_236),
        .a(_T_234),
        .b(_WTEMP_415)
    );
    wire _T_237;
    BITWISEOR #(.width(1)) bitwiseor_2979 (
        .y(_T_237),
        .a(_T_232),
        .b(_T_236)
    );
    wire _T_239;
    MUX_UNSIGNED #(.width(1)) u_mux_2980 (
        .y(_T_239),
        .sel(_T_228),
        .a(_T_237),
        .b(1'h0)
    );
    wire _T_240;
    EQ_UNSIGNED #(.width(2)) u_eq_2981 (
        .y(_T_240),
        .a(io_roundingMode),
        .b(2'h2)
    );
    wire _T_241;
    BITWISEAND #(.width(1)) bitwiseand_2982 (
        .y(_T_241),
        .a(sign),
        .b(roundInexact)
    );
    wire _T_243;
    MUX_UNSIGNED #(.width(1)) u_mux_2983 (
        .y(_T_243),
        .sel(_T_240),
        .a(_T_241),
        .b(1'h0)
    );
    wire _T_244;
    BITWISEOR #(.width(1)) bitwiseor_2984 (
        .y(_T_244),
        .a(_T_239),
        .b(_T_243)
    );
    wire _T_245;
    EQ_UNSIGNED #(.width(2)) u_eq_2985 (
        .y(_T_245),
        .a(io_roundingMode),
        .b(2'h3)
    );
    wire _T_247;
    EQ_UNSIGNED #(.width(1)) u_eq_2986 (
        .y(_T_247),
        .a(sign),
        .b(1'h0)
    );
    wire _T_248;
    BITWISEAND #(.width(1)) bitwiseand_2987 (
        .y(_T_248),
        .a(_T_247),
        .b(roundInexact)
    );
    wire _T_250;
    MUX_UNSIGNED #(.width(1)) u_mux_2988 (
        .y(_T_250),
        .sel(_T_245),
        .a(_T_248),
        .b(1'h0)
    );
    wire round;
    BITWISEOR #(.width(1)) bitwiseor_2989 (
        .y(round),
        .a(_T_244),
        .b(_T_250)
    );
    wire [52:0] _T_252;
    BITS #(.width(64), .high(63), .low(11)) bits_2990 (
        .y(_T_252),
        .in(normAbsIn)
    );
    wire [53:0] unroundedNorm;
    CAT #(.width_a(1), .width_b(53)) cat_2991 (
        .y(unroundedNorm),
        .a(1'h0),
        .b(_T_252)
    );
    wire [54:0] _T_255;
    wire [53:0] _WTEMP_416;
    PAD_UNSIGNED #(.width(1), .n(54)) u_pad_2992 (
        .y(_WTEMP_416),
        .in(1'h1)
    );
    ADD_UNSIGNED #(.width(54)) u_add_2993 (
        .y(_T_255),
        .a(unroundedNorm),
        .b(_WTEMP_416)
    );
    wire [53:0] _T_256;
    TAIL #(.width(55), .n(1)) tail_2994 (
        .y(_T_256),
        .in(_T_255)
    );
    wire [53:0] roundedNorm;
    MUX_UNSIGNED #(.width(54)) u_mux_2995 (
        .y(roundedNorm),
        .sel(round),
        .a(_T_256),
        .b(unroundedNorm)
    );
    wire [5:0] _T_257;
    BITWISENOT #(.width(6)) bitwisenot_2996 (
        .y(_T_257),
        .in(normCount)
    );
    wire [9:0] unroundedExp;
    CAT #(.width_a(4), .width_b(6)) cat_2997 (
        .y(unroundedExp),
        .a(4'h0),
        .b(_T_257)
    );
    wire [10:0] _T_260;
    CAT #(.width_a(1), .width_b(10)) cat_2998 (
        .y(_T_260),
        .a(1'h0),
        .b(unroundedExp)
    );
    wire _T_261;
    BITS #(.width(54), .high(53), .low(53)) bits_2999 (
        .y(_T_261),
        .in(roundedNorm)
    );
    wire [11:0] _T_262;
    wire [10:0] _WTEMP_417;
    PAD_UNSIGNED #(.width(1), .n(11)) u_pad_3000 (
        .y(_WTEMP_417),
        .in(_T_261)
    );
    ADD_UNSIGNED #(.width(11)) u_add_3001 (
        .y(_T_262),
        .a(_T_260),
        .b(_WTEMP_417)
    );
    wire [10:0] roundedExp;
    TAIL #(.width(12), .n(1)) tail_3002 (
        .y(roundedExp),
        .in(_T_262)
    );
    wire _T_263;
    BITS #(.width(64), .high(63), .low(63)) bits_3003 (
        .y(_T_263),
        .in(normAbsIn)
    );
    wire [10:0] _T_265;
    BITS #(.width(11), .high(10), .low(0)) bits_3004 (
        .y(_T_265),
        .in(roundedExp)
    );
    wire [10:0] _T_266;
    assign _T_266 = _T_265;
    wire [11:0] expOut;
    CAT #(.width_a(1), .width_b(11)) cat_3005 (
        .y(expOut),
        .a(_T_263),
        .b(_T_266)
    );
    wire overflow;
    assign overflow = 1'h0;
    wire inexact;
    BITWISEOR #(.width(1)) bitwiseor_3006 (
        .y(inexact),
        .a(roundInexact),
        .b(overflow)
    );
    wire [51:0] _T_267;
    BITS #(.width(54), .high(51), .low(0)) bits_3007 (
        .y(_T_267),
        .in(roundedNorm)
    );
    wire [12:0] _T_268;
    CAT #(.width_a(1), .width_b(12)) cat_3008 (
        .y(_T_268),
        .a(sign),
        .b(expOut)
    );
    wire [64:0] _T_269;
    CAT #(.width_a(13), .width_b(52)) cat_3009 (
        .y(_T_269),
        .a(_T_268),
        .b(_T_267)
    );
    wire [1:0] _T_272;
    CAT #(.width_a(1), .width_b(1)) cat_3010 (
        .y(_T_272),
        .a(1'h0),
        .b(inexact)
    );
    wire [2:0] _T_273;
    assign _T_273 = 3'h0;
    wire [4:0] _T_274;
    CAT #(.width_a(3), .width_b(2)) cat_3011 (
        .y(_T_274),
        .a(_T_273),
        .b(_T_272)
    );
    assign io_exceptionFlags = _T_274;
    assign io_out = _T_269;
endmodule //INToRecFN_1
module FPToFP(
    input clock,
    input reset,
    input io_in_valid,
    input [4:0] io_in_bits_cmd,
    input io_in_bits_ldst,
    input io_in_bits_wen,
    input io_in_bits_ren1,
    input io_in_bits_ren2,
    input io_in_bits_ren3,
    input io_in_bits_swap12,
    input io_in_bits_swap23,
    input io_in_bits_single,
    input io_in_bits_fromint,
    input io_in_bits_toint,
    input io_in_bits_fastpipe,
    input io_in_bits_fma,
    input io_in_bits_div,
    input io_in_bits_sqrt,
    input io_in_bits_wflags,
    input [2:0] io_in_bits_rm,
    input [1:0] io_in_bits_typ,
    input [64:0] io_in_bits_in1,
    input [64:0] io_in_bits_in2,
    input [64:0] io_in_bits_in3,
    output io_out_valid,
    output [64:0] io_out_bits_data,
    output [4:0] io_out_bits_exc,
    input io_lt
);
    wire __T_134__q;
    wire __T_134__d;
    DFF_POSCLK #(.width(1)) _T_134 (
        .q(__T_134__q),
        .d(__T_134__d),
        .clk(clock)
    );
    wire _WTEMP_423;
    MUX_UNSIGNED #(.width(1)) u_mux_3057 (
        .y(__T_134__d),
        .sel(reset),
        .a(1'h0),
        .b(_WTEMP_423)
    );
    wire [4:0] __T_157_cmd__q;
    wire [4:0] __T_157_cmd__d;
    DFF_POSCLK #(.width(5)) _T_157_cmd (
        .q(__T_157_cmd__q),
        .d(__T_157_cmd__d),
        .clk(clock)
    );
    wire __T_157_ldst__q;
    wire __T_157_ldst__d;
    DFF_POSCLK #(.width(1)) _T_157_ldst (
        .q(__T_157_ldst__q),
        .d(__T_157_ldst__d),
        .clk(clock)
    );
    wire __T_157_wen__q;
    wire __T_157_wen__d;
    DFF_POSCLK #(.width(1)) _T_157_wen (
        .q(__T_157_wen__q),
        .d(__T_157_wen__d),
        .clk(clock)
    );
    wire __T_157_ren1__q;
    wire __T_157_ren1__d;
    DFF_POSCLK #(.width(1)) _T_157_ren1 (
        .q(__T_157_ren1__q),
        .d(__T_157_ren1__d),
        .clk(clock)
    );
    wire __T_157_ren2__q;
    wire __T_157_ren2__d;
    DFF_POSCLK #(.width(1)) _T_157_ren2 (
        .q(__T_157_ren2__q),
        .d(__T_157_ren2__d),
        .clk(clock)
    );
    wire __T_157_ren3__q;
    wire __T_157_ren3__d;
    DFF_POSCLK #(.width(1)) _T_157_ren3 (
        .q(__T_157_ren3__q),
        .d(__T_157_ren3__d),
        .clk(clock)
    );
    wire __T_157_swap12__q;
    wire __T_157_swap12__d;
    DFF_POSCLK #(.width(1)) _T_157_swap12 (
        .q(__T_157_swap12__q),
        .d(__T_157_swap12__d),
        .clk(clock)
    );
    wire __T_157_swap23__q;
    wire __T_157_swap23__d;
    DFF_POSCLK #(.width(1)) _T_157_swap23 (
        .q(__T_157_swap23__q),
        .d(__T_157_swap23__d),
        .clk(clock)
    );
    wire __T_157_single__q;
    wire __T_157_single__d;
    DFF_POSCLK #(.width(1)) _T_157_single (
        .q(__T_157_single__q),
        .d(__T_157_single__d),
        .clk(clock)
    );
    wire __T_157_fromint__q;
    wire __T_157_fromint__d;
    DFF_POSCLK #(.width(1)) _T_157_fromint (
        .q(__T_157_fromint__q),
        .d(__T_157_fromint__d),
        .clk(clock)
    );
    wire __T_157_toint__q;
    wire __T_157_toint__d;
    DFF_POSCLK #(.width(1)) _T_157_toint (
        .q(__T_157_toint__q),
        .d(__T_157_toint__d),
        .clk(clock)
    );
    wire __T_157_fastpipe__q;
    wire __T_157_fastpipe__d;
    DFF_POSCLK #(.width(1)) _T_157_fastpipe (
        .q(__T_157_fastpipe__q),
        .d(__T_157_fastpipe__d),
        .clk(clock)
    );
    wire __T_157_fma__q;
    wire __T_157_fma__d;
    DFF_POSCLK #(.width(1)) _T_157_fma (
        .q(__T_157_fma__q),
        .d(__T_157_fma__d),
        .clk(clock)
    );
    wire __T_157_div__q;
    wire __T_157_div__d;
    DFF_POSCLK #(.width(1)) _T_157_div (
        .q(__T_157_div__q),
        .d(__T_157_div__d),
        .clk(clock)
    );
    wire __T_157_sqrt__q;
    wire __T_157_sqrt__d;
    DFF_POSCLK #(.width(1)) _T_157_sqrt (
        .q(__T_157_sqrt__q),
        .d(__T_157_sqrt__d),
        .clk(clock)
    );
    wire __T_157_wflags__q;
    wire __T_157_wflags__d;
    DFF_POSCLK #(.width(1)) _T_157_wflags (
        .q(__T_157_wflags__q),
        .d(__T_157_wflags__d),
        .clk(clock)
    );
    wire [2:0] __T_157_rm__q;
    wire [2:0] __T_157_rm__d;
    DFF_POSCLK #(.width(3)) _T_157_rm (
        .q(__T_157_rm__q),
        .d(__T_157_rm__d),
        .clk(clock)
    );
    wire [1:0] __T_157_typ__q;
    wire [1:0] __T_157_typ__d;
    DFF_POSCLK #(.width(2)) _T_157_typ (
        .q(__T_157_typ__q),
        .d(__T_157_typ__d),
        .clk(clock)
    );
    wire [64:0] __T_157_in1__q;
    wire [64:0] __T_157_in1__d;
    DFF_POSCLK #(.width(65)) _T_157_in1 (
        .q(__T_157_in1__q),
        .d(__T_157_in1__d),
        .clk(clock)
    );
    wire [64:0] __T_157_in2__q;
    wire [64:0] __T_157_in2__d;
    DFF_POSCLK #(.width(65)) _T_157_in2 (
        .q(__T_157_in2__q),
        .d(__T_157_in2__d),
        .clk(clock)
    );
    wire [64:0] __T_157_in3__q;
    wire [64:0] __T_157_in3__d;
    DFF_POSCLK #(.width(65)) _T_157_in3 (
        .q(__T_157_in3__q),
        .d(__T_157_in3__d),
        .clk(clock)
    );
    wire in_valid;
    wire [4:0] in_bits_cmd;
    wire in_bits_ldst;
    wire in_bits_wen;
    wire in_bits_ren1;
    wire in_bits_ren2;
    wire in_bits_ren3;
    wire in_bits_swap12;
    wire in_bits_swap23;
    wire in_bits_single;
    wire in_bits_fromint;
    wire in_bits_toint;
    wire in_bits_fastpipe;
    wire in_bits_fma;
    wire in_bits_div;
    wire in_bits_sqrt;
    wire in_bits_wflags;
    wire [2:0] in_bits_rm;
    wire [1:0] in_bits_typ;
    wire [64:0] in_bits_in1;
    wire [64:0] in_bits_in2;
    wire [64:0] in_bits_in3;
    wire _T_272;
    BITS #(.width(3), .high(1), .low(1)) bits_3058 (
        .y(_T_272),
        .in(in_bits_rm)
    );
    wire [64:0] _T_273;
    BITWISEXOR #(.width(65)) bitwisexor_3059 (
        .y(_T_273),
        .a(in_bits_in1),
        .b(in_bits_in2)
    );
    wire _T_274;
    BITS #(.width(3), .high(0), .low(0)) bits_3060 (
        .y(_T_274),
        .in(in_bits_rm)
    );
    wire [64:0] _T_275;
    BITWISENOT #(.width(65)) bitwisenot_3061 (
        .y(_T_275),
        .in(in_bits_in2)
    );
    wire [64:0] _T_276;
    MUX_UNSIGNED #(.width(65)) u_mux_3062 (
        .y(_T_276),
        .sel(_T_274),
        .a(_T_275),
        .b(in_bits_in2)
    );
    wire [64:0] signNum;
    MUX_UNSIGNED #(.width(65)) u_mux_3063 (
        .y(signNum),
        .sel(_T_272),
        .a(_T_273),
        .b(_T_276)
    );
    wire _T_277;
    BITS #(.width(65), .high(32), .low(32)) bits_3064 (
        .y(_T_277),
        .in(signNum)
    );
    wire [31:0] _T_278;
    BITS #(.width(65), .high(31), .low(0)) bits_3065 (
        .y(_T_278),
        .in(in_bits_in1)
    );
    wire [32:0] fsgnj_s;
    CAT #(.width_a(1), .width_b(32)) cat_3066 (
        .y(fsgnj_s),
        .a(_T_277),
        .b(_T_278)
    );
    wire [31:0] _T_279;
    SHR_UNSIGNED #(.width(65), .n(33)) u_shr_3067 (
        .y(_T_279),
        .in(in_bits_in1)
    );
    wire [64:0] _T_280;
    CAT #(.width_a(32), .width_b(33)) cat_3068 (
        .y(_T_280),
        .a(_T_279),
        .b(fsgnj_s)
    );
    wire _T_281;
    BITS #(.width(65), .high(64), .low(64)) bits_3069 (
        .y(_T_281),
        .in(signNum)
    );
    wire [63:0] _T_282;
    BITS #(.width(65), .high(63), .low(0)) bits_3070 (
        .y(_T_282),
        .in(in_bits_in1)
    );
    wire [64:0] _T_283;
    CAT #(.width_a(1), .width_b(64)) cat_3071 (
        .y(_T_283),
        .a(_T_281),
        .b(_T_282)
    );
    wire [64:0] fsgnj;
    MUX_UNSIGNED #(.width(65)) u_mux_3072 (
        .y(fsgnj),
        .sel(in_bits_single),
        .a(_T_280),
        .b(_T_283)
    );
    wire [64:0] mux_data;
    wire [4:0] mux_exc;
    wire [4:0] _T_292;
    wire [4:0] _WTEMP_424;
    PAD_UNSIGNED #(.width(4), .n(5)) u_pad_3073 (
        .y(_WTEMP_424),
        .in(4'hD)
    );
    BITWISEAND #(.width(5)) bitwiseand_3074 (
        .y(_T_292),
        .a(in_bits_cmd),
        .b(_WTEMP_424)
    );
    wire _T_293;
    wire [4:0] _WTEMP_425;
    PAD_UNSIGNED #(.width(3), .n(5)) u_pad_3075 (
        .y(_WTEMP_425),
        .in(3'h5)
    );
    EQ_UNSIGNED #(.width(5)) u_eq_3076 (
        .y(_T_293),
        .a(_WTEMP_425),
        .b(_T_292)
    );
    wire [2:0] _T_294;
    BITS #(.width(65), .high(31), .low(29)) bits_3077 (
        .y(_T_294),
        .in(in_bits_in1)
    );
    wire [2:0] _T_295;
    BITWISENOT #(.width(3)) bitwisenot_3078 (
        .y(_T_295),
        .in(_T_294)
    );
    wire _T_297;
    wire [2:0] _WTEMP_426;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_3079 (
        .y(_WTEMP_426),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(3)) u_eq_3080 (
        .y(_T_297),
        .a(_T_295),
        .b(_WTEMP_426)
    );
    wire [2:0] _T_298;
    BITS #(.width(65), .high(31), .low(29)) bits_3081 (
        .y(_T_298),
        .in(in_bits_in2)
    );
    wire [2:0] _T_299;
    BITWISENOT #(.width(3)) bitwisenot_3082 (
        .y(_T_299),
        .in(_T_298)
    );
    wire _T_301;
    wire [2:0] _WTEMP_427;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_3083 (
        .y(_WTEMP_427),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(3)) u_eq_3084 (
        .y(_T_301),
        .a(_T_299),
        .b(_WTEMP_427)
    );
    wire [2:0] _T_302;
    BITS #(.width(65), .high(31), .low(29)) bits_3085 (
        .y(_T_302),
        .in(in_bits_in1)
    );
    wire [2:0] _T_303;
    BITWISENOT #(.width(3)) bitwisenot_3086 (
        .y(_T_303),
        .in(_T_302)
    );
    wire _T_305;
    wire [2:0] _WTEMP_428;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_3087 (
        .y(_WTEMP_428),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(3)) u_eq_3088 (
        .y(_T_305),
        .a(_T_303),
        .b(_WTEMP_428)
    );
    wire _T_306;
    BITS #(.width(65), .high(22), .low(22)) bits_3089 (
        .y(_T_306),
        .in(in_bits_in1)
    );
    wire _T_308;
    EQ_UNSIGNED #(.width(1)) u_eq_3090 (
        .y(_T_308),
        .a(_T_306),
        .b(1'h0)
    );
    wire _T_309;
    BITWISEAND #(.width(1)) bitwiseand_3091 (
        .y(_T_309),
        .a(_T_305),
        .b(_T_308)
    );
    wire [2:0] _T_310;
    BITS #(.width(65), .high(31), .low(29)) bits_3092 (
        .y(_T_310),
        .in(in_bits_in2)
    );
    wire [2:0] _T_311;
    BITWISENOT #(.width(3)) bitwisenot_3093 (
        .y(_T_311),
        .in(_T_310)
    );
    wire _T_313;
    wire [2:0] _WTEMP_429;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_3094 (
        .y(_WTEMP_429),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(3)) u_eq_3095 (
        .y(_T_313),
        .a(_T_311),
        .b(_WTEMP_429)
    );
    wire _T_314;
    BITS #(.width(65), .high(22), .low(22)) bits_3096 (
        .y(_T_314),
        .in(in_bits_in2)
    );
    wire _T_316;
    EQ_UNSIGNED #(.width(1)) u_eq_3097 (
        .y(_T_316),
        .a(_T_314),
        .b(1'h0)
    );
    wire _T_317;
    BITWISEAND #(.width(1)) bitwiseand_3098 (
        .y(_T_317),
        .a(_T_313),
        .b(_T_316)
    );
    wire _T_318;
    BITWISEOR #(.width(1)) bitwiseor_3099 (
        .y(_T_318),
        .a(_T_309),
        .b(_T_317)
    );
    wire _T_319;
    BITWISEAND #(.width(1)) bitwiseand_3100 (
        .y(_T_319),
        .a(_T_297),
        .b(_T_301)
    );
    wire _T_320;
    BITWISEOR #(.width(1)) bitwiseor_3101 (
        .y(_T_320),
        .a(_T_318),
        .b(_T_319)
    );
    wire [65:0] _T_323;
    assign _T_323 = 66'hE0080000E0400000;
    wire [64:0] _T_324;
    assign _T_324 = 65'hE0080000E0400000;
    wire _T_325;
    BITS #(.width(3), .high(0), .low(0)) bits_3102 (
        .y(_T_325),
        .in(in_bits_rm)
    );
    wire _T_326;
    NEQ_UNSIGNED #(.width(1)) u_neq_3103 (
        .y(_T_326),
        .a(_T_325),
        .b(io_lt)
    );
    wire _T_328;
    EQ_UNSIGNED #(.width(1)) u_eq_3104 (
        .y(_T_328),
        .a(_T_297),
        .b(1'h0)
    );
    wire _T_329;
    BITWISEAND #(.width(1)) bitwiseand_3105 (
        .y(_T_329),
        .a(_T_326),
        .b(_T_328)
    );
    wire _T_330;
    BITWISEOR #(.width(1)) bitwiseor_3106 (
        .y(_T_330),
        .a(_T_301),
        .b(_T_329)
    );
    wire [2:0] _T_331;
    BITS #(.width(65), .high(63), .low(61)) bits_3107 (
        .y(_T_331),
        .in(in_bits_in1)
    );
    wire [2:0] _T_332;
    BITWISENOT #(.width(3)) bitwisenot_3108 (
        .y(_T_332),
        .in(_T_331)
    );
    wire _T_334;
    wire [2:0] _WTEMP_430;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_3109 (
        .y(_WTEMP_430),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(3)) u_eq_3110 (
        .y(_T_334),
        .a(_T_332),
        .b(_WTEMP_430)
    );
    wire [2:0] _T_335;
    BITS #(.width(65), .high(63), .low(61)) bits_3111 (
        .y(_T_335),
        .in(in_bits_in2)
    );
    wire [2:0] _T_336;
    BITWISENOT #(.width(3)) bitwisenot_3112 (
        .y(_T_336),
        .in(_T_335)
    );
    wire _T_338;
    wire [2:0] _WTEMP_431;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_3113 (
        .y(_WTEMP_431),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(3)) u_eq_3114 (
        .y(_T_338),
        .a(_T_336),
        .b(_WTEMP_431)
    );
    wire [2:0] _T_339;
    BITS #(.width(65), .high(63), .low(61)) bits_3115 (
        .y(_T_339),
        .in(in_bits_in1)
    );
    wire [2:0] _T_340;
    BITWISENOT #(.width(3)) bitwisenot_3116 (
        .y(_T_340),
        .in(_T_339)
    );
    wire _T_342;
    wire [2:0] _WTEMP_432;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_3117 (
        .y(_WTEMP_432),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(3)) u_eq_3118 (
        .y(_T_342),
        .a(_T_340),
        .b(_WTEMP_432)
    );
    wire _T_343;
    BITS #(.width(65), .high(51), .low(51)) bits_3119 (
        .y(_T_343),
        .in(in_bits_in1)
    );
    wire _T_345;
    EQ_UNSIGNED #(.width(1)) u_eq_3120 (
        .y(_T_345),
        .a(_T_343),
        .b(1'h0)
    );
    wire _T_346;
    BITWISEAND #(.width(1)) bitwiseand_3121 (
        .y(_T_346),
        .a(_T_342),
        .b(_T_345)
    );
    wire [2:0] _T_347;
    BITS #(.width(65), .high(63), .low(61)) bits_3122 (
        .y(_T_347),
        .in(in_bits_in2)
    );
    wire [2:0] _T_348;
    BITWISENOT #(.width(3)) bitwisenot_3123 (
        .y(_T_348),
        .in(_T_347)
    );
    wire _T_350;
    wire [2:0] _WTEMP_433;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_3124 (
        .y(_WTEMP_433),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(3)) u_eq_3125 (
        .y(_T_350),
        .a(_T_348),
        .b(_WTEMP_433)
    );
    wire _T_351;
    BITS #(.width(65), .high(51), .low(51)) bits_3126 (
        .y(_T_351),
        .in(in_bits_in2)
    );
    wire _T_353;
    EQ_UNSIGNED #(.width(1)) u_eq_3127 (
        .y(_T_353),
        .a(_T_351),
        .b(1'h0)
    );
    wire _T_354;
    BITWISEAND #(.width(1)) bitwiseand_3128 (
        .y(_T_354),
        .a(_T_350),
        .b(_T_353)
    );
    wire _T_355;
    BITWISEOR #(.width(1)) bitwiseor_3129 (
        .y(_T_355),
        .a(_T_346),
        .b(_T_354)
    );
    wire _T_356;
    BITWISEAND #(.width(1)) bitwiseand_3130 (
        .y(_T_356),
        .a(_T_334),
        .b(_T_338)
    );
    wire _T_357;
    BITWISEOR #(.width(1)) bitwiseor_3131 (
        .y(_T_357),
        .a(_T_355),
        .b(_T_356)
    );
    wire _T_359;
    BITS #(.width(3), .high(0), .low(0)) bits_3132 (
        .y(_T_359),
        .in(in_bits_rm)
    );
    wire _T_360;
    NEQ_UNSIGNED #(.width(1)) u_neq_3133 (
        .y(_T_360),
        .a(_T_359),
        .b(io_lt)
    );
    wire _T_362;
    EQ_UNSIGNED #(.width(1)) u_eq_3134 (
        .y(_T_362),
        .a(_T_334),
        .b(1'h0)
    );
    wire _T_363;
    BITWISEAND #(.width(1)) bitwiseand_3135 (
        .y(_T_363),
        .a(_T_360),
        .b(_T_362)
    );
    wire _T_364;
    BITWISEOR #(.width(1)) bitwiseor_3136 (
        .y(_T_364),
        .a(_T_338),
        .b(_T_363)
    );
    wire _T_365;
    MUX_UNSIGNED #(.width(1)) u_mux_3137 (
        .y(_T_365),
        .sel(in_bits_single),
        .a(_T_330),
        .b(_T_364)
    );
    wire _T_366;
    MUX_UNSIGNED #(.width(1)) u_mux_3138 (
        .y(_T_366),
        .sel(in_bits_single),
        .a(_T_318),
        .b(_T_355)
    );
    wire _T_367;
    MUX_UNSIGNED #(.width(1)) u_mux_3139 (
        .y(_T_367),
        .sel(in_bits_single),
        .a(_T_320),
        .b(_T_357)
    );
    wire [64:0] _T_368;
    MUX_UNSIGNED #(.width(65)) u_mux_3140 (
        .y(_T_368),
        .sel(in_bits_single),
        .a(_T_324),
        .b(65'hE008000000000000)
    );
    wire [4:0] _T_369;
    SHL_UNSIGNED #(.width(1), .n(4)) u_shl_3141 (
        .y(_T_369),
        .in(_T_366)
    );
    wire [64:0] _T_370;
    MUX_UNSIGNED #(.width(65)) u_mux_3142 (
        .y(_T_370),
        .sel(_T_365),
        .a(in_bits_in1),
        .b(in_bits_in2)
    );
    wire [64:0] _T_371;
    MUX_UNSIGNED #(.width(65)) u_mux_3143 (
        .y(_T_371),
        .sel(_T_367),
        .a(_T_368),
        .b(_T_370)
    );
    wire [4:0] _T_374;
    wire [4:0] _WTEMP_434;
    PAD_UNSIGNED #(.width(3), .n(5)) u_pad_3144 (
        .y(_WTEMP_434),
        .in(3'h4)
    );
    BITWISEAND #(.width(5)) bitwiseand_3145 (
        .y(_T_374),
        .a(in_bits_cmd),
        .b(_WTEMP_434)
    );
    wire _T_375;
    wire [4:0] _WTEMP_435;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_3146 (
        .y(_WTEMP_435),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(5)) u_eq_3147 (
        .y(_T_375),
        .a(_WTEMP_435),
        .b(_T_374)
    );
    wire _RecFNToRecFN__clock;
    wire _RecFNToRecFN__reset;
    wire [64:0] _RecFNToRecFN__io_in;
    wire [1:0] _RecFNToRecFN__io_roundingMode;
    wire [32:0] _RecFNToRecFN__io_out;
    wire [4:0] _RecFNToRecFN__io_exceptionFlags;
    RecFNToRecFN RecFNToRecFN (
        .clock(_RecFNToRecFN__clock),
        .reset(_RecFNToRecFN__reset),
        .io_in(_RecFNToRecFN__io_in),
        .io_roundingMode(_RecFNToRecFN__io_roundingMode),
        .io_out(_RecFNToRecFN__io_out),
        .io_exceptionFlags(_RecFNToRecFN__io_exceptionFlags)
    );
    wire _RecFNToRecFN_1__clock;
    wire _RecFNToRecFN_1__reset;
    wire [32:0] _RecFNToRecFN_1__io_in;
    wire [1:0] _RecFNToRecFN_1__io_roundingMode;
    wire [64:0] _RecFNToRecFN_1__io_out;
    wire [4:0] _RecFNToRecFN_1__io_exceptionFlags;
    RecFNToRecFN_1 RecFNToRecFN_1 (
        .clock(_RecFNToRecFN_1__clock),
        .reset(_RecFNToRecFN_1__reset),
        .io_in(_RecFNToRecFN_1__io_in),
        .io_roundingMode(_RecFNToRecFN_1__io_roundingMode),
        .io_out(_RecFNToRecFN_1__io_out),
        .io_exceptionFlags(_RecFNToRecFN_1__io_exceptionFlags)
    );
    wire [31:0] _T_376;
    SHR_UNSIGNED #(.width(65), .n(33)) u_shr_3435 (
        .y(_T_376),
        .in(_RecFNToRecFN_1__io_out)
    );
    wire [64:0] _T_377;
    CAT #(.width_a(32), .width_b(33)) cat_3436 (
        .y(_T_377),
        .a(_T_376),
        .b(_RecFNToRecFN__io_out)
    );
    wire [64:0] _node_30;
    MUX_UNSIGNED #(.width(65)) u_mux_3437 (
        .y(_node_30),
        .sel(_T_293),
        .a(_T_371),
        .b(fsgnj)
    );
    wire [4:0] _node_31;
    wire [4:0] _WTEMP_474;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_3438 (
        .y(_WTEMP_474),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(5)) u_mux_3439 (
        .y(_node_31),
        .sel(_T_293),
        .a(_T_369),
        .b(_WTEMP_474)
    );
    wire _T_379;
    EQ_UNSIGNED #(.width(1)) u_eq_3440 (
        .y(_T_379),
        .a(in_bits_single),
        .b(1'h0)
    );
    wire [64:0] _node_32;
    MUX_UNSIGNED #(.width(65)) u_mux_3441 (
        .y(_node_32),
        .sel(in_bits_single),
        .a(_T_377),
        .b(_node_30)
    );
    wire [4:0] _node_33;
    MUX_UNSIGNED #(.width(5)) u_mux_3442 (
        .y(_node_33),
        .sel(in_bits_single),
        .a(_RecFNToRecFN__io_exceptionFlags),
        .b(_node_31)
    );
    wire [64:0] _node_34;
    MUX_UNSIGNED #(.width(65)) u_mux_3443 (
        .y(_node_34),
        .sel(_T_379),
        .a(_RecFNToRecFN_1__io_out),
        .b(_node_32)
    );
    wire [64:0] _node_35;
    MUX_UNSIGNED #(.width(65)) u_mux_3444 (
        .y(_node_35),
        .sel(_T_293),
        .a(_T_371),
        .b(fsgnj)
    );
    wire [4:0] _node_36;
    MUX_UNSIGNED #(.width(5)) u_mux_3445 (
        .y(_node_36),
        .sel(_T_379),
        .a(_RecFNToRecFN_1__io_exceptionFlags),
        .b(_node_33)
    );
    wire [4:0] _node_37;
    wire [4:0] _WTEMP_475;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_3446 (
        .y(_WTEMP_475),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(5)) u_mux_3447 (
        .y(_node_37),
        .sel(_T_293),
        .a(_T_369),
        .b(_WTEMP_475)
    );
    wire __T_382__q;
    wire __T_382__d;
    DFF_POSCLK #(.width(1)) _T_382 (
        .q(__T_382__q),
        .d(__T_382__d),
        .clk(clock)
    );
    wire _WTEMP_476;
    MUX_UNSIGNED #(.width(1)) u_mux_3448 (
        .y(__T_382__d),
        .sel(reset),
        .a(1'h0),
        .b(_WTEMP_476)
    );
    wire [64:0] __T_386_data__q;
    wire [64:0] __T_386_data__d;
    DFF_POSCLK #(.width(65)) _T_386_data (
        .q(__T_386_data__q),
        .d(__T_386_data__d),
        .clk(clock)
    );
    wire [4:0] __T_386_exc__q;
    wire [4:0] __T_386_exc__d;
    DFF_POSCLK #(.width(5)) _T_386_exc (
        .q(__T_386_exc__q),
        .d(__T_386_exc__d),
        .clk(clock)
    );
    wire _T_398_valid;
    wire [64:0] _T_398_bits_data;
    wire [4:0] _T_398_bits_exc;
    assign _RecFNToRecFN__clock = clock;
    assign _RecFNToRecFN__io_in = in_bits_in1;
    BITS #(.width(3), .high(1), .low(0)) bits_3449 (
        .y(_RecFNToRecFN__io_roundingMode),
        .in(in_bits_rm)
    );
    assign _RecFNToRecFN__reset = reset;
    assign _RecFNToRecFN_1__clock = clock;
    BITS #(.width(65), .high(32), .low(0)) bits_3450 (
        .y(_RecFNToRecFN_1__io_in),
        .in(in_bits_in1)
    );
    BITS #(.width(3), .high(1), .low(0)) bits_3451 (
        .y(_RecFNToRecFN_1__io_roundingMode),
        .in(in_bits_rm)
    );
    assign _RecFNToRecFN_1__reset = reset;
    assign _WTEMP_423 = io_in_valid;
    MUX_UNSIGNED #(.width(5)) u_mux_3452 (
        .y(__T_157_cmd__d),
        .sel(io_in_valid),
        .a(io_in_bits_cmd),
        .b(__T_157_cmd__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_3453 (
        .y(__T_157_div__d),
        .sel(io_in_valid),
        .a(io_in_bits_div),
        .b(__T_157_div__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_3454 (
        .y(__T_157_fastpipe__d),
        .sel(io_in_valid),
        .a(io_in_bits_fastpipe),
        .b(__T_157_fastpipe__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_3455 (
        .y(__T_157_fma__d),
        .sel(io_in_valid),
        .a(io_in_bits_fma),
        .b(__T_157_fma__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_3456 (
        .y(__T_157_fromint__d),
        .sel(io_in_valid),
        .a(io_in_bits_fromint),
        .b(__T_157_fromint__q)
    );
    MUX_UNSIGNED #(.width(65)) u_mux_3457 (
        .y(__T_157_in1__d),
        .sel(io_in_valid),
        .a(io_in_bits_in1),
        .b(__T_157_in1__q)
    );
    MUX_UNSIGNED #(.width(65)) u_mux_3458 (
        .y(__T_157_in2__d),
        .sel(io_in_valid),
        .a(io_in_bits_in2),
        .b(__T_157_in2__q)
    );
    MUX_UNSIGNED #(.width(65)) u_mux_3459 (
        .y(__T_157_in3__d),
        .sel(io_in_valid),
        .a(io_in_bits_in3),
        .b(__T_157_in3__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_3460 (
        .y(__T_157_ldst__d),
        .sel(io_in_valid),
        .a(io_in_bits_ldst),
        .b(__T_157_ldst__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_3461 (
        .y(__T_157_ren1__d),
        .sel(io_in_valid),
        .a(io_in_bits_ren1),
        .b(__T_157_ren1__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_3462 (
        .y(__T_157_ren2__d),
        .sel(io_in_valid),
        .a(io_in_bits_ren2),
        .b(__T_157_ren2__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_3463 (
        .y(__T_157_ren3__d),
        .sel(io_in_valid),
        .a(io_in_bits_ren3),
        .b(__T_157_ren3__q)
    );
    MUX_UNSIGNED #(.width(3)) u_mux_3464 (
        .y(__T_157_rm__d),
        .sel(io_in_valid),
        .a(io_in_bits_rm),
        .b(__T_157_rm__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_3465 (
        .y(__T_157_single__d),
        .sel(io_in_valid),
        .a(io_in_bits_single),
        .b(__T_157_single__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_3466 (
        .y(__T_157_sqrt__d),
        .sel(io_in_valid),
        .a(io_in_bits_sqrt),
        .b(__T_157_sqrt__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_3467 (
        .y(__T_157_swap12__d),
        .sel(io_in_valid),
        .a(io_in_bits_swap12),
        .b(__T_157_swap12__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_3468 (
        .y(__T_157_swap23__d),
        .sel(io_in_valid),
        .a(io_in_bits_swap23),
        .b(__T_157_swap23__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_3469 (
        .y(__T_157_toint__d),
        .sel(io_in_valid),
        .a(io_in_bits_toint),
        .b(__T_157_toint__q)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_3470 (
        .y(__T_157_typ__d),
        .sel(io_in_valid),
        .a(io_in_bits_typ),
        .b(__T_157_typ__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_3471 (
        .y(__T_157_wen__d),
        .sel(io_in_valid),
        .a(io_in_bits_wen),
        .b(__T_157_wen__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_3472 (
        .y(__T_157_wflags__d),
        .sel(io_in_valid),
        .a(io_in_bits_wflags),
        .b(__T_157_wflags__q)
    );
    assign _WTEMP_476 = in_valid;
    MUX_UNSIGNED #(.width(65)) u_mux_3473 (
        .y(__T_386_data__d),
        .sel(in_valid),
        .a(mux_data),
        .b(__T_386_data__q)
    );
    MUX_UNSIGNED #(.width(5)) u_mux_3474 (
        .y(__T_386_exc__d),
        .sel(in_valid),
        .a(mux_exc),
        .b(__T_386_exc__q)
    );
    assign _T_398_bits_data = __T_386_data__q;
    assign _T_398_bits_exc = __T_386_exc__q;
    assign _T_398_valid = __T_382__q;
    assign in_bits_cmd = __T_157_cmd__q;
    assign in_bits_div = __T_157_div__q;
    assign in_bits_fastpipe = __T_157_fastpipe__q;
    assign in_bits_fma = __T_157_fma__q;
    assign in_bits_fromint = __T_157_fromint__q;
    assign in_bits_in1 = __T_157_in1__q;
    assign in_bits_in2 = __T_157_in2__q;
    assign in_bits_in3 = __T_157_in3__q;
    assign in_bits_ldst = __T_157_ldst__q;
    assign in_bits_ren1 = __T_157_ren1__q;
    assign in_bits_ren2 = __T_157_ren2__q;
    assign in_bits_ren3 = __T_157_ren3__q;
    assign in_bits_rm = __T_157_rm__q;
    assign in_bits_single = __T_157_single__q;
    assign in_bits_sqrt = __T_157_sqrt__q;
    assign in_bits_swap12 = __T_157_swap12__q;
    assign in_bits_swap23 = __T_157_swap23__q;
    assign in_bits_toint = __T_157_toint__q;
    assign in_bits_typ = __T_157_typ__q;
    assign in_bits_wen = __T_157_wen__q;
    assign in_bits_wflags = __T_157_wflags__q;
    assign in_valid = __T_134__q;
    assign io_out_bits_data = _T_398_bits_data;
    assign io_out_bits_exc = _T_398_bits_exc;
    assign io_out_valid = _T_398_valid;
    MUX_UNSIGNED #(.width(65)) u_mux_3475 (
        .y(mux_data),
        .sel(_T_375),
        .a(_node_34),
        .b(_node_35)
    );
    MUX_UNSIGNED #(.width(5)) u_mux_3476 (
        .y(mux_exc),
        .sel(_T_375),
        .a(_node_36),
        .b(_node_37)
    );
endmodule //FPToFP
module RecFNToRecFN(
    input clock,
    input reset,
    input [64:0] io_in,
    input [1:0] io_roundingMode,
    output [32:0] io_out,
    output [4:0] io_exceptionFlags
);
    wire [11:0] _T_10;
    BITS #(.width(65), .high(63), .low(52)) bits_3148 (
        .y(_T_10),
        .in(io_in)
    );
    wire [2:0] _T_11;
    BITS #(.width(12), .high(11), .low(9)) bits_3149 (
        .y(_T_11),
        .in(_T_10)
    );
    wire _T_13;
    wire [2:0] _WTEMP_436;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_3150 (
        .y(_WTEMP_436),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(3)) u_eq_3151 (
        .y(_T_13),
        .a(_T_11),
        .b(_WTEMP_436)
    );
    wire [1:0] _T_14;
    BITS #(.width(12), .high(11), .low(10)) bits_3152 (
        .y(_T_14),
        .in(_T_10)
    );
    wire _T_16;
    EQ_UNSIGNED #(.width(2)) u_eq_3153 (
        .y(_T_16),
        .a(_T_14),
        .b(2'h3)
    );
    wire _T_24_sign;
    wire _T_24_isNaN;
    wire _T_24_isInf;
    wire _T_24_isZero;
    wire [12:0] _T_24_sExp;
    wire [55:0] _T_24_sig;
    wire _T_31;
    BITS #(.width(65), .high(64), .low(64)) bits_3154 (
        .y(_T_31),
        .in(io_in)
    );
    wire _T_32;
    BITS #(.width(12), .high(9), .low(9)) bits_3155 (
        .y(_T_32),
        .in(_T_10)
    );
    wire _T_33;
    BITWISEAND #(.width(1)) bitwiseand_3156 (
        .y(_T_33),
        .a(_T_16),
        .b(_T_32)
    );
    wire _T_34;
    BITS #(.width(12), .high(9), .low(9)) bits_3157 (
        .y(_T_34),
        .in(_T_10)
    );
    wire _T_36;
    EQ_UNSIGNED #(.width(1)) u_eq_3158 (
        .y(_T_36),
        .a(_T_34),
        .b(1'h0)
    );
    wire _T_37;
    BITWISEAND #(.width(1)) bitwiseand_3159 (
        .y(_T_37),
        .a(_T_16),
        .b(_T_36)
    );
    wire [12:0] _T_38;
    CVT_UNSIGNED #(.width(12)) u_cvt_3160 (
        .y(_T_38),
        .in(_T_10)
    );
    wire _T_41;
    EQ_UNSIGNED #(.width(1)) u_eq_3161 (
        .y(_T_41),
        .a(_T_13),
        .b(1'h0)
    );
    wire [51:0] _T_42;
    BITS #(.width(65), .high(51), .low(0)) bits_3162 (
        .y(_T_42),
        .in(io_in)
    );
    wire [53:0] _T_44;
    CAT #(.width_a(52), .width_b(2)) cat_3163 (
        .y(_T_44),
        .a(_T_42),
        .b(2'h0)
    );
    wire [1:0] _T_45;
    CAT #(.width_a(1), .width_b(1)) cat_3164 (
        .y(_T_45),
        .a(1'h0),
        .b(_T_41)
    );
    wire [55:0] _T_46;
    CAT #(.width_a(2), .width_b(54)) cat_3165 (
        .y(_T_46),
        .a(_T_45),
        .b(_T_44)
    );
    wire [13:0] _T_48;
    wire [12:0] _WTEMP_437;
    PAD_SIGNED #(.width(12), .n(13)) s_pad_3166 (
        .y(_WTEMP_437),
        .in(-12'sh700)
    );
    ADD_SIGNED #(.width(13)) s_add_3167 (
        .y(_T_48),
        .a(_T_24_sExp),
        .b(_WTEMP_437)
    );
    wire outRawFloat_sign;
    wire outRawFloat_isNaN;
    wire outRawFloat_isInf;
    wire outRawFloat_isZero;
    wire [9:0] outRawFloat_sExp;
    wire [26:0] outRawFloat_sig;
    wire _T_63;
    wire [13:0] _WTEMP_438;
    PAD_SIGNED #(.width(1), .n(14)) s_pad_3168 (
        .y(_WTEMP_438),
        .in(1'sh0)
    );
    LT_SIGNED #(.width(14)) s_lt_3169 (
        .y(_T_63),
        .a(_T_48),
        .b(_WTEMP_438)
    );
    wire [3:0] _T_64;
    BITS #(.width(14), .high(12), .low(9)) bits_3170 (
        .y(_T_64),
        .in(_T_48)
    );
    wire _T_66;
    wire [3:0] _WTEMP_439;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_3171 (
        .y(_WTEMP_439),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_3172 (
        .y(_T_66),
        .a(_T_64),
        .b(_WTEMP_439)
    );
    wire [6:0] _T_71;
    assign _T_71 = 7'h7F;
    wire [8:0] _T_73;
    assign _T_73 = 9'h1FC;
    wire [8:0] _T_74;
    BITS #(.width(14), .high(8), .low(0)) bits_3173 (
        .y(_T_74),
        .in(_T_48)
    );
    wire [8:0] _T_75;
    MUX_UNSIGNED #(.width(9)) u_mux_3174 (
        .y(_T_75),
        .sel(_T_66),
        .a(_T_73),
        .b(_T_74)
    );
    wire [9:0] _T_76;
    CAT #(.width_a(1), .width_b(9)) cat_3175 (
        .y(_T_76),
        .a(_T_63),
        .b(_T_75)
    );
    wire [9:0] _T_77;
    ASSINT #(.width(10)) assint_3176 (
        .y(_T_77),
        .in(_T_76)
    );
    wire [25:0] _T_78;
    BITS #(.width(56), .high(55), .low(30)) bits_3177 (
        .y(_T_78),
        .in(_T_24_sig)
    );
    wire [29:0] _T_79;
    BITS #(.width(56), .high(29), .low(0)) bits_3178 (
        .y(_T_79),
        .in(_T_24_sig)
    );
    wire _T_81;
    wire [29:0] _WTEMP_440;
    PAD_UNSIGNED #(.width(1), .n(30)) u_pad_3179 (
        .y(_WTEMP_440),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(30)) u_neq_3180 (
        .y(_T_81),
        .a(_T_79),
        .b(_WTEMP_440)
    );
    wire [26:0] _T_82;
    CAT #(.width_a(26), .width_b(1)) cat_3181 (
        .y(_T_82),
        .a(_T_78),
        .b(_T_81)
    );
    wire _T_83;
    BITS #(.width(27), .high(24), .low(24)) bits_3182 (
        .y(_T_83),
        .in(outRawFloat_sig)
    );
    wire _T_85;
    EQ_UNSIGNED #(.width(1)) u_eq_3183 (
        .y(_T_85),
        .a(_T_83),
        .b(1'h0)
    );
    wire invalidExc;
    BITWISEAND #(.width(1)) bitwiseand_3184 (
        .y(invalidExc),
        .a(outRawFloat_isNaN),
        .b(_T_85)
    );
    wire _RoundRawFNToRecFN__clock;
    wire _RoundRawFNToRecFN__reset;
    wire _RoundRawFNToRecFN__io_invalidExc;
    wire _RoundRawFNToRecFN__io_infiniteExc;
    wire _RoundRawFNToRecFN__io_in_sign;
    wire _RoundRawFNToRecFN__io_in_isNaN;
    wire _RoundRawFNToRecFN__io_in_isInf;
    wire _RoundRawFNToRecFN__io_in_isZero;
    wire [9:0] _RoundRawFNToRecFN__io_in_sExp;
    wire [26:0] _RoundRawFNToRecFN__io_in_sig;
    wire [1:0] _RoundRawFNToRecFN__io_roundingMode;
    wire [32:0] _RoundRawFNToRecFN__io_out;
    wire [4:0] _RoundRawFNToRecFN__io_exceptionFlags;
    RoundRawFNToRecFN RoundRawFNToRecFN (
        .clock(_RoundRawFNToRecFN__clock),
        .reset(_RoundRawFNToRecFN__reset),
        .io_invalidExc(_RoundRawFNToRecFN__io_invalidExc),
        .io_infiniteExc(_RoundRawFNToRecFN__io_infiniteExc),
        .io_in_sign(_RoundRawFNToRecFN__io_in_sign),
        .io_in_isNaN(_RoundRawFNToRecFN__io_in_isNaN),
        .io_in_isInf(_RoundRawFNToRecFN__io_in_isInf),
        .io_in_isZero(_RoundRawFNToRecFN__io_in_isZero),
        .io_in_sExp(_RoundRawFNToRecFN__io_in_sExp),
        .io_in_sig(_RoundRawFNToRecFN__io_in_sig),
        .io_roundingMode(_RoundRawFNToRecFN__io_roundingMode),
        .io_out(_RoundRawFNToRecFN__io_out),
        .io_exceptionFlags(_RoundRawFNToRecFN__io_exceptionFlags)
    );
    assign _RoundRawFNToRecFN__clock = clock;
    assign _RoundRawFNToRecFN__io_in_isInf = outRawFloat_isInf;
    assign _RoundRawFNToRecFN__io_in_isNaN = outRawFloat_isNaN;
    assign _RoundRawFNToRecFN__io_in_isZero = outRawFloat_isZero;
    assign _RoundRawFNToRecFN__io_in_sExp = outRawFloat_sExp;
    assign _RoundRawFNToRecFN__io_in_sig = outRawFloat_sig;
    assign _RoundRawFNToRecFN__io_in_sign = outRawFloat_sign;
    assign _RoundRawFNToRecFN__io_infiniteExc = 1'h0;
    assign _RoundRawFNToRecFN__io_invalidExc = invalidExc;
    assign _RoundRawFNToRecFN__io_roundingMode = io_roundingMode;
    assign _RoundRawFNToRecFN__reset = reset;
    assign _T_24_isInf = _T_37;
    assign _T_24_isNaN = _T_33;
    assign _T_24_isZero = _T_13;
    assign _T_24_sExp = _T_38;
    assign _T_24_sig = _T_46;
    assign _T_24_sign = _T_31;
    assign io_exceptionFlags = _RoundRawFNToRecFN__io_exceptionFlags;
    assign io_out = _RoundRawFNToRecFN__io_out;
    assign outRawFloat_isInf = _T_24_isInf;
    assign outRawFloat_isNaN = _T_24_isNaN;
    assign outRawFloat_isZero = _T_24_isZero;
    assign outRawFloat_sExp = _T_77;
    assign outRawFloat_sig = _T_82;
    assign outRawFloat_sign = _T_24_sign;
endmodule //RecFNToRecFN
module ADD_SIGNED(y, a, b);
    parameter width = 4;
    output [width:0] y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = $signed(a) + $signed(b);
endmodule // ADD_SIGNED
module RoundRawFNToRecFN(
    input clock,
    input reset,
    input io_invalidExc,
    input io_infiniteExc,
    input io_in_sign,
    input io_in_isNaN,
    input io_in_isInf,
    input io_in_isZero,
    input [9:0] io_in_sExp,
    input [26:0] io_in_sig,
    input [1:0] io_roundingMode,
    output [32:0] io_out,
    output [4:0] io_exceptionFlags
);
    wire roundingMode_nearest_even;
    EQ_UNSIGNED #(.width(2)) u_eq_3185 (
        .y(roundingMode_nearest_even),
        .a(io_roundingMode),
        .b(2'h0)
    );
    wire roundingMode_minMag;
    EQ_UNSIGNED #(.width(2)) u_eq_3186 (
        .y(roundingMode_minMag),
        .a(io_roundingMode),
        .b(2'h1)
    );
    wire roundingMode_min;
    EQ_UNSIGNED #(.width(2)) u_eq_3187 (
        .y(roundingMode_min),
        .a(io_roundingMode),
        .b(2'h2)
    );
    wire roundingMode_max;
    EQ_UNSIGNED #(.width(2)) u_eq_3188 (
        .y(roundingMode_max),
        .a(io_roundingMode),
        .b(2'h3)
    );
    wire _T_26;
    BITWISEAND #(.width(1)) bitwiseand_3189 (
        .y(_T_26),
        .a(roundingMode_min),
        .b(io_in_sign)
    );
    wire _T_28;
    EQ_UNSIGNED #(.width(1)) u_eq_3190 (
        .y(_T_28),
        .a(io_in_sign),
        .b(1'h0)
    );
    wire _T_29;
    BITWISEAND #(.width(1)) bitwiseand_3191 (
        .y(_T_29),
        .a(roundingMode_max),
        .b(_T_28)
    );
    wire roundMagUp;
    BITWISEOR #(.width(1)) bitwiseor_3192 (
        .y(roundMagUp),
        .a(_T_26),
        .b(_T_29)
    );
    wire doShiftSigDown1;
    BITS #(.width(27), .high(26), .low(26)) bits_3193 (
        .y(doShiftSigDown1),
        .in(io_in_sig)
    );
    wire isNegExp;
    wire [9:0] _WTEMP_441;
    PAD_SIGNED #(.width(1), .n(10)) s_pad_3194 (
        .y(_WTEMP_441),
        .in(1'sh0)
    );
    LT_SIGNED #(.width(10)) s_lt_3195 (
        .y(isNegExp),
        .a(io_in_sExp),
        .b(_WTEMP_441)
    );
    wire _T_31;
    BITS #(.width(1), .high(0), .low(0)) bits_3196 (
        .y(_T_31),
        .in(isNegExp)
    );
    wire [24:0] _T_34;
    MUX_UNSIGNED #(.width(25)) u_mux_3197 (
        .y(_T_34),
        .sel(_T_31),
        .a(25'h1FFFFFF),
        .b(25'h0)
    );
    wire [8:0] _T_35;
    BITS #(.width(10), .high(8), .low(0)) bits_3198 (
        .y(_T_35),
        .in(io_in_sExp)
    );
    wire [8:0] _T_36;
    BITWISENOT #(.width(9)) bitwisenot_3199 (
        .y(_T_36),
        .in(_T_35)
    );
    wire _T_37;
    BITS #(.width(9), .high(8), .low(8)) bits_3200 (
        .y(_T_37),
        .in(_T_36)
    );
    wire [7:0] _T_38;
    BITS #(.width(9), .high(7), .low(0)) bits_3201 (
        .y(_T_38),
        .in(_T_36)
    );
    wire _T_39;
    BITS #(.width(8), .high(7), .low(7)) bits_3202 (
        .y(_T_39),
        .in(_T_38)
    );
    wire [6:0] _T_40;
    BITS #(.width(8), .high(6), .low(0)) bits_3203 (
        .y(_T_40),
        .in(_T_38)
    );
    wire _T_41;
    BITS #(.width(7), .high(6), .low(6)) bits_3204 (
        .y(_T_41),
        .in(_T_40)
    );
    wire [5:0] _T_42;
    BITS #(.width(7), .high(5), .low(0)) bits_3205 (
        .y(_T_42),
        .in(_T_40)
    );
    wire [64:0] _T_45;
    DSHR_SIGNED #(.width_in(65), .width_n(6)) s_dshr_3206 (
        .y(_T_45),
        .in(-65'sh10000000000000000),
        .n(_T_42)
    );
    wire [21:0] _T_46;
    BITS #(.width(65), .high(63), .low(42)) bits_3207 (
        .y(_T_46),
        .in(_T_45)
    );
    wire [15:0] _T_47;
    BITS #(.width(22), .high(15), .low(0)) bits_3208 (
        .y(_T_47),
        .in(_T_46)
    );
    wire [15:0] _T_50;
    assign _T_50 = 16'hFF00;
    wire [15:0] _T_51;
    assign _T_51 = 16'hFF;
    wire [7:0] _T_52;
    SHR_UNSIGNED #(.width(16), .n(8)) u_shr_3209 (
        .y(_T_52),
        .in(_T_47)
    );
    wire [15:0] _T_53;
    wire [15:0] _WTEMP_442;
    PAD_UNSIGNED #(.width(8), .n(16)) u_pad_3210 (
        .y(_WTEMP_442),
        .in(_T_52)
    );
    BITWISEAND #(.width(16)) bitwiseand_3211 (
        .y(_T_53),
        .a(_WTEMP_442),
        .b(_T_51)
    );
    wire [7:0] _T_54;
    BITS #(.width(16), .high(7), .low(0)) bits_3212 (
        .y(_T_54),
        .in(_T_47)
    );
    wire [15:0] _T_55;
    SHL_UNSIGNED #(.width(8), .n(8)) u_shl_3213 (
        .y(_T_55),
        .in(_T_54)
    );
    wire [15:0] _T_56;
    assign _T_56 = 16'hFF00;
    wire [15:0] _T_57;
    BITWISEAND #(.width(16)) bitwiseand_3214 (
        .y(_T_57),
        .a(_T_55),
        .b(_T_56)
    );
    wire [15:0] _T_58;
    BITWISEOR #(.width(16)) bitwiseor_3215 (
        .y(_T_58),
        .a(_T_53),
        .b(_T_57)
    );
    wire [11:0] _T_59;
    assign _T_59 = 12'hFF;
    wire [15:0] _T_60;
    assign _T_60 = 16'hFF0;
    wire [15:0] _T_61;
    assign _T_61 = 16'hF0F;
    wire [11:0] _T_62;
    SHR_UNSIGNED #(.width(16), .n(4)) u_shr_3216 (
        .y(_T_62),
        .in(_T_58)
    );
    wire [15:0] _T_63;
    wire [15:0] _WTEMP_443;
    PAD_UNSIGNED #(.width(12), .n(16)) u_pad_3217 (
        .y(_WTEMP_443),
        .in(_T_62)
    );
    BITWISEAND #(.width(16)) bitwiseand_3218 (
        .y(_T_63),
        .a(_WTEMP_443),
        .b(_T_61)
    );
    wire [11:0] _T_64;
    BITS #(.width(16), .high(11), .low(0)) bits_3219 (
        .y(_T_64),
        .in(_T_58)
    );
    wire [15:0] _T_65;
    SHL_UNSIGNED #(.width(12), .n(4)) u_shl_3220 (
        .y(_T_65),
        .in(_T_64)
    );
    wire [15:0] _T_66;
    assign _T_66 = 16'hF0F0;
    wire [15:0] _T_67;
    BITWISEAND #(.width(16)) bitwiseand_3221 (
        .y(_T_67),
        .a(_T_65),
        .b(_T_66)
    );
    wire [15:0] _T_68;
    BITWISEOR #(.width(16)) bitwiseor_3222 (
        .y(_T_68),
        .a(_T_63),
        .b(_T_67)
    );
    wire [13:0] _T_69;
    assign _T_69 = 14'hF0F;
    wire [15:0] _T_70;
    assign _T_70 = 16'h3C3C;
    wire [15:0] _T_71;
    assign _T_71 = 16'h3333;
    wire [13:0] _T_72;
    SHR_UNSIGNED #(.width(16), .n(2)) u_shr_3223 (
        .y(_T_72),
        .in(_T_68)
    );
    wire [15:0] _T_73;
    wire [15:0] _WTEMP_444;
    PAD_UNSIGNED #(.width(14), .n(16)) u_pad_3224 (
        .y(_WTEMP_444),
        .in(_T_72)
    );
    BITWISEAND #(.width(16)) bitwiseand_3225 (
        .y(_T_73),
        .a(_WTEMP_444),
        .b(_T_71)
    );
    wire [13:0] _T_74;
    BITS #(.width(16), .high(13), .low(0)) bits_3226 (
        .y(_T_74),
        .in(_T_68)
    );
    wire [15:0] _T_75;
    SHL_UNSIGNED #(.width(14), .n(2)) u_shl_3227 (
        .y(_T_75),
        .in(_T_74)
    );
    wire [15:0] _T_76;
    assign _T_76 = 16'hCCCC;
    wire [15:0] _T_77;
    BITWISEAND #(.width(16)) bitwiseand_3228 (
        .y(_T_77),
        .a(_T_75),
        .b(_T_76)
    );
    wire [15:0] _T_78;
    BITWISEOR #(.width(16)) bitwiseor_3229 (
        .y(_T_78),
        .a(_T_73),
        .b(_T_77)
    );
    wire [14:0] _T_79;
    assign _T_79 = 15'h3333;
    wire [15:0] _T_80;
    assign _T_80 = 16'h6666;
    wire [15:0] _T_81;
    assign _T_81 = 16'h5555;
    wire [14:0] _T_82;
    SHR_UNSIGNED #(.width(16), .n(1)) u_shr_3230 (
        .y(_T_82),
        .in(_T_78)
    );
    wire [15:0] _T_83;
    wire [15:0] _WTEMP_445;
    PAD_UNSIGNED #(.width(15), .n(16)) u_pad_3231 (
        .y(_WTEMP_445),
        .in(_T_82)
    );
    BITWISEAND #(.width(16)) bitwiseand_3232 (
        .y(_T_83),
        .a(_WTEMP_445),
        .b(_T_81)
    );
    wire [14:0] _T_84;
    BITS #(.width(16), .high(14), .low(0)) bits_3233 (
        .y(_T_84),
        .in(_T_78)
    );
    wire [15:0] _T_85;
    SHL_UNSIGNED #(.width(15), .n(1)) u_shl_3234 (
        .y(_T_85),
        .in(_T_84)
    );
    wire [15:0] _T_86;
    assign _T_86 = 16'hAAAA;
    wire [15:0] _T_87;
    BITWISEAND #(.width(16)) bitwiseand_3235 (
        .y(_T_87),
        .a(_T_85),
        .b(_T_86)
    );
    wire [15:0] _T_88;
    BITWISEOR #(.width(16)) bitwiseor_3236 (
        .y(_T_88),
        .a(_T_83),
        .b(_T_87)
    );
    wire [5:0] _T_89;
    BITS #(.width(22), .high(21), .low(16)) bits_3237 (
        .y(_T_89),
        .in(_T_46)
    );
    wire [3:0] _T_90;
    BITS #(.width(6), .high(3), .low(0)) bits_3238 (
        .y(_T_90),
        .in(_T_89)
    );
    wire [1:0] _T_91;
    BITS #(.width(4), .high(1), .low(0)) bits_3239 (
        .y(_T_91),
        .in(_T_90)
    );
    wire _T_92;
    BITS #(.width(2), .high(0), .low(0)) bits_3240 (
        .y(_T_92),
        .in(_T_91)
    );
    wire _T_93;
    BITS #(.width(2), .high(1), .low(1)) bits_3241 (
        .y(_T_93),
        .in(_T_91)
    );
    wire [1:0] _T_94;
    CAT #(.width_a(1), .width_b(1)) cat_3242 (
        .y(_T_94),
        .a(_T_92),
        .b(_T_93)
    );
    wire [1:0] _T_95;
    BITS #(.width(4), .high(3), .low(2)) bits_3243 (
        .y(_T_95),
        .in(_T_90)
    );
    wire _T_96;
    BITS #(.width(2), .high(0), .low(0)) bits_3244 (
        .y(_T_96),
        .in(_T_95)
    );
    wire _T_97;
    BITS #(.width(2), .high(1), .low(1)) bits_3245 (
        .y(_T_97),
        .in(_T_95)
    );
    wire [1:0] _T_98;
    CAT #(.width_a(1), .width_b(1)) cat_3246 (
        .y(_T_98),
        .a(_T_96),
        .b(_T_97)
    );
    wire [3:0] _T_99;
    CAT #(.width_a(2), .width_b(2)) cat_3247 (
        .y(_T_99),
        .a(_T_94),
        .b(_T_98)
    );
    wire [1:0] _T_100;
    BITS #(.width(6), .high(5), .low(4)) bits_3248 (
        .y(_T_100),
        .in(_T_89)
    );
    wire _T_101;
    BITS #(.width(2), .high(0), .low(0)) bits_3249 (
        .y(_T_101),
        .in(_T_100)
    );
    wire _T_102;
    BITS #(.width(2), .high(1), .low(1)) bits_3250 (
        .y(_T_102),
        .in(_T_100)
    );
    wire [1:0] _T_103;
    CAT #(.width_a(1), .width_b(1)) cat_3251 (
        .y(_T_103),
        .a(_T_101),
        .b(_T_102)
    );
    wire [5:0] _T_104;
    CAT #(.width_a(4), .width_b(2)) cat_3252 (
        .y(_T_104),
        .a(_T_99),
        .b(_T_103)
    );
    wire [21:0] _T_105;
    CAT #(.width_a(16), .width_b(6)) cat_3253 (
        .y(_T_105),
        .a(_T_88),
        .b(_T_104)
    );
    wire [21:0] _T_106;
    BITWISENOT #(.width(22)) bitwisenot_3254 (
        .y(_T_106),
        .in(_T_105)
    );
    wire [21:0] _T_107;
    wire [21:0] _WTEMP_446;
    PAD_UNSIGNED #(.width(1), .n(22)) u_pad_3255 (
        .y(_WTEMP_446),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(22)) u_mux_3256 (
        .y(_T_107),
        .sel(_T_41),
        .a(_WTEMP_446),
        .b(_T_106)
    );
    wire [21:0] _T_108;
    BITWISENOT #(.width(22)) bitwisenot_3257 (
        .y(_T_108),
        .in(_T_107)
    );
    wire [24:0] _T_110;
    CAT #(.width_a(22), .width_b(3)) cat_3258 (
        .y(_T_110),
        .a(_T_108),
        .b(3'h7)
    );
    wire _T_111;
    BITS #(.width(7), .high(6), .low(6)) bits_3259 (
        .y(_T_111),
        .in(_T_40)
    );
    wire [5:0] _T_112;
    BITS #(.width(7), .high(5), .low(0)) bits_3260 (
        .y(_T_112),
        .in(_T_40)
    );
    wire [64:0] _T_114;
    DSHR_SIGNED #(.width_in(65), .width_n(6)) s_dshr_3261 (
        .y(_T_114),
        .in(-65'sh10000000000000000),
        .n(_T_112)
    );
    wire [2:0] _T_115;
    BITS #(.width(65), .high(2), .low(0)) bits_3262 (
        .y(_T_115),
        .in(_T_114)
    );
    wire [1:0] _T_116;
    BITS #(.width(3), .high(1), .low(0)) bits_3263 (
        .y(_T_116),
        .in(_T_115)
    );
    wire _T_117;
    BITS #(.width(2), .high(0), .low(0)) bits_3264 (
        .y(_T_117),
        .in(_T_116)
    );
    wire _T_118;
    BITS #(.width(2), .high(1), .low(1)) bits_3265 (
        .y(_T_118),
        .in(_T_116)
    );
    wire [1:0] _T_119;
    CAT #(.width_a(1), .width_b(1)) cat_3266 (
        .y(_T_119),
        .a(_T_117),
        .b(_T_118)
    );
    wire _T_120;
    BITS #(.width(3), .high(2), .low(2)) bits_3267 (
        .y(_T_120),
        .in(_T_115)
    );
    wire [2:0] _T_121;
    CAT #(.width_a(2), .width_b(1)) cat_3268 (
        .y(_T_121),
        .a(_T_119),
        .b(_T_120)
    );
    wire [2:0] _T_123;
    wire [2:0] _WTEMP_447;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_3269 (
        .y(_WTEMP_447),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(3)) u_mux_3270 (
        .y(_T_123),
        .sel(_T_111),
        .a(_T_121),
        .b(_WTEMP_447)
    );
    wire [24:0] _T_124;
    wire [24:0] _WTEMP_448;
    PAD_UNSIGNED #(.width(3), .n(25)) u_pad_3271 (
        .y(_WTEMP_448),
        .in(_T_123)
    );
    MUX_UNSIGNED #(.width(25)) u_mux_3272 (
        .y(_T_124),
        .sel(_T_39),
        .a(_T_110),
        .b(_WTEMP_448)
    );
    wire [24:0] _T_126;
    wire [24:0] _WTEMP_449;
    PAD_UNSIGNED #(.width(1), .n(25)) u_pad_3273 (
        .y(_WTEMP_449),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(25)) u_mux_3274 (
        .y(_T_126),
        .sel(_T_37),
        .a(_T_124),
        .b(_WTEMP_449)
    );
    wire [24:0] _T_127;
    BITWISEOR #(.width(25)) bitwiseor_3275 (
        .y(_T_127),
        .a(_T_34),
        .b(_T_126)
    );
    wire [24:0] _T_128;
    wire [24:0] _WTEMP_450;
    PAD_UNSIGNED #(.width(1), .n(25)) u_pad_3276 (
        .y(_WTEMP_450),
        .in(doShiftSigDown1)
    );
    BITWISEOR #(.width(25)) bitwiseor_3277 (
        .y(_T_128),
        .a(_T_127),
        .b(_WTEMP_450)
    );
    wire [26:0] roundMask;
    CAT #(.width_a(25), .width_b(2)) cat_3278 (
        .y(roundMask),
        .a(_T_128),
        .b(2'h3)
    );
    wire [27:0] _T_130;
    CAT #(.width_a(1), .width_b(27)) cat_3279 (
        .y(_T_130),
        .a(isNegExp),
        .b(roundMask)
    );
    wire [26:0] shiftedRoundMask;
    SHR_UNSIGNED #(.width(28), .n(1)) u_shr_3280 (
        .y(shiftedRoundMask),
        .in(_T_130)
    );
    wire [26:0] _T_131;
    BITWISENOT #(.width(27)) bitwisenot_3281 (
        .y(_T_131),
        .in(shiftedRoundMask)
    );
    wire [26:0] roundPosMask;
    BITWISEAND #(.width(27)) bitwiseand_3282 (
        .y(roundPosMask),
        .a(_T_131),
        .b(roundMask)
    );
    wire [26:0] _T_132;
    BITWISEAND #(.width(27)) bitwiseand_3283 (
        .y(_T_132),
        .a(io_in_sig),
        .b(roundPosMask)
    );
    wire roundPosBit;
    wire [26:0] _WTEMP_451;
    PAD_UNSIGNED #(.width(1), .n(27)) u_pad_3284 (
        .y(_WTEMP_451),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(27)) u_neq_3285 (
        .y(roundPosBit),
        .a(_T_132),
        .b(_WTEMP_451)
    );
    wire [26:0] _T_134;
    BITWISEAND #(.width(27)) bitwiseand_3286 (
        .y(_T_134),
        .a(io_in_sig),
        .b(shiftedRoundMask)
    );
    wire anyRoundExtra;
    wire [26:0] _WTEMP_452;
    PAD_UNSIGNED #(.width(1), .n(27)) u_pad_3287 (
        .y(_WTEMP_452),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(27)) u_neq_3288 (
        .y(anyRoundExtra),
        .a(_T_134),
        .b(_WTEMP_452)
    );
    wire anyRound;
    BITWISEOR #(.width(1)) bitwiseor_3289 (
        .y(anyRound),
        .a(roundPosBit),
        .b(anyRoundExtra)
    );
    wire _T_136;
    BITWISEAND #(.width(1)) bitwiseand_3290 (
        .y(_T_136),
        .a(roundingMode_nearest_even),
        .b(roundPosBit)
    );
    wire _T_137;
    BITWISEAND #(.width(1)) bitwiseand_3291 (
        .y(_T_137),
        .a(roundMagUp),
        .b(anyRound)
    );
    wire _T_138;
    BITWISEOR #(.width(1)) bitwiseor_3292 (
        .y(_T_138),
        .a(_T_136),
        .b(_T_137)
    );
    wire [26:0] _T_139;
    BITWISEOR #(.width(27)) bitwiseor_3293 (
        .y(_T_139),
        .a(io_in_sig),
        .b(roundMask)
    );
    wire [24:0] _T_140;
    SHR_UNSIGNED #(.width(27), .n(2)) u_shr_3294 (
        .y(_T_140),
        .in(_T_139)
    );
    wire [25:0] _T_142;
    wire [24:0] _WTEMP_453;
    PAD_UNSIGNED #(.width(1), .n(25)) u_pad_3295 (
        .y(_WTEMP_453),
        .in(1'h1)
    );
    ADD_UNSIGNED #(.width(25)) u_add_3296 (
        .y(_T_142),
        .a(_T_140),
        .b(_WTEMP_453)
    );
    wire _T_143;
    BITWISEAND #(.width(1)) bitwiseand_3297 (
        .y(_T_143),
        .a(roundingMode_nearest_even),
        .b(roundPosBit)
    );
    wire _T_145;
    EQ_UNSIGNED #(.width(1)) u_eq_3298 (
        .y(_T_145),
        .a(anyRoundExtra),
        .b(1'h0)
    );
    wire _T_146;
    BITWISEAND #(.width(1)) bitwiseand_3299 (
        .y(_T_146),
        .a(_T_143),
        .b(_T_145)
    );
    wire [25:0] _T_147;
    SHR_UNSIGNED #(.width(27), .n(1)) u_shr_3300 (
        .y(_T_147),
        .in(roundMask)
    );
    wire [25:0] _T_149;
    MUX_UNSIGNED #(.width(26)) u_mux_3301 (
        .y(_T_149),
        .sel(_T_146),
        .a(_T_147),
        .b(26'h0)
    );
    wire [25:0] _T_150;
    BITWISENOT #(.width(26)) bitwisenot_3302 (
        .y(_T_150),
        .in(_T_149)
    );
    wire [25:0] _T_151;
    BITWISEAND #(.width(26)) bitwiseand_3303 (
        .y(_T_151),
        .a(_T_142),
        .b(_T_150)
    );
    wire [26:0] _T_152;
    BITWISENOT #(.width(27)) bitwisenot_3304 (
        .y(_T_152),
        .in(roundMask)
    );
    wire [26:0] _T_153;
    BITWISEAND #(.width(27)) bitwiseand_3305 (
        .y(_T_153),
        .a(io_in_sig),
        .b(_T_152)
    );
    wire [24:0] _T_154;
    SHR_UNSIGNED #(.width(27), .n(2)) u_shr_3306 (
        .y(_T_154),
        .in(_T_153)
    );
    wire [25:0] roundedSig;
    wire [25:0] _WTEMP_454;
    PAD_UNSIGNED #(.width(25), .n(26)) u_pad_3307 (
        .y(_WTEMP_454),
        .in(_T_154)
    );
    MUX_UNSIGNED #(.width(26)) u_mux_3308 (
        .y(roundedSig),
        .sel(_T_138),
        .a(_T_151),
        .b(_WTEMP_454)
    );
    wire [1:0] _T_155;
    SHR_UNSIGNED #(.width(26), .n(24)) u_shr_3309 (
        .y(_T_155),
        .in(roundedSig)
    );
    wire [2:0] _T_156;
    CVT_UNSIGNED #(.width(2)) u_cvt_3310 (
        .y(_T_156),
        .in(_T_155)
    );
    wire [10:0] sRoundedExp;
    wire [9:0] _WTEMP_455;
    PAD_SIGNED #(.width(3), .n(10)) s_pad_3311 (
        .y(_WTEMP_455),
        .in(_T_156)
    );
    ADD_SIGNED #(.width(10)) s_add_3312 (
        .y(sRoundedExp),
        .a(io_in_sExp),
        .b(_WTEMP_455)
    );
    wire [8:0] common_expOut;
    BITS #(.width(11), .high(8), .low(0)) bits_3313 (
        .y(common_expOut),
        .in(sRoundedExp)
    );
    wire [22:0] _T_157;
    BITS #(.width(26), .high(23), .low(1)) bits_3314 (
        .y(_T_157),
        .in(roundedSig)
    );
    wire [22:0] _T_158;
    BITS #(.width(26), .high(22), .low(0)) bits_3315 (
        .y(_T_158),
        .in(roundedSig)
    );
    wire [22:0] common_fractOut;
    MUX_UNSIGNED #(.width(23)) u_mux_3316 (
        .y(common_fractOut),
        .sel(doShiftSigDown1),
        .a(_T_157),
        .b(_T_158)
    );
    wire [3:0] _T_159;
    SHR_SIGNED #(.width(11), .n(7)) s_shr_3317 (
        .y(_T_159),
        .in(sRoundedExp)
    );
    wire common_overflow;
    wire [3:0] _WTEMP_456;
    PAD_SIGNED #(.width(3), .n(4)) s_pad_3318 (
        .y(_WTEMP_456),
        .in(3'sh3)
    );
    GEQ_SIGNED #(.width(4)) s_geq_3319 (
        .y(common_overflow),
        .a(_T_159),
        .b(_WTEMP_456)
    );
    wire common_totalUnderflow;
    wire [10:0] _WTEMP_457;
    PAD_SIGNED #(.width(8), .n(11)) s_pad_3320 (
        .y(_WTEMP_457),
        .in(8'sh6B)
    );
    LT_SIGNED #(.width(11)) s_lt_3321 (
        .y(common_totalUnderflow),
        .a(sRoundedExp),
        .b(_WTEMP_457)
    );
    wire [8:0] _T_164;
    MUX_SIGNED #(.width(9)) s_mux_3322 (
        .y(_T_164),
        .sel(doShiftSigDown1),
        .a(9'sh81),
        .b(9'sh82)
    );
    wire _T_165;
    wire [9:0] _WTEMP_458;
    PAD_SIGNED #(.width(9), .n(10)) s_pad_3323 (
        .y(_WTEMP_458),
        .in(_T_164)
    );
    LT_SIGNED #(.width(10)) s_lt_3324 (
        .y(_T_165),
        .a(io_in_sExp),
        .b(_WTEMP_458)
    );
    wire common_underflow;
    BITWISEAND #(.width(1)) bitwiseand_3325 (
        .y(common_underflow),
        .a(anyRound),
        .b(_T_165)
    );
    wire isNaNOut;
    BITWISEOR #(.width(1)) bitwiseor_3326 (
        .y(isNaNOut),
        .a(io_invalidExc),
        .b(io_in_isNaN)
    );
    wire notNaN_isSpecialInfOut;
    BITWISEOR #(.width(1)) bitwiseor_3327 (
        .y(notNaN_isSpecialInfOut),
        .a(io_infiniteExc),
        .b(io_in_isInf)
    );
    wire _T_167;
    EQ_UNSIGNED #(.width(1)) u_eq_3328 (
        .y(_T_167),
        .a(isNaNOut),
        .b(1'h0)
    );
    wire _T_169;
    EQ_UNSIGNED #(.width(1)) u_eq_3329 (
        .y(_T_169),
        .a(notNaN_isSpecialInfOut),
        .b(1'h0)
    );
    wire _T_170;
    BITWISEAND #(.width(1)) bitwiseand_3330 (
        .y(_T_170),
        .a(_T_167),
        .b(_T_169)
    );
    wire _T_172;
    EQ_UNSIGNED #(.width(1)) u_eq_3331 (
        .y(_T_172),
        .a(io_in_isZero),
        .b(1'h0)
    );
    wire commonCase;
    BITWISEAND #(.width(1)) bitwiseand_3332 (
        .y(commonCase),
        .a(_T_170),
        .b(_T_172)
    );
    wire overflow;
    BITWISEAND #(.width(1)) bitwiseand_3333 (
        .y(overflow),
        .a(commonCase),
        .b(common_overflow)
    );
    wire underflow;
    BITWISEAND #(.width(1)) bitwiseand_3334 (
        .y(underflow),
        .a(commonCase),
        .b(common_underflow)
    );
    wire _T_173;
    BITWISEAND #(.width(1)) bitwiseand_3335 (
        .y(_T_173),
        .a(commonCase),
        .b(anyRound)
    );
    wire inexact;
    BITWISEOR #(.width(1)) bitwiseor_3336 (
        .y(inexact),
        .a(overflow),
        .b(_T_173)
    );
    wire overflow_roundMagUp;
    BITWISEOR #(.width(1)) bitwiseor_3337 (
        .y(overflow_roundMagUp),
        .a(roundingMode_nearest_even),
        .b(roundMagUp)
    );
    wire _T_174;
    BITWISEAND #(.width(1)) bitwiseand_3338 (
        .y(_T_174),
        .a(commonCase),
        .b(common_totalUnderflow)
    );
    wire pegMinNonzeroMagOut;
    BITWISEAND #(.width(1)) bitwiseand_3339 (
        .y(pegMinNonzeroMagOut),
        .a(_T_174),
        .b(roundMagUp)
    );
    wire _T_175;
    BITWISEAND #(.width(1)) bitwiseand_3340 (
        .y(_T_175),
        .a(commonCase),
        .b(overflow)
    );
    wire _T_177;
    EQ_UNSIGNED #(.width(1)) u_eq_3341 (
        .y(_T_177),
        .a(overflow_roundMagUp),
        .b(1'h0)
    );
    wire pegMaxFiniteMagOut;
    BITWISEAND #(.width(1)) bitwiseand_3342 (
        .y(pegMaxFiniteMagOut),
        .a(_T_175),
        .b(_T_177)
    );
    wire _T_178;
    BITWISEAND #(.width(1)) bitwiseand_3343 (
        .y(_T_178),
        .a(overflow),
        .b(overflow_roundMagUp)
    );
    wire notNaN_isInfOut;
    BITWISEOR #(.width(1)) bitwiseor_3344 (
        .y(notNaN_isInfOut),
        .a(notNaN_isSpecialInfOut),
        .b(_T_178)
    );
    wire signOut;
    MUX_UNSIGNED #(.width(1)) u_mux_3345 (
        .y(signOut),
        .sel(isNaNOut),
        .a(1'h0),
        .b(io_in_sign)
    );
    wire _T_180;
    BITWISEOR #(.width(1)) bitwiseor_3346 (
        .y(_T_180),
        .a(io_in_isZero),
        .b(common_totalUnderflow)
    );
    wire [8:0] _T_183;
    wire [8:0] _WTEMP_459;
    PAD_UNSIGNED #(.width(1), .n(9)) u_pad_3347 (
        .y(_WTEMP_459),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(9)) u_mux_3348 (
        .y(_T_183),
        .sel(_T_180),
        .a(9'h1C0),
        .b(_WTEMP_459)
    );
    wire [8:0] _T_184;
    BITWISENOT #(.width(9)) bitwisenot_3349 (
        .y(_T_184),
        .in(_T_183)
    );
    wire [8:0] _T_185;
    BITWISEAND #(.width(9)) bitwiseand_3350 (
        .y(_T_185),
        .a(common_expOut),
        .b(_T_184)
    );
    wire [8:0] _T_187;
    assign _T_187 = 9'h194;
    wire [8:0] _T_189;
    wire [8:0] _WTEMP_460;
    PAD_UNSIGNED #(.width(1), .n(9)) u_pad_3351 (
        .y(_WTEMP_460),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(9)) u_mux_3352 (
        .y(_T_189),
        .sel(pegMinNonzeroMagOut),
        .a(_T_187),
        .b(_WTEMP_460)
    );
    wire [8:0] _T_190;
    BITWISENOT #(.width(9)) bitwisenot_3353 (
        .y(_T_190),
        .in(_T_189)
    );
    wire [8:0] _T_191;
    BITWISEAND #(.width(9)) bitwiseand_3354 (
        .y(_T_191),
        .a(_T_185),
        .b(_T_190)
    );
    wire [8:0] _T_194;
    wire [8:0] _WTEMP_461;
    PAD_UNSIGNED #(.width(1), .n(9)) u_pad_3355 (
        .y(_WTEMP_461),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(9)) u_mux_3356 (
        .y(_T_194),
        .sel(pegMaxFiniteMagOut),
        .a(9'h80),
        .b(_WTEMP_461)
    );
    wire [8:0] _T_195;
    BITWISENOT #(.width(9)) bitwisenot_3357 (
        .y(_T_195),
        .in(_T_194)
    );
    wire [8:0] _T_196;
    BITWISEAND #(.width(9)) bitwiseand_3358 (
        .y(_T_196),
        .a(_T_191),
        .b(_T_195)
    );
    wire [8:0] _T_199;
    wire [8:0] _WTEMP_462;
    PAD_UNSIGNED #(.width(1), .n(9)) u_pad_3359 (
        .y(_WTEMP_462),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(9)) u_mux_3360 (
        .y(_T_199),
        .sel(notNaN_isInfOut),
        .a(9'h40),
        .b(_WTEMP_462)
    );
    wire [8:0] _T_200;
    BITWISENOT #(.width(9)) bitwisenot_3361 (
        .y(_T_200),
        .in(_T_199)
    );
    wire [8:0] _T_201;
    BITWISEAND #(.width(9)) bitwiseand_3362 (
        .y(_T_201),
        .a(_T_196),
        .b(_T_200)
    );
    wire [8:0] _T_204;
    wire [8:0] _WTEMP_463;
    PAD_UNSIGNED #(.width(1), .n(9)) u_pad_3363 (
        .y(_WTEMP_463),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(9)) u_mux_3364 (
        .y(_T_204),
        .sel(pegMinNonzeroMagOut),
        .a(9'h6B),
        .b(_WTEMP_463)
    );
    wire [8:0] _T_205;
    BITWISEOR #(.width(9)) bitwiseor_3365 (
        .y(_T_205),
        .a(_T_201),
        .b(_T_204)
    );
    wire [8:0] _T_208;
    wire [8:0] _WTEMP_464;
    PAD_UNSIGNED #(.width(1), .n(9)) u_pad_3366 (
        .y(_WTEMP_464),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(9)) u_mux_3367 (
        .y(_T_208),
        .sel(pegMaxFiniteMagOut),
        .a(9'h17F),
        .b(_WTEMP_464)
    );
    wire [8:0] _T_209;
    BITWISEOR #(.width(9)) bitwiseor_3368 (
        .y(_T_209),
        .a(_T_205),
        .b(_T_208)
    );
    wire [8:0] _T_212;
    wire [8:0] _WTEMP_465;
    PAD_UNSIGNED #(.width(1), .n(9)) u_pad_3369 (
        .y(_WTEMP_465),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(9)) u_mux_3370 (
        .y(_T_212),
        .sel(notNaN_isInfOut),
        .a(9'h180),
        .b(_WTEMP_465)
    );
    wire [8:0] _T_213;
    BITWISEOR #(.width(9)) bitwiseor_3371 (
        .y(_T_213),
        .a(_T_209),
        .b(_T_212)
    );
    wire [8:0] _T_216;
    wire [8:0] _WTEMP_466;
    PAD_UNSIGNED #(.width(1), .n(9)) u_pad_3372 (
        .y(_WTEMP_466),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(9)) u_mux_3373 (
        .y(_T_216),
        .sel(isNaNOut),
        .a(9'h1C0),
        .b(_WTEMP_466)
    );
    wire [8:0] expOut;
    BITWISEOR #(.width(9)) bitwiseor_3374 (
        .y(expOut),
        .a(_T_213),
        .b(_T_216)
    );
    wire _T_217;
    BITWISEOR #(.width(1)) bitwiseor_3375 (
        .y(_T_217),
        .a(common_totalUnderflow),
        .b(isNaNOut)
    );
    wire [22:0] _T_219;
    assign _T_219 = 23'h400000;
    wire [22:0] _T_221;
    wire [22:0] _WTEMP_467;
    PAD_UNSIGNED #(.width(1), .n(23)) u_pad_3376 (
        .y(_WTEMP_467),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(23)) u_mux_3377 (
        .y(_T_221),
        .sel(isNaNOut),
        .a(_T_219),
        .b(_WTEMP_467)
    );
    wire [22:0] _T_222;
    MUX_UNSIGNED #(.width(23)) u_mux_3378 (
        .y(_T_222),
        .sel(_T_217),
        .a(_T_221),
        .b(common_fractOut)
    );
    wire _T_223;
    BITS #(.width(1), .high(0), .low(0)) bits_3379 (
        .y(_T_223),
        .in(pegMaxFiniteMagOut)
    );
    wire [22:0] _T_226;
    MUX_UNSIGNED #(.width(23)) u_mux_3380 (
        .y(_T_226),
        .sel(_T_223),
        .a(23'h7FFFFF),
        .b(23'h0)
    );
    wire [22:0] fractOut;
    BITWISEOR #(.width(23)) bitwiseor_3381 (
        .y(fractOut),
        .a(_T_222),
        .b(_T_226)
    );
    wire [9:0] _T_227;
    CAT #(.width_a(1), .width_b(9)) cat_3382 (
        .y(_T_227),
        .a(signOut),
        .b(expOut)
    );
    wire [32:0] _T_228;
    CAT #(.width_a(10), .width_b(23)) cat_3383 (
        .y(_T_228),
        .a(_T_227),
        .b(fractOut)
    );
    wire [1:0] _T_229;
    CAT #(.width_a(1), .width_b(1)) cat_3384 (
        .y(_T_229),
        .a(underflow),
        .b(inexact)
    );
    wire [1:0] _T_230;
    CAT #(.width_a(1), .width_b(1)) cat_3385 (
        .y(_T_230),
        .a(io_invalidExc),
        .b(io_infiniteExc)
    );
    wire [2:0] _T_231;
    CAT #(.width_a(2), .width_b(1)) cat_3386 (
        .y(_T_231),
        .a(_T_230),
        .b(overflow)
    );
    wire [4:0] _T_232;
    CAT #(.width_a(3), .width_b(2)) cat_3387 (
        .y(_T_232),
        .a(_T_231),
        .b(_T_229)
    );
    assign io_exceptionFlags = _T_232;
    assign io_out = _T_228;
endmodule //RoundRawFNToRecFN
module SHR_SIGNED(y, in);
    parameter width = 4;
    parameter n = 2;
    output [(n < width ? (width-n-1) : 0):0] y;
    input [width-1:0] in;
    assign y = n < width ? in[width-1:n] : in[width-1:width-1];
endmodule // SHR_SIGNED
module GEQ_SIGNED(y, a, b);
    parameter width = 4;
    output y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = $signed(a) >= $signed(b);
endmodule // GEQ_SIGNED
module RecFNToRecFN_1(
    input clock,
    input reset,
    input [32:0] io_in,
    input [1:0] io_roundingMode,
    output [64:0] io_out,
    output [4:0] io_exceptionFlags
);
    wire [8:0] _T_10;
    BITS #(.width(33), .high(31), .low(23)) bits_3388 (
        .y(_T_10),
        .in(io_in)
    );
    wire [2:0] _T_11;
    BITS #(.width(9), .high(8), .low(6)) bits_3389 (
        .y(_T_11),
        .in(_T_10)
    );
    wire _T_13;
    wire [2:0] _WTEMP_468;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_3390 (
        .y(_WTEMP_468),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(3)) u_eq_3391 (
        .y(_T_13),
        .a(_T_11),
        .b(_WTEMP_468)
    );
    wire [1:0] _T_14;
    BITS #(.width(9), .high(8), .low(7)) bits_3392 (
        .y(_T_14),
        .in(_T_10)
    );
    wire _T_16;
    EQ_UNSIGNED #(.width(2)) u_eq_3393 (
        .y(_T_16),
        .a(_T_14),
        .b(2'h3)
    );
    wire _T_24_sign;
    wire _T_24_isNaN;
    wire _T_24_isInf;
    wire _T_24_isZero;
    wire [9:0] _T_24_sExp;
    wire [26:0] _T_24_sig;
    wire _T_31;
    BITS #(.width(33), .high(32), .low(32)) bits_3394 (
        .y(_T_31),
        .in(io_in)
    );
    wire _T_32;
    BITS #(.width(9), .high(6), .low(6)) bits_3395 (
        .y(_T_32),
        .in(_T_10)
    );
    wire _T_33;
    BITWISEAND #(.width(1)) bitwiseand_3396 (
        .y(_T_33),
        .a(_T_16),
        .b(_T_32)
    );
    wire _T_34;
    BITS #(.width(9), .high(6), .low(6)) bits_3397 (
        .y(_T_34),
        .in(_T_10)
    );
    wire _T_36;
    EQ_UNSIGNED #(.width(1)) u_eq_3398 (
        .y(_T_36),
        .a(_T_34),
        .b(1'h0)
    );
    wire _T_37;
    BITWISEAND #(.width(1)) bitwiseand_3399 (
        .y(_T_37),
        .a(_T_16),
        .b(_T_36)
    );
    wire [9:0] _T_38;
    CVT_UNSIGNED #(.width(9)) u_cvt_3400 (
        .y(_T_38),
        .in(_T_10)
    );
    wire _T_41;
    EQ_UNSIGNED #(.width(1)) u_eq_3401 (
        .y(_T_41),
        .a(_T_13),
        .b(1'h0)
    );
    wire [22:0] _T_42;
    BITS #(.width(33), .high(22), .low(0)) bits_3402 (
        .y(_T_42),
        .in(io_in)
    );
    wire [24:0] _T_44;
    CAT #(.width_a(23), .width_b(2)) cat_3403 (
        .y(_T_44),
        .a(_T_42),
        .b(2'h0)
    );
    wire [1:0] _T_45;
    CAT #(.width_a(1), .width_b(1)) cat_3404 (
        .y(_T_45),
        .a(1'h0),
        .b(_T_41)
    );
    wire [26:0] _T_46;
    CAT #(.width_a(2), .width_b(25)) cat_3405 (
        .y(_T_46),
        .a(_T_45),
        .b(_T_44)
    );
    wire [12:0] _T_48;
    wire [11:0] _WTEMP_469;
    PAD_SIGNED #(.width(10), .n(12)) s_pad_3406 (
        .y(_WTEMP_469),
        .in(_T_24_sExp)
    );
    ADD_SIGNED #(.width(12)) s_add_3407 (
        .y(_T_48),
        .a(_WTEMP_469),
        .b(12'sh700)
    );
    wire outRawFloat_sign;
    wire outRawFloat_isNaN;
    wire outRawFloat_isInf;
    wire outRawFloat_isZero;
    wire [12:0] outRawFloat_sExp;
    wire [55:0] outRawFloat_sig;
    wire [55:0] _T_62;
    SHL_UNSIGNED #(.width(27), .n(29)) u_shl_3408 (
        .y(_T_62),
        .in(_T_24_sig)
    );
    wire _T_63;
    BITS #(.width(56), .high(53), .low(53)) bits_3409 (
        .y(_T_63),
        .in(outRawFloat_sig)
    );
    wire _T_65;
    EQ_UNSIGNED #(.width(1)) u_eq_3410 (
        .y(_T_65),
        .a(_T_63),
        .b(1'h0)
    );
    wire invalidExc;
    BITWISEAND #(.width(1)) bitwiseand_3411 (
        .y(invalidExc),
        .a(outRawFloat_isNaN),
        .b(_T_65)
    );
    wire _T_67;
    EQ_UNSIGNED #(.width(1)) u_eq_3412 (
        .y(_T_67),
        .a(outRawFloat_isNaN),
        .b(1'h0)
    );
    wire _T_68;
    BITWISEAND #(.width(1)) bitwiseand_3413 (
        .y(_T_68),
        .a(outRawFloat_sign),
        .b(_T_67)
    );
    wire [11:0] _T_69;
    BITS #(.width(13), .high(11), .low(0)) bits_3414 (
        .y(_T_69),
        .in(outRawFloat_sExp)
    );
    wire [11:0] _T_72;
    wire [11:0] _WTEMP_470;
    PAD_UNSIGNED #(.width(1), .n(12)) u_pad_3415 (
        .y(_WTEMP_470),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(12)) u_mux_3416 (
        .y(_T_72),
        .sel(outRawFloat_isZero),
        .a(12'hC00),
        .b(_WTEMP_470)
    );
    wire [11:0] _T_73;
    BITWISENOT #(.width(12)) bitwisenot_3417 (
        .y(_T_73),
        .in(_T_72)
    );
    wire [11:0] _T_74;
    BITWISEAND #(.width(12)) bitwiseand_3418 (
        .y(_T_74),
        .a(_T_69),
        .b(_T_73)
    );
    wire _T_75;
    BITWISEOR #(.width(1)) bitwiseor_3419 (
        .y(_T_75),
        .a(outRawFloat_isZero),
        .b(outRawFloat_isInf)
    );
    wire [11:0] _T_78;
    wire [11:0] _WTEMP_471;
    PAD_UNSIGNED #(.width(1), .n(12)) u_pad_3420 (
        .y(_WTEMP_471),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(12)) u_mux_3421 (
        .y(_T_78),
        .sel(_T_75),
        .a(12'h200),
        .b(_WTEMP_471)
    );
    wire [11:0] _T_79;
    BITWISENOT #(.width(12)) bitwisenot_3422 (
        .y(_T_79),
        .in(_T_78)
    );
    wire [11:0] _T_80;
    BITWISEAND #(.width(12)) bitwiseand_3423 (
        .y(_T_80),
        .a(_T_74),
        .b(_T_79)
    );
    wire [11:0] _T_83;
    wire [11:0] _WTEMP_472;
    PAD_UNSIGNED #(.width(1), .n(12)) u_pad_3424 (
        .y(_WTEMP_472),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(12)) u_mux_3425 (
        .y(_T_83),
        .sel(outRawFloat_isInf),
        .a(12'hC00),
        .b(_WTEMP_472)
    );
    wire [11:0] _T_84;
    BITWISEOR #(.width(12)) bitwiseor_3426 (
        .y(_T_84),
        .a(_T_80),
        .b(_T_83)
    );
    wire [11:0] _T_87;
    wire [11:0] _WTEMP_473;
    PAD_UNSIGNED #(.width(1), .n(12)) u_pad_3427 (
        .y(_WTEMP_473),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(12)) u_mux_3428 (
        .y(_T_87),
        .sel(outRawFloat_isNaN),
        .a(12'hE00),
        .b(_WTEMP_473)
    );
    wire [11:0] _T_88;
    BITWISEOR #(.width(12)) bitwiseor_3429 (
        .y(_T_88),
        .a(_T_84),
        .b(_T_87)
    );
    wire [51:0] _T_90;
    assign _T_90 = 52'h8000000000000;
    wire [51:0] _T_91;
    BITS #(.width(56), .high(53), .low(2)) bits_3430 (
        .y(_T_91),
        .in(outRawFloat_sig)
    );
    wire [51:0] _T_92;
    MUX_UNSIGNED #(.width(52)) u_mux_3431 (
        .y(_T_92),
        .sel(outRawFloat_isNaN),
        .a(_T_90),
        .b(_T_91)
    );
    wire [12:0] _T_93;
    CAT #(.width_a(1), .width_b(12)) cat_3432 (
        .y(_T_93),
        .a(_T_68),
        .b(_T_88)
    );
    wire [64:0] _T_94;
    CAT #(.width_a(13), .width_b(52)) cat_3433 (
        .y(_T_94),
        .a(_T_93),
        .b(_T_92)
    );
    wire [4:0] _T_96;
    CAT #(.width_a(1), .width_b(4)) cat_3434 (
        .y(_T_96),
        .a(invalidExc),
        .b(4'h0)
    );
    assign _T_24_isInf = _T_37;
    assign _T_24_isNaN = _T_33;
    assign _T_24_isZero = _T_13;
    assign _T_24_sExp = _T_38;
    assign _T_24_sig = _T_46;
    assign _T_24_sign = _T_31;
    assign io_exceptionFlags = _T_96;
    assign io_out = _T_94;
    assign outRawFloat_isInf = _T_24_isInf;
    assign outRawFloat_isNaN = _T_24_isNaN;
    assign outRawFloat_isZero = _T_24_isZero;
    assign outRawFloat_sExp = _T_48;
    assign outRawFloat_sig = _T_62;
    assign outRawFloat_sign = _T_24_sign;
endmodule //RecFNToRecFN_1
module FPUFMAPipe_1(
    input clock,
    input reset,
    input io_in_valid,
    input [4:0] io_in_bits_cmd,
    input io_in_bits_ldst,
    input io_in_bits_wen,
    input io_in_bits_ren1,
    input io_in_bits_ren2,
    input io_in_bits_ren3,
    input io_in_bits_swap12,
    input io_in_bits_swap23,
    input io_in_bits_single,
    input io_in_bits_fromint,
    input io_in_bits_toint,
    input io_in_bits_fastpipe,
    input io_in_bits_fma,
    input io_in_bits_div,
    input io_in_bits_sqrt,
    input io_in_bits_wflags,
    input [2:0] io_in_bits_rm,
    input [1:0] io_in_bits_typ,
    input [64:0] io_in_bits_in1,
    input [64:0] io_in_bits_in2,
    input [64:0] io_in_bits_in3,
    output io_out_valid,
    output [64:0] io_out_bits_data,
    output [4:0] io_out_bits_exc
);
    wire [63:0] one;
    assign one = 64'h8000000000000000;
    wire _T_131;
    BITS #(.width(65), .high(64), .low(64)) bits_3479 (
        .y(_T_131),
        .in(io_in_bits_in1)
    );
    wire _T_132;
    BITS #(.width(65), .high(64), .low(64)) bits_3480 (
        .y(_T_132),
        .in(io_in_bits_in2)
    );
    wire _T_133;
    BITWISEXOR #(.width(1)) bitwisexor_3481 (
        .y(_T_133),
        .a(_T_131),
        .b(_T_132)
    );
    wire [64:0] zero;
    SHL_UNSIGNED #(.width(1), .n(64)) u_shl_3482 (
        .y(zero),
        .in(_T_133)
    );
    wire _valid__q;
    wire _valid__d;
    DFF_POSCLK #(.width(1)) valid (
        .q(_valid__q),
        .d(_valid__d),
        .clk(clock)
    );
    wire [4:0] _in_cmd__q;
    wire [4:0] _in_cmd__d;
    DFF_POSCLK #(.width(5)) in_cmd (
        .q(_in_cmd__q),
        .d(_in_cmd__d),
        .clk(clock)
    );
    wire _in_ldst__q;
    wire _in_ldst__d;
    DFF_POSCLK #(.width(1)) in_ldst (
        .q(_in_ldst__q),
        .d(_in_ldst__d),
        .clk(clock)
    );
    wire _in_wen__q;
    wire _in_wen__d;
    DFF_POSCLK #(.width(1)) in_wen (
        .q(_in_wen__q),
        .d(_in_wen__d),
        .clk(clock)
    );
    wire _in_ren1__q;
    wire _in_ren1__d;
    DFF_POSCLK #(.width(1)) in_ren1 (
        .q(_in_ren1__q),
        .d(_in_ren1__d),
        .clk(clock)
    );
    wire _in_ren2__q;
    wire _in_ren2__d;
    DFF_POSCLK #(.width(1)) in_ren2 (
        .q(_in_ren2__q),
        .d(_in_ren2__d),
        .clk(clock)
    );
    wire _in_ren3__q;
    wire _in_ren3__d;
    DFF_POSCLK #(.width(1)) in_ren3 (
        .q(_in_ren3__q),
        .d(_in_ren3__d),
        .clk(clock)
    );
    wire _in_swap12__q;
    wire _in_swap12__d;
    DFF_POSCLK #(.width(1)) in_swap12 (
        .q(_in_swap12__q),
        .d(_in_swap12__d),
        .clk(clock)
    );
    wire _in_swap23__q;
    wire _in_swap23__d;
    DFF_POSCLK #(.width(1)) in_swap23 (
        .q(_in_swap23__q),
        .d(_in_swap23__d),
        .clk(clock)
    );
    wire _in_single__q;
    wire _in_single__d;
    DFF_POSCLK #(.width(1)) in_single (
        .q(_in_single__q),
        .d(_in_single__d),
        .clk(clock)
    );
    wire _in_fromint__q;
    wire _in_fromint__d;
    DFF_POSCLK #(.width(1)) in_fromint (
        .q(_in_fromint__q),
        .d(_in_fromint__d),
        .clk(clock)
    );
    wire _in_toint__q;
    wire _in_toint__d;
    DFF_POSCLK #(.width(1)) in_toint (
        .q(_in_toint__q),
        .d(_in_toint__d),
        .clk(clock)
    );
    wire _in_fastpipe__q;
    wire _in_fastpipe__d;
    DFF_POSCLK #(.width(1)) in_fastpipe (
        .q(_in_fastpipe__q),
        .d(_in_fastpipe__d),
        .clk(clock)
    );
    wire _in_fma__q;
    wire _in_fma__d;
    DFF_POSCLK #(.width(1)) in_fma (
        .q(_in_fma__q),
        .d(_in_fma__d),
        .clk(clock)
    );
    wire _in_div__q;
    wire _in_div__d;
    DFF_POSCLK #(.width(1)) in_div (
        .q(_in_div__q),
        .d(_in_div__d),
        .clk(clock)
    );
    wire _in_sqrt__q;
    wire _in_sqrt__d;
    DFF_POSCLK #(.width(1)) in_sqrt (
        .q(_in_sqrt__q),
        .d(_in_sqrt__d),
        .clk(clock)
    );
    wire _in_wflags__q;
    wire _in_wflags__d;
    DFF_POSCLK #(.width(1)) in_wflags (
        .q(_in_wflags__q),
        .d(_in_wflags__d),
        .clk(clock)
    );
    wire [2:0] _in_rm__q;
    wire [2:0] _in_rm__d;
    DFF_POSCLK #(.width(3)) in_rm (
        .q(_in_rm__q),
        .d(_in_rm__d),
        .clk(clock)
    );
    wire [1:0] _in_typ__q;
    wire [1:0] _in_typ__d;
    DFF_POSCLK #(.width(2)) in_typ (
        .q(_in_typ__q),
        .d(_in_typ__d),
        .clk(clock)
    );
    wire [64:0] _in_in1__q;
    wire [64:0] _in_in1__d;
    DFF_POSCLK #(.width(65)) in_in1 (
        .q(_in_in1__q),
        .d(_in_in1__d),
        .clk(clock)
    );
    wire [64:0] _in_in2__q;
    wire [64:0] _in_in2__d;
    DFF_POSCLK #(.width(65)) in_in2 (
        .q(_in_in2__q),
        .d(_in_in2__d),
        .clk(clock)
    );
    wire [64:0] _in_in3__q;
    wire [64:0] _in_in3__d;
    DFF_POSCLK #(.width(65)) in_in3 (
        .q(_in_in3__q),
        .d(_in_in3__d),
        .clk(clock)
    );
    wire _T_177;
    BITS #(.width(5), .high(1), .low(1)) bits_3483 (
        .y(_T_177),
        .in(io_in_bits_cmd)
    );
    wire _T_178;
    BITWISEOR #(.width(1)) bitwiseor_3484 (
        .y(_T_178),
        .a(io_in_bits_ren3),
        .b(io_in_bits_swap23)
    );
    wire _T_179;
    BITWISEAND #(.width(1)) bitwiseand_3485 (
        .y(_T_179),
        .a(_T_177),
        .b(_T_178)
    );
    wire _T_180;
    BITS #(.width(5), .high(0), .low(0)) bits_3486 (
        .y(_T_180),
        .in(io_in_bits_cmd)
    );
    wire [1:0] _T_181;
    CAT #(.width_a(1), .width_b(1)) cat_3487 (
        .y(_T_181),
        .a(_T_179),
        .b(_T_180)
    );
    wire _T_182;
    BITWISEOR #(.width(1)) bitwiseor_3488 (
        .y(_T_182),
        .a(io_in_bits_ren3),
        .b(io_in_bits_swap23)
    );
    wire _T_184;
    EQ_UNSIGNED #(.width(1)) u_eq_3489 (
        .y(_T_184),
        .a(_T_182),
        .b(1'h0)
    );
    wire [64:0] _node_38;
    wire [64:0] _WTEMP_478;
    PAD_UNSIGNED #(.width(64), .n(65)) u_pad_3490 (
        .y(_WTEMP_478),
        .in(64'h8000000000000000)
    );
    MUX_UNSIGNED #(.width(65)) u_mux_3491 (
        .y(_node_38),
        .sel(io_in_bits_swap23),
        .a(_WTEMP_478),
        .b(io_in_bits_in2)
    );
    wire [64:0] _node_39;
    MUX_UNSIGNED #(.width(65)) u_mux_3492 (
        .y(_node_39),
        .sel(_T_184),
        .a(zero),
        .b(io_in_bits_in3)
    );
    wire _fma__clock;
    wire _fma__reset;
    wire [1:0] _fma__io_op;
    wire [64:0] _fma__io_a;
    wire [64:0] _fma__io_b;
    wire [64:0] _fma__io_c;
    wire [1:0] _fma__io_roundingMode;
    wire [64:0] _fma__io_out;
    wire [4:0] _fma__io_exceptionFlags;
    MulAddRecFN_1 fma (
        .clock(_fma__clock),
        .reset(_fma__reset),
        .io_op(_fma__io_op),
        .io_a(_fma__io_a),
        .io_b(_fma__io_b),
        .io_c(_fma__io_c),
        .io_roundingMode(_fma__io_roundingMode),
        .io_out(_fma__io_out),
        .io_exceptionFlags(_fma__io_exceptionFlags)
    );
    wire [64:0] res_data;
    wire [4:0] res_exc;
    wire __T_192__q;
    wire __T_192__d;
    DFF_POSCLK #(.width(1)) _T_192 (
        .q(__T_192__q),
        .d(__T_192__d),
        .clk(clock)
    );
    wire _WTEMP_642;
    MUX_UNSIGNED #(.width(1)) u_mux_4661 (
        .y(__T_192__d),
        .sel(reset),
        .a(1'h0),
        .b(_WTEMP_642)
    );
    wire [64:0] __T_196_data__q;
    wire [64:0] __T_196_data__d;
    DFF_POSCLK #(.width(65)) _T_196_data (
        .q(__T_196_data__q),
        .d(__T_196_data__d),
        .clk(clock)
    );
    wire [4:0] __T_196_exc__q;
    wire [4:0] __T_196_exc__d;
    DFF_POSCLK #(.width(5)) _T_196_exc (
        .q(__T_196_exc__q),
        .d(__T_196_exc__d),
        .clk(clock)
    );
    wire __T_201__q;
    wire __T_201__d;
    DFF_POSCLK #(.width(1)) _T_201 (
        .q(__T_201__q),
        .d(__T_201__d),
        .clk(clock)
    );
    wire _WTEMP_643;
    MUX_UNSIGNED #(.width(1)) u_mux_4662 (
        .y(__T_201__d),
        .sel(reset),
        .a(1'h0),
        .b(_WTEMP_643)
    );
    wire [64:0] __T_205_data__q;
    wire [64:0] __T_205_data__d;
    DFF_POSCLK #(.width(65)) _T_205_data (
        .q(__T_205_data__q),
        .d(__T_205_data__d),
        .clk(clock)
    );
    wire [4:0] __T_205_exc__q;
    wire [4:0] __T_205_exc__d;
    DFF_POSCLK #(.width(5)) _T_205_exc (
        .q(__T_205_exc__q),
        .d(__T_205_exc__d),
        .clk(clock)
    );
    wire __T_210__q;
    wire __T_210__d;
    DFF_POSCLK #(.width(1)) _T_210 (
        .q(__T_210__q),
        .d(__T_210__d),
        .clk(clock)
    );
    wire _WTEMP_644;
    MUX_UNSIGNED #(.width(1)) u_mux_4663 (
        .y(__T_210__d),
        .sel(reset),
        .a(1'h0),
        .b(_WTEMP_644)
    );
    wire [64:0] __T_214_data__q;
    wire [64:0] __T_214_data__d;
    DFF_POSCLK #(.width(65)) _T_214_data (
        .q(__T_214_data__q),
        .d(__T_214_data__d),
        .clk(clock)
    );
    wire [4:0] __T_214_exc__q;
    wire [4:0] __T_214_exc__d;
    DFF_POSCLK #(.width(5)) _T_214_exc (
        .q(__T_214_exc__q),
        .d(__T_214_exc__d),
        .clk(clock)
    );
    wire _T_226_valid;
    wire [64:0] _T_226_bits_data;
    wire [4:0] _T_226_bits_exc;
    assign _WTEMP_642 = _valid__q;
    MUX_UNSIGNED #(.width(65)) u_mux_4664 (
        .y(__T_196_data__d),
        .sel(_valid__q),
        .a(res_data),
        .b(__T_196_data__q)
    );
    MUX_UNSIGNED #(.width(5)) u_mux_4665 (
        .y(__T_196_exc__d),
        .sel(_valid__q),
        .a(res_exc),
        .b(__T_196_exc__q)
    );
    assign _WTEMP_643 = __T_192__q;
    MUX_UNSIGNED #(.width(65)) u_mux_4666 (
        .y(__T_205_data__d),
        .sel(__T_192__q),
        .a(__T_196_data__q),
        .b(__T_205_data__q)
    );
    MUX_UNSIGNED #(.width(5)) u_mux_4667 (
        .y(__T_205_exc__d),
        .sel(__T_192__q),
        .a(__T_196_exc__q),
        .b(__T_205_exc__q)
    );
    assign _WTEMP_644 = __T_201__q;
    MUX_UNSIGNED #(.width(65)) u_mux_4668 (
        .y(__T_214_data__d),
        .sel(__T_201__q),
        .a(__T_205_data__q),
        .b(__T_214_data__q)
    );
    MUX_UNSIGNED #(.width(5)) u_mux_4669 (
        .y(__T_214_exc__d),
        .sel(__T_201__q),
        .a(__T_205_exc__q),
        .b(__T_214_exc__q)
    );
    assign _T_226_bits_data = __T_214_data__q;
    assign _T_226_bits_exc = __T_214_exc__q;
    assign _T_226_valid = __T_210__q;
    assign _fma__clock = clock;
    assign _fma__io_a = _in_in1__q;
    assign _fma__io_b = _in_in2__q;
    assign _fma__io_c = _in_in3__q;
    BITS #(.width(5), .high(1), .low(0)) bits_4670 (
        .y(_fma__io_op),
        .in(_in_cmd__q)
    );
    BITS #(.width(3), .high(1), .low(0)) bits_4671 (
        .y(_fma__io_roundingMode),
        .in(_in_rm__q)
    );
    assign _fma__reset = reset;
    wire [4:0] _WTEMP_645;
    PAD_UNSIGNED #(.width(2), .n(5)) u_pad_4672 (
        .y(_WTEMP_645),
        .in(_T_181)
    );
    MUX_UNSIGNED #(.width(5)) u_mux_4673 (
        .y(_in_cmd__d),
        .sel(io_in_valid),
        .a(_WTEMP_645),
        .b(_in_cmd__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_4674 (
        .y(_in_div__d),
        .sel(io_in_valid),
        .a(io_in_bits_div),
        .b(_in_div__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_4675 (
        .y(_in_fastpipe__d),
        .sel(io_in_valid),
        .a(io_in_bits_fastpipe),
        .b(_in_fastpipe__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_4676 (
        .y(_in_fma__d),
        .sel(io_in_valid),
        .a(io_in_bits_fma),
        .b(_in_fma__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_4677 (
        .y(_in_fromint__d),
        .sel(io_in_valid),
        .a(io_in_bits_fromint),
        .b(_in_fromint__q)
    );
    MUX_UNSIGNED #(.width(65)) u_mux_4678 (
        .y(_in_in1__d),
        .sel(io_in_valid),
        .a(io_in_bits_in1),
        .b(_in_in1__q)
    );
    MUX_UNSIGNED #(.width(65)) u_mux_4679 (
        .y(_in_in2__d),
        .sel(io_in_valid),
        .a(_node_38),
        .b(_in_in2__q)
    );
    MUX_UNSIGNED #(.width(65)) u_mux_4680 (
        .y(_in_in3__d),
        .sel(io_in_valid),
        .a(_node_39),
        .b(_in_in3__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_4681 (
        .y(_in_ldst__d),
        .sel(io_in_valid),
        .a(io_in_bits_ldst),
        .b(_in_ldst__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_4682 (
        .y(_in_ren1__d),
        .sel(io_in_valid),
        .a(io_in_bits_ren1),
        .b(_in_ren1__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_4683 (
        .y(_in_ren2__d),
        .sel(io_in_valid),
        .a(io_in_bits_ren2),
        .b(_in_ren2__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_4684 (
        .y(_in_ren3__d),
        .sel(io_in_valid),
        .a(io_in_bits_ren3),
        .b(_in_ren3__q)
    );
    MUX_UNSIGNED #(.width(3)) u_mux_4685 (
        .y(_in_rm__d),
        .sel(io_in_valid),
        .a(io_in_bits_rm),
        .b(_in_rm__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_4686 (
        .y(_in_single__d),
        .sel(io_in_valid),
        .a(io_in_bits_single),
        .b(_in_single__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_4687 (
        .y(_in_sqrt__d),
        .sel(io_in_valid),
        .a(io_in_bits_sqrt),
        .b(_in_sqrt__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_4688 (
        .y(_in_swap12__d),
        .sel(io_in_valid),
        .a(io_in_bits_swap12),
        .b(_in_swap12__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_4689 (
        .y(_in_swap23__d),
        .sel(io_in_valid),
        .a(io_in_bits_swap23),
        .b(_in_swap23__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_4690 (
        .y(_in_toint__d),
        .sel(io_in_valid),
        .a(io_in_bits_toint),
        .b(_in_toint__q)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_4691 (
        .y(_in_typ__d),
        .sel(io_in_valid),
        .a(io_in_bits_typ),
        .b(_in_typ__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_4692 (
        .y(_in_wen__d),
        .sel(io_in_valid),
        .a(io_in_bits_wen),
        .b(_in_wen__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_4693 (
        .y(_in_wflags__d),
        .sel(io_in_valid),
        .a(io_in_bits_wflags),
        .b(_in_wflags__q)
    );
    assign io_out_bits_data = _T_226_bits_data;
    assign io_out_bits_exc = _T_226_bits_exc;
    assign io_out_valid = _T_226_valid;
    assign res_data = _fma__io_out;
    assign res_exc = _fma__io_exceptionFlags;
    assign _valid__d = io_in_valid;
endmodule //FPUFMAPipe_1
module MulAddRecFN_1(
    input clock,
    input reset,
    input [1:0] io_op,
    input [64:0] io_a,
    input [64:0] io_b,
    input [64:0] io_c,
    input [1:0] io_roundingMode,
    output [64:0] io_out,
    output [4:0] io_exceptionFlags
);
    wire _mulAddRecFN_preMul__clock;
    wire _mulAddRecFN_preMul__reset;
    wire [1:0] _mulAddRecFN_preMul__io_op;
    wire [64:0] _mulAddRecFN_preMul__io_a;
    wire [64:0] _mulAddRecFN_preMul__io_b;
    wire [64:0] _mulAddRecFN_preMul__io_c;
    wire [1:0] _mulAddRecFN_preMul__io_roundingMode;
    wire [52:0] _mulAddRecFN_preMul__io_mulAddA;
    wire [52:0] _mulAddRecFN_preMul__io_mulAddB;
    wire [105:0] _mulAddRecFN_preMul__io_mulAddC;
    wire [2:0] _mulAddRecFN_preMul__io_toPostMul_highExpA;
    wire _mulAddRecFN_preMul__io_toPostMul_isNaN_isQuietNaNA;
    wire [2:0] _mulAddRecFN_preMul__io_toPostMul_highExpB;
    wire _mulAddRecFN_preMul__io_toPostMul_isNaN_isQuietNaNB;
    wire _mulAddRecFN_preMul__io_toPostMul_signProd;
    wire _mulAddRecFN_preMul__io_toPostMul_isZeroProd;
    wire _mulAddRecFN_preMul__io_toPostMul_opSignC;
    wire [2:0] _mulAddRecFN_preMul__io_toPostMul_highExpC;
    wire _mulAddRecFN_preMul__io_toPostMul_isNaN_isQuietNaNC;
    wire _mulAddRecFN_preMul__io_toPostMul_isCDominant;
    wire _mulAddRecFN_preMul__io_toPostMul_CAlignDist_0;
    wire [7:0] _mulAddRecFN_preMul__io_toPostMul_CAlignDist;
    wire _mulAddRecFN_preMul__io_toPostMul_bit0AlignedNegSigC;
    wire [54:0] _mulAddRecFN_preMul__io_toPostMul_highAlignedNegSigC;
    wire [13:0] _mulAddRecFN_preMul__io_toPostMul_sExpSum;
    wire [1:0] _mulAddRecFN_preMul__io_toPostMul_roundingMode;
    MulAddRecFN_preMul_1 mulAddRecFN_preMul (
        .clock(_mulAddRecFN_preMul__clock),
        .reset(_mulAddRecFN_preMul__reset),
        .io_op(_mulAddRecFN_preMul__io_op),
        .io_a(_mulAddRecFN_preMul__io_a),
        .io_b(_mulAddRecFN_preMul__io_b),
        .io_c(_mulAddRecFN_preMul__io_c),
        .io_roundingMode(_mulAddRecFN_preMul__io_roundingMode),
        .io_mulAddA(_mulAddRecFN_preMul__io_mulAddA),
        .io_mulAddB(_mulAddRecFN_preMul__io_mulAddB),
        .io_mulAddC(_mulAddRecFN_preMul__io_mulAddC),
        .io_toPostMul_highExpA(_mulAddRecFN_preMul__io_toPostMul_highExpA),
        .io_toPostMul_isNaN_isQuietNaNA(_mulAddRecFN_preMul__io_toPostMul_isNaN_isQuietNaNA),
        .io_toPostMul_highExpB(_mulAddRecFN_preMul__io_toPostMul_highExpB),
        .io_toPostMul_isNaN_isQuietNaNB(_mulAddRecFN_preMul__io_toPostMul_isNaN_isQuietNaNB),
        .io_toPostMul_signProd(_mulAddRecFN_preMul__io_toPostMul_signProd),
        .io_toPostMul_isZeroProd(_mulAddRecFN_preMul__io_toPostMul_isZeroProd),
        .io_toPostMul_opSignC(_mulAddRecFN_preMul__io_toPostMul_opSignC),
        .io_toPostMul_highExpC(_mulAddRecFN_preMul__io_toPostMul_highExpC),
        .io_toPostMul_isNaN_isQuietNaNC(_mulAddRecFN_preMul__io_toPostMul_isNaN_isQuietNaNC),
        .io_toPostMul_isCDominant(_mulAddRecFN_preMul__io_toPostMul_isCDominant),
        .io_toPostMul_CAlignDist_0(_mulAddRecFN_preMul__io_toPostMul_CAlignDist_0),
        .io_toPostMul_CAlignDist(_mulAddRecFN_preMul__io_toPostMul_CAlignDist),
        .io_toPostMul_bit0AlignedNegSigC(_mulAddRecFN_preMul__io_toPostMul_bit0AlignedNegSigC),
        .io_toPostMul_highAlignedNegSigC(_mulAddRecFN_preMul__io_toPostMul_highAlignedNegSigC),
        .io_toPostMul_sExpSum(_mulAddRecFN_preMul__io_toPostMul_sExpSum),
        .io_toPostMul_roundingMode(_mulAddRecFN_preMul__io_toPostMul_roundingMode)
    );
    wire _mulAddRecFN_postMul__clock;
    wire _mulAddRecFN_postMul__reset;
    wire [2:0] _mulAddRecFN_postMul__io_fromPreMul_highExpA;
    wire _mulAddRecFN_postMul__io_fromPreMul_isNaN_isQuietNaNA;
    wire [2:0] _mulAddRecFN_postMul__io_fromPreMul_highExpB;
    wire _mulAddRecFN_postMul__io_fromPreMul_isNaN_isQuietNaNB;
    wire _mulAddRecFN_postMul__io_fromPreMul_signProd;
    wire _mulAddRecFN_postMul__io_fromPreMul_isZeroProd;
    wire _mulAddRecFN_postMul__io_fromPreMul_opSignC;
    wire [2:0] _mulAddRecFN_postMul__io_fromPreMul_highExpC;
    wire _mulAddRecFN_postMul__io_fromPreMul_isNaN_isQuietNaNC;
    wire _mulAddRecFN_postMul__io_fromPreMul_isCDominant;
    wire _mulAddRecFN_postMul__io_fromPreMul_CAlignDist_0;
    wire [7:0] _mulAddRecFN_postMul__io_fromPreMul_CAlignDist;
    wire _mulAddRecFN_postMul__io_fromPreMul_bit0AlignedNegSigC;
    wire [54:0] _mulAddRecFN_postMul__io_fromPreMul_highAlignedNegSigC;
    wire [13:0] _mulAddRecFN_postMul__io_fromPreMul_sExpSum;
    wire [1:0] _mulAddRecFN_postMul__io_fromPreMul_roundingMode;
    wire [106:0] _mulAddRecFN_postMul__io_mulAddResult;
    wire [64:0] _mulAddRecFN_postMul__io_out;
    wire [4:0] _mulAddRecFN_postMul__io_exceptionFlags;
    MulAddRecFN_postMul_1 mulAddRecFN_postMul (
        .clock(_mulAddRecFN_postMul__clock),
        .reset(_mulAddRecFN_postMul__reset),
        .io_fromPreMul_highExpA(_mulAddRecFN_postMul__io_fromPreMul_highExpA),
        .io_fromPreMul_isNaN_isQuietNaNA(_mulAddRecFN_postMul__io_fromPreMul_isNaN_isQuietNaNA),
        .io_fromPreMul_highExpB(_mulAddRecFN_postMul__io_fromPreMul_highExpB),
        .io_fromPreMul_isNaN_isQuietNaNB(_mulAddRecFN_postMul__io_fromPreMul_isNaN_isQuietNaNB),
        .io_fromPreMul_signProd(_mulAddRecFN_postMul__io_fromPreMul_signProd),
        .io_fromPreMul_isZeroProd(_mulAddRecFN_postMul__io_fromPreMul_isZeroProd),
        .io_fromPreMul_opSignC(_mulAddRecFN_postMul__io_fromPreMul_opSignC),
        .io_fromPreMul_highExpC(_mulAddRecFN_postMul__io_fromPreMul_highExpC),
        .io_fromPreMul_isNaN_isQuietNaNC(_mulAddRecFN_postMul__io_fromPreMul_isNaN_isQuietNaNC),
        .io_fromPreMul_isCDominant(_mulAddRecFN_postMul__io_fromPreMul_isCDominant),
        .io_fromPreMul_CAlignDist_0(_mulAddRecFN_postMul__io_fromPreMul_CAlignDist_0),
        .io_fromPreMul_CAlignDist(_mulAddRecFN_postMul__io_fromPreMul_CAlignDist),
        .io_fromPreMul_bit0AlignedNegSigC(_mulAddRecFN_postMul__io_fromPreMul_bit0AlignedNegSigC),
        .io_fromPreMul_highAlignedNegSigC(_mulAddRecFN_postMul__io_fromPreMul_highAlignedNegSigC),
        .io_fromPreMul_sExpSum(_mulAddRecFN_postMul__io_fromPreMul_sExpSum),
        .io_fromPreMul_roundingMode(_mulAddRecFN_postMul__io_fromPreMul_roundingMode),
        .io_mulAddResult(_mulAddRecFN_postMul__io_mulAddResult),
        .io_out(_mulAddRecFN_postMul__io_out),
        .io_exceptionFlags(_mulAddRecFN_postMul__io_exceptionFlags)
    );
    wire [105:0] _T_16;
    MUL2_UNSIGNED #(.width_a(53), .width_b(53)) u_mul2_4656 (
        .y(_T_16),
        .a(_mulAddRecFN_preMul__io_mulAddA),
        .b(_mulAddRecFN_preMul__io_mulAddB)
    );
    wire [106:0] _T_18;
    CAT #(.width_a(1), .width_b(106)) cat_4657 (
        .y(_T_18),
        .a(1'h0),
        .b(_mulAddRecFN_preMul__io_mulAddC)
    );
    wire [107:0] _T_19;
    wire [106:0] _WTEMP_641;
    PAD_UNSIGNED #(.width(106), .n(107)) u_pad_4658 (
        .y(_WTEMP_641),
        .in(_T_16)
    );
    ADD_UNSIGNED #(.width(107)) u_add_4659 (
        .y(_T_19),
        .a(_WTEMP_641),
        .b(_T_18)
    );
    wire [106:0] _T_20;
    TAIL #(.width(108), .n(1)) tail_4660 (
        .y(_T_20),
        .in(_T_19)
    );
    assign io_exceptionFlags = _mulAddRecFN_postMul__io_exceptionFlags;
    assign io_out = _mulAddRecFN_postMul__io_out;
    assign _mulAddRecFN_postMul__clock = clock;
    assign _mulAddRecFN_postMul__io_fromPreMul_CAlignDist = _mulAddRecFN_preMul__io_toPostMul_CAlignDist;
    assign _mulAddRecFN_postMul__io_fromPreMul_CAlignDist_0 = _mulAddRecFN_preMul__io_toPostMul_CAlignDist_0;
    assign _mulAddRecFN_postMul__io_fromPreMul_bit0AlignedNegSigC = _mulAddRecFN_preMul__io_toPostMul_bit0AlignedNegSigC;
    assign _mulAddRecFN_postMul__io_fromPreMul_highAlignedNegSigC = _mulAddRecFN_preMul__io_toPostMul_highAlignedNegSigC;
    assign _mulAddRecFN_postMul__io_fromPreMul_highExpA = _mulAddRecFN_preMul__io_toPostMul_highExpA;
    assign _mulAddRecFN_postMul__io_fromPreMul_highExpB = _mulAddRecFN_preMul__io_toPostMul_highExpB;
    assign _mulAddRecFN_postMul__io_fromPreMul_highExpC = _mulAddRecFN_preMul__io_toPostMul_highExpC;
    assign _mulAddRecFN_postMul__io_fromPreMul_isCDominant = _mulAddRecFN_preMul__io_toPostMul_isCDominant;
    assign _mulAddRecFN_postMul__io_fromPreMul_isNaN_isQuietNaNA = _mulAddRecFN_preMul__io_toPostMul_isNaN_isQuietNaNA;
    assign _mulAddRecFN_postMul__io_fromPreMul_isNaN_isQuietNaNB = _mulAddRecFN_preMul__io_toPostMul_isNaN_isQuietNaNB;
    assign _mulAddRecFN_postMul__io_fromPreMul_isNaN_isQuietNaNC = _mulAddRecFN_preMul__io_toPostMul_isNaN_isQuietNaNC;
    assign _mulAddRecFN_postMul__io_fromPreMul_isZeroProd = _mulAddRecFN_preMul__io_toPostMul_isZeroProd;
    assign _mulAddRecFN_postMul__io_fromPreMul_opSignC = _mulAddRecFN_preMul__io_toPostMul_opSignC;
    assign _mulAddRecFN_postMul__io_fromPreMul_roundingMode = _mulAddRecFN_preMul__io_toPostMul_roundingMode;
    assign _mulAddRecFN_postMul__io_fromPreMul_sExpSum = _mulAddRecFN_preMul__io_toPostMul_sExpSum;
    assign _mulAddRecFN_postMul__io_fromPreMul_signProd = _mulAddRecFN_preMul__io_toPostMul_signProd;
    assign _mulAddRecFN_postMul__io_mulAddResult = _T_20;
    assign _mulAddRecFN_postMul__reset = reset;
    assign _mulAddRecFN_preMul__clock = clock;
    assign _mulAddRecFN_preMul__io_a = io_a;
    assign _mulAddRecFN_preMul__io_b = io_b;
    assign _mulAddRecFN_preMul__io_c = io_c;
    assign _mulAddRecFN_preMul__io_op = io_op;
    assign _mulAddRecFN_preMul__io_roundingMode = io_roundingMode;
    assign _mulAddRecFN_preMul__reset = reset;
endmodule //MulAddRecFN_1
module MulAddRecFN_preMul_1(
    input clock,
    input reset,
    input [1:0] io_op,
    input [64:0] io_a,
    input [64:0] io_b,
    input [64:0] io_c,
    input [1:0] io_roundingMode,
    output [52:0] io_mulAddA,
    output [52:0] io_mulAddB,
    output [105:0] io_mulAddC,
    output [2:0] io_toPostMul_highExpA,
    output io_toPostMul_isNaN_isQuietNaNA,
    output [2:0] io_toPostMul_highExpB,
    output io_toPostMul_isNaN_isQuietNaNB,
    output io_toPostMul_signProd,
    output io_toPostMul_isZeroProd,
    output io_toPostMul_opSignC,
    output [2:0] io_toPostMul_highExpC,
    output io_toPostMul_isNaN_isQuietNaNC,
    output io_toPostMul_isCDominant,
    output io_toPostMul_CAlignDist_0,
    output [7:0] io_toPostMul_CAlignDist,
    output io_toPostMul_bit0AlignedNegSigC,
    output [54:0] io_toPostMul_highAlignedNegSigC,
    output [13:0] io_toPostMul_sExpSum,
    output [1:0] io_toPostMul_roundingMode
);
    wire signA;
    BITS #(.width(65), .high(64), .low(64)) bits_3493 (
        .y(signA),
        .in(io_a)
    );
    wire [11:0] expA;
    BITS #(.width(65), .high(63), .low(52)) bits_3494 (
        .y(expA),
        .in(io_a)
    );
    wire [51:0] fractA;
    BITS #(.width(65), .high(51), .low(0)) bits_3495 (
        .y(fractA),
        .in(io_a)
    );
    wire [2:0] _T_52;
    BITS #(.width(12), .high(11), .low(9)) bits_3496 (
        .y(_T_52),
        .in(expA)
    );
    wire isZeroA;
    wire [2:0] _WTEMP_479;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_3497 (
        .y(_WTEMP_479),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(3)) u_eq_3498 (
        .y(isZeroA),
        .a(_T_52),
        .b(_WTEMP_479)
    );
    wire _T_55;
    EQ_UNSIGNED #(.width(1)) u_eq_3499 (
        .y(_T_55),
        .a(isZeroA),
        .b(1'h0)
    );
    wire [52:0] sigA;
    CAT #(.width_a(1), .width_b(52)) cat_3500 (
        .y(sigA),
        .a(_T_55),
        .b(fractA)
    );
    wire signB;
    BITS #(.width(65), .high(64), .low(64)) bits_3501 (
        .y(signB),
        .in(io_b)
    );
    wire [11:0] expB;
    BITS #(.width(65), .high(63), .low(52)) bits_3502 (
        .y(expB),
        .in(io_b)
    );
    wire [51:0] fractB;
    BITS #(.width(65), .high(51), .low(0)) bits_3503 (
        .y(fractB),
        .in(io_b)
    );
    wire [2:0] _T_56;
    BITS #(.width(12), .high(11), .low(9)) bits_3504 (
        .y(_T_56),
        .in(expB)
    );
    wire isZeroB;
    wire [2:0] _WTEMP_480;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_3505 (
        .y(_WTEMP_480),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(3)) u_eq_3506 (
        .y(isZeroB),
        .a(_T_56),
        .b(_WTEMP_480)
    );
    wire _T_59;
    EQ_UNSIGNED #(.width(1)) u_eq_3507 (
        .y(_T_59),
        .a(isZeroB),
        .b(1'h0)
    );
    wire [52:0] sigB;
    CAT #(.width_a(1), .width_b(52)) cat_3508 (
        .y(sigB),
        .a(_T_59),
        .b(fractB)
    );
    wire _T_60;
    BITS #(.width(65), .high(64), .low(64)) bits_3509 (
        .y(_T_60),
        .in(io_c)
    );
    wire _T_61;
    BITS #(.width(2), .high(0), .low(0)) bits_3510 (
        .y(_T_61),
        .in(io_op)
    );
    wire opSignC;
    BITWISEXOR #(.width(1)) bitwisexor_3511 (
        .y(opSignC),
        .a(_T_60),
        .b(_T_61)
    );
    wire [11:0] expC;
    BITS #(.width(65), .high(63), .low(52)) bits_3512 (
        .y(expC),
        .in(io_c)
    );
    wire [51:0] fractC;
    BITS #(.width(65), .high(51), .low(0)) bits_3513 (
        .y(fractC),
        .in(io_c)
    );
    wire [2:0] _T_62;
    BITS #(.width(12), .high(11), .low(9)) bits_3514 (
        .y(_T_62),
        .in(expC)
    );
    wire isZeroC;
    wire [2:0] _WTEMP_481;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_3515 (
        .y(_WTEMP_481),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(3)) u_eq_3516 (
        .y(isZeroC),
        .a(_T_62),
        .b(_WTEMP_481)
    );
    wire _T_65;
    EQ_UNSIGNED #(.width(1)) u_eq_3517 (
        .y(_T_65),
        .a(isZeroC),
        .b(1'h0)
    );
    wire [52:0] sigC;
    CAT #(.width_a(1), .width_b(52)) cat_3518 (
        .y(sigC),
        .a(_T_65),
        .b(fractC)
    );
    wire _T_66;
    BITWISEXOR #(.width(1)) bitwisexor_3519 (
        .y(_T_66),
        .a(signA),
        .b(signB)
    );
    wire _T_67;
    BITS #(.width(2), .high(1), .low(1)) bits_3520 (
        .y(_T_67),
        .in(io_op)
    );
    wire signProd;
    BITWISEXOR #(.width(1)) bitwisexor_3521 (
        .y(signProd),
        .a(_T_66),
        .b(_T_67)
    );
    wire isZeroProd;
    BITWISEOR #(.width(1)) bitwiseor_3522 (
        .y(isZeroProd),
        .a(isZeroA),
        .b(isZeroB)
    );
    wire _T_68;
    BITS #(.width(12), .high(11), .low(11)) bits_3523 (
        .y(_T_68),
        .in(expB)
    );
    wire _T_70;
    EQ_UNSIGNED #(.width(1)) u_eq_3524 (
        .y(_T_70),
        .a(_T_68),
        .b(1'h0)
    );
    wire _T_71;
    BITS #(.width(1), .high(0), .low(0)) bits_3525 (
        .y(_T_71),
        .in(_T_70)
    );
    wire [2:0] _T_74;
    MUX_UNSIGNED #(.width(3)) u_mux_3526 (
        .y(_T_74),
        .sel(_T_71),
        .a(3'h7),
        .b(3'h0)
    );
    wire [10:0] _T_75;
    BITS #(.width(12), .high(10), .low(0)) bits_3527 (
        .y(_T_75),
        .in(expB)
    );
    wire [13:0] _T_76;
    CAT #(.width_a(3), .width_b(11)) cat_3528 (
        .y(_T_76),
        .a(_T_74),
        .b(_T_75)
    );
    wire [14:0] _T_77;
    wire [13:0] _WTEMP_482;
    PAD_UNSIGNED #(.width(12), .n(14)) u_pad_3529 (
        .y(_WTEMP_482),
        .in(expA)
    );
    ADD_UNSIGNED #(.width(14)) u_add_3530 (
        .y(_T_77),
        .a(_WTEMP_482),
        .b(_T_76)
    );
    wire [13:0] _T_78;
    TAIL #(.width(15), .n(1)) tail_3531 (
        .y(_T_78),
        .in(_T_77)
    );
    wire [14:0] _T_80;
    wire [13:0] _WTEMP_483;
    PAD_UNSIGNED #(.width(6), .n(14)) u_pad_3532 (
        .y(_WTEMP_483),
        .in(6'h38)
    );
    ADD_UNSIGNED #(.width(14)) u_add_3533 (
        .y(_T_80),
        .a(_T_78),
        .b(_WTEMP_483)
    );
    wire [13:0] sExpAlignedProd;
    TAIL #(.width(15), .n(1)) tail_3534 (
        .y(sExpAlignedProd),
        .in(_T_80)
    );
    wire doSubMags;
    BITWISEXOR #(.width(1)) bitwisexor_3535 (
        .y(doSubMags),
        .a(signProd),
        .b(opSignC)
    );
    wire [14:0] _T_81;
    wire [13:0] _WTEMP_484;
    PAD_UNSIGNED #(.width(12), .n(14)) u_pad_3536 (
        .y(_WTEMP_484),
        .in(expC)
    );
    SUB_UNSIGNED #(.width(14)) u_sub_3537 (
        .y(_T_81),
        .a(sExpAlignedProd),
        .b(_WTEMP_484)
    );
    wire [14:0] _T_82;
    ASUINT #(.width(15)) asuint_3538 (
        .y(_T_82),
        .in(_T_81)
    );
    wire [13:0] sNatCAlignDist;
    TAIL #(.width(15), .n(1)) tail_3539 (
        .y(sNatCAlignDist),
        .in(_T_82)
    );
    wire _T_83;
    BITS #(.width(14), .high(13), .low(13)) bits_3540 (
        .y(_T_83),
        .in(sNatCAlignDist)
    );
    wire CAlignDist_floor;
    BITWISEOR #(.width(1)) bitwiseor_3541 (
        .y(CAlignDist_floor),
        .a(isZeroProd),
        .b(_T_83)
    );
    wire [12:0] _T_84;
    BITS #(.width(14), .high(12), .low(0)) bits_3542 (
        .y(_T_84),
        .in(sNatCAlignDist)
    );
    wire _T_86;
    wire [12:0] _WTEMP_485;
    PAD_UNSIGNED #(.width(1), .n(13)) u_pad_3543 (
        .y(_WTEMP_485),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(13)) u_eq_3544 (
        .y(_T_86),
        .a(_T_84),
        .b(_WTEMP_485)
    );
    wire CAlignDist_0;
    BITWISEOR #(.width(1)) bitwiseor_3545 (
        .y(CAlignDist_0),
        .a(CAlignDist_floor),
        .b(_T_86)
    );
    wire _T_88;
    EQ_UNSIGNED #(.width(1)) u_eq_3546 (
        .y(_T_88),
        .a(isZeroC),
        .b(1'h0)
    );
    wire [12:0] _T_89;
    BITS #(.width(14), .high(12), .low(0)) bits_3547 (
        .y(_T_89),
        .in(sNatCAlignDist)
    );
    wire _T_91;
    wire [12:0] _WTEMP_486;
    PAD_UNSIGNED #(.width(6), .n(13)) u_pad_3548 (
        .y(_WTEMP_486),
        .in(6'h36)
    );
    LT_UNSIGNED #(.width(13)) u_lt_3549 (
        .y(_T_91),
        .a(_T_89),
        .b(_WTEMP_486)
    );
    wire _T_92;
    BITWISEOR #(.width(1)) bitwiseor_3550 (
        .y(_T_92),
        .a(CAlignDist_floor),
        .b(_T_91)
    );
    wire isCDominant;
    BITWISEAND #(.width(1)) bitwiseand_3551 (
        .y(isCDominant),
        .a(_T_88),
        .b(_T_92)
    );
    wire [12:0] _T_94;
    BITS #(.width(14), .high(12), .low(0)) bits_3552 (
        .y(_T_94),
        .in(sNatCAlignDist)
    );
    wire _T_96;
    wire [12:0] _WTEMP_487;
    PAD_UNSIGNED #(.width(8), .n(13)) u_pad_3553 (
        .y(_WTEMP_487),
        .in(8'hA1)
    );
    LT_UNSIGNED #(.width(13)) u_lt_3554 (
        .y(_T_96),
        .a(_T_94),
        .b(_WTEMP_487)
    );
    wire [7:0] _T_97;
    BITS #(.width(14), .high(7), .low(0)) bits_3555 (
        .y(_T_97),
        .in(sNatCAlignDist)
    );
    wire [7:0] _T_99;
    MUX_UNSIGNED #(.width(8)) u_mux_3556 (
        .y(_T_99),
        .sel(_T_96),
        .a(_T_97),
        .b(8'hA1)
    );
    wire [7:0] CAlignDist;
    wire [7:0] _WTEMP_488;
    PAD_UNSIGNED #(.width(1), .n(8)) u_pad_3557 (
        .y(_WTEMP_488),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(8)) u_mux_3558 (
        .y(CAlignDist),
        .sel(CAlignDist_floor),
        .a(_WTEMP_488),
        .b(_T_99)
    );
    wire [13:0] sExpSum;
    wire [13:0] _WTEMP_489;
    PAD_UNSIGNED #(.width(12), .n(14)) u_pad_3559 (
        .y(_WTEMP_489),
        .in(expC)
    );
    MUX_UNSIGNED #(.width(14)) u_mux_3560 (
        .y(sExpSum),
        .sel(CAlignDist_floor),
        .a(_WTEMP_489),
        .b(sExpAlignedProd)
    );
    wire _T_100;
    BITS #(.width(8), .high(7), .low(7)) bits_3561 (
        .y(_T_100),
        .in(CAlignDist)
    );
    wire [6:0] _T_101;
    BITS #(.width(8), .high(6), .low(0)) bits_3562 (
        .y(_T_101),
        .in(CAlignDist)
    );
    wire _T_102;
    BITS #(.width(7), .high(6), .low(6)) bits_3563 (
        .y(_T_102),
        .in(_T_101)
    );
    wire [5:0] _T_103;
    BITS #(.width(7), .high(5), .low(0)) bits_3564 (
        .y(_T_103),
        .in(_T_101)
    );
    wire [64:0] _T_106;
    DSHR_SIGNED #(.width_in(65), .width_n(6)) s_dshr_3565 (
        .y(_T_106),
        .in(-65'sh10000000000000000),
        .n(_T_103)
    );
    wire [32:0] _T_107;
    BITS #(.width(65), .high(63), .low(31)) bits_3566 (
        .y(_T_107),
        .in(_T_106)
    );
    wire [31:0] _T_108;
    BITS #(.width(33), .high(31), .low(0)) bits_3567 (
        .y(_T_108),
        .in(_T_107)
    );
    wire [31:0] _T_111;
    assign _T_111 = 32'hFFFF0000;
    wire [31:0] _T_112;
    assign _T_112 = 32'hFFFF;
    wire [15:0] _T_113;
    SHR_UNSIGNED #(.width(32), .n(16)) u_shr_3568 (
        .y(_T_113),
        .in(_T_108)
    );
    wire [31:0] _T_114;
    wire [31:0] _WTEMP_490;
    PAD_UNSIGNED #(.width(16), .n(32)) u_pad_3569 (
        .y(_WTEMP_490),
        .in(_T_113)
    );
    BITWISEAND #(.width(32)) bitwiseand_3570 (
        .y(_T_114),
        .a(_WTEMP_490),
        .b(_T_112)
    );
    wire [15:0] _T_115;
    BITS #(.width(32), .high(15), .low(0)) bits_3571 (
        .y(_T_115),
        .in(_T_108)
    );
    wire [31:0] _T_116;
    SHL_UNSIGNED #(.width(16), .n(16)) u_shl_3572 (
        .y(_T_116),
        .in(_T_115)
    );
    wire [31:0] _T_117;
    assign _T_117 = 32'hFFFF0000;
    wire [31:0] _T_118;
    BITWISEAND #(.width(32)) bitwiseand_3573 (
        .y(_T_118),
        .a(_T_116),
        .b(_T_117)
    );
    wire [31:0] _T_119;
    BITWISEOR #(.width(32)) bitwiseor_3574 (
        .y(_T_119),
        .a(_T_114),
        .b(_T_118)
    );
    wire [23:0] _T_120;
    assign _T_120 = 24'hFFFF;
    wire [31:0] _T_121;
    assign _T_121 = 32'hFFFF00;
    wire [31:0] _T_122;
    assign _T_122 = 32'hFF00FF;
    wire [23:0] _T_123;
    SHR_UNSIGNED #(.width(32), .n(8)) u_shr_3575 (
        .y(_T_123),
        .in(_T_119)
    );
    wire [31:0] _T_124;
    wire [31:0] _WTEMP_491;
    PAD_UNSIGNED #(.width(24), .n(32)) u_pad_3576 (
        .y(_WTEMP_491),
        .in(_T_123)
    );
    BITWISEAND #(.width(32)) bitwiseand_3577 (
        .y(_T_124),
        .a(_WTEMP_491),
        .b(_T_122)
    );
    wire [23:0] _T_125;
    BITS #(.width(32), .high(23), .low(0)) bits_3578 (
        .y(_T_125),
        .in(_T_119)
    );
    wire [31:0] _T_126;
    SHL_UNSIGNED #(.width(24), .n(8)) u_shl_3579 (
        .y(_T_126),
        .in(_T_125)
    );
    wire [31:0] _T_127;
    assign _T_127 = 32'hFF00FF00;
    wire [31:0] _T_128;
    BITWISEAND #(.width(32)) bitwiseand_3580 (
        .y(_T_128),
        .a(_T_126),
        .b(_T_127)
    );
    wire [31:0] _T_129;
    BITWISEOR #(.width(32)) bitwiseor_3581 (
        .y(_T_129),
        .a(_T_124),
        .b(_T_128)
    );
    wire [27:0] _T_130;
    assign _T_130 = 28'hFF00FF;
    wire [31:0] _T_131;
    assign _T_131 = 32'hFF00FF0;
    wire [31:0] _T_132;
    assign _T_132 = 32'hF0F0F0F;
    wire [27:0] _T_133;
    SHR_UNSIGNED #(.width(32), .n(4)) u_shr_3582 (
        .y(_T_133),
        .in(_T_129)
    );
    wire [31:0] _T_134;
    wire [31:0] _WTEMP_492;
    PAD_UNSIGNED #(.width(28), .n(32)) u_pad_3583 (
        .y(_WTEMP_492),
        .in(_T_133)
    );
    BITWISEAND #(.width(32)) bitwiseand_3584 (
        .y(_T_134),
        .a(_WTEMP_492),
        .b(_T_132)
    );
    wire [27:0] _T_135;
    BITS #(.width(32), .high(27), .low(0)) bits_3585 (
        .y(_T_135),
        .in(_T_129)
    );
    wire [31:0] _T_136;
    SHL_UNSIGNED #(.width(28), .n(4)) u_shl_3586 (
        .y(_T_136),
        .in(_T_135)
    );
    wire [31:0] _T_137;
    assign _T_137 = 32'hF0F0F0F0;
    wire [31:0] _T_138;
    BITWISEAND #(.width(32)) bitwiseand_3587 (
        .y(_T_138),
        .a(_T_136),
        .b(_T_137)
    );
    wire [31:0] _T_139;
    BITWISEOR #(.width(32)) bitwiseor_3588 (
        .y(_T_139),
        .a(_T_134),
        .b(_T_138)
    );
    wire [29:0] _T_140;
    assign _T_140 = 30'hF0F0F0F;
    wire [31:0] _T_141;
    assign _T_141 = 32'h3C3C3C3C;
    wire [31:0] _T_142;
    assign _T_142 = 32'h33333333;
    wire [29:0] _T_143;
    SHR_UNSIGNED #(.width(32), .n(2)) u_shr_3589 (
        .y(_T_143),
        .in(_T_139)
    );
    wire [31:0] _T_144;
    wire [31:0] _WTEMP_493;
    PAD_UNSIGNED #(.width(30), .n(32)) u_pad_3590 (
        .y(_WTEMP_493),
        .in(_T_143)
    );
    BITWISEAND #(.width(32)) bitwiseand_3591 (
        .y(_T_144),
        .a(_WTEMP_493),
        .b(_T_142)
    );
    wire [29:0] _T_145;
    BITS #(.width(32), .high(29), .low(0)) bits_3592 (
        .y(_T_145),
        .in(_T_139)
    );
    wire [31:0] _T_146;
    SHL_UNSIGNED #(.width(30), .n(2)) u_shl_3593 (
        .y(_T_146),
        .in(_T_145)
    );
    wire [31:0] _T_147;
    assign _T_147 = 32'hCCCCCCCC;
    wire [31:0] _T_148;
    BITWISEAND #(.width(32)) bitwiseand_3594 (
        .y(_T_148),
        .a(_T_146),
        .b(_T_147)
    );
    wire [31:0] _T_149;
    BITWISEOR #(.width(32)) bitwiseor_3595 (
        .y(_T_149),
        .a(_T_144),
        .b(_T_148)
    );
    wire [30:0] _T_150;
    assign _T_150 = 31'h33333333;
    wire [31:0] _T_151;
    assign _T_151 = 32'h66666666;
    wire [31:0] _T_152;
    assign _T_152 = 32'h55555555;
    wire [30:0] _T_153;
    SHR_UNSIGNED #(.width(32), .n(1)) u_shr_3596 (
        .y(_T_153),
        .in(_T_149)
    );
    wire [31:0] _T_154;
    wire [31:0] _WTEMP_494;
    PAD_UNSIGNED #(.width(31), .n(32)) u_pad_3597 (
        .y(_WTEMP_494),
        .in(_T_153)
    );
    BITWISEAND #(.width(32)) bitwiseand_3598 (
        .y(_T_154),
        .a(_WTEMP_494),
        .b(_T_152)
    );
    wire [30:0] _T_155;
    BITS #(.width(32), .high(30), .low(0)) bits_3599 (
        .y(_T_155),
        .in(_T_149)
    );
    wire [31:0] _T_156;
    SHL_UNSIGNED #(.width(31), .n(1)) u_shl_3600 (
        .y(_T_156),
        .in(_T_155)
    );
    wire [31:0] _T_157;
    assign _T_157 = 32'hAAAAAAAA;
    wire [31:0] _T_158;
    BITWISEAND #(.width(32)) bitwiseand_3601 (
        .y(_T_158),
        .a(_T_156),
        .b(_T_157)
    );
    wire [31:0] _T_159;
    BITWISEOR #(.width(32)) bitwiseor_3602 (
        .y(_T_159),
        .a(_T_154),
        .b(_T_158)
    );
    wire _T_160;
    BITS #(.width(33), .high(32), .low(32)) bits_3603 (
        .y(_T_160),
        .in(_T_107)
    );
    wire [32:0] _T_161;
    CAT #(.width_a(32), .width_b(1)) cat_3604 (
        .y(_T_161),
        .a(_T_159),
        .b(_T_160)
    );
    wire [32:0] _T_162;
    BITWISENOT #(.width(33)) bitwisenot_3605 (
        .y(_T_162),
        .in(_T_161)
    );
    wire [32:0] _T_163;
    wire [32:0] _WTEMP_495;
    PAD_UNSIGNED #(.width(1), .n(33)) u_pad_3606 (
        .y(_WTEMP_495),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(33)) u_mux_3607 (
        .y(_T_163),
        .sel(_T_102),
        .a(_WTEMP_495),
        .b(_T_162)
    );
    wire [32:0] _T_164;
    BITWISENOT #(.width(33)) bitwisenot_3608 (
        .y(_T_164),
        .in(_T_163)
    );
    wire [52:0] _T_166;
    CAT #(.width_a(33), .width_b(20)) cat_3609 (
        .y(_T_166),
        .a(_T_164),
        .b(20'hFFFFF)
    );
    wire _T_167;
    BITS #(.width(7), .high(6), .low(6)) bits_3610 (
        .y(_T_167),
        .in(_T_101)
    );
    wire [5:0] _T_168;
    BITS #(.width(7), .high(5), .low(0)) bits_3611 (
        .y(_T_168),
        .in(_T_101)
    );
    wire [64:0] _T_170;
    DSHR_SIGNED #(.width_in(65), .width_n(6)) s_dshr_3612 (
        .y(_T_170),
        .in(-65'sh10000000000000000),
        .n(_T_168)
    );
    wire [19:0] _T_171;
    BITS #(.width(65), .high(19), .low(0)) bits_3613 (
        .y(_T_171),
        .in(_T_170)
    );
    wire [15:0] _T_172;
    BITS #(.width(20), .high(15), .low(0)) bits_3614 (
        .y(_T_172),
        .in(_T_171)
    );
    wire [15:0] _T_175;
    assign _T_175 = 16'hFF00;
    wire [15:0] _T_176;
    assign _T_176 = 16'hFF;
    wire [7:0] _T_177;
    SHR_UNSIGNED #(.width(16), .n(8)) u_shr_3615 (
        .y(_T_177),
        .in(_T_172)
    );
    wire [15:0] _T_178;
    wire [15:0] _WTEMP_496;
    PAD_UNSIGNED #(.width(8), .n(16)) u_pad_3616 (
        .y(_WTEMP_496),
        .in(_T_177)
    );
    BITWISEAND #(.width(16)) bitwiseand_3617 (
        .y(_T_178),
        .a(_WTEMP_496),
        .b(_T_176)
    );
    wire [7:0] _T_179;
    BITS #(.width(16), .high(7), .low(0)) bits_3618 (
        .y(_T_179),
        .in(_T_172)
    );
    wire [15:0] _T_180;
    SHL_UNSIGNED #(.width(8), .n(8)) u_shl_3619 (
        .y(_T_180),
        .in(_T_179)
    );
    wire [15:0] _T_181;
    assign _T_181 = 16'hFF00;
    wire [15:0] _T_182;
    BITWISEAND #(.width(16)) bitwiseand_3620 (
        .y(_T_182),
        .a(_T_180),
        .b(_T_181)
    );
    wire [15:0] _T_183;
    BITWISEOR #(.width(16)) bitwiseor_3621 (
        .y(_T_183),
        .a(_T_178),
        .b(_T_182)
    );
    wire [11:0] _T_184;
    assign _T_184 = 12'hFF;
    wire [15:0] _T_185;
    assign _T_185 = 16'hFF0;
    wire [15:0] _T_186;
    assign _T_186 = 16'hF0F;
    wire [11:0] _T_187;
    SHR_UNSIGNED #(.width(16), .n(4)) u_shr_3622 (
        .y(_T_187),
        .in(_T_183)
    );
    wire [15:0] _T_188;
    wire [15:0] _WTEMP_497;
    PAD_UNSIGNED #(.width(12), .n(16)) u_pad_3623 (
        .y(_WTEMP_497),
        .in(_T_187)
    );
    BITWISEAND #(.width(16)) bitwiseand_3624 (
        .y(_T_188),
        .a(_WTEMP_497),
        .b(_T_186)
    );
    wire [11:0] _T_189;
    BITS #(.width(16), .high(11), .low(0)) bits_3625 (
        .y(_T_189),
        .in(_T_183)
    );
    wire [15:0] _T_190;
    SHL_UNSIGNED #(.width(12), .n(4)) u_shl_3626 (
        .y(_T_190),
        .in(_T_189)
    );
    wire [15:0] _T_191;
    assign _T_191 = 16'hF0F0;
    wire [15:0] _T_192;
    BITWISEAND #(.width(16)) bitwiseand_3627 (
        .y(_T_192),
        .a(_T_190),
        .b(_T_191)
    );
    wire [15:0] _T_193;
    BITWISEOR #(.width(16)) bitwiseor_3628 (
        .y(_T_193),
        .a(_T_188),
        .b(_T_192)
    );
    wire [13:0] _T_194;
    assign _T_194 = 14'hF0F;
    wire [15:0] _T_195;
    assign _T_195 = 16'h3C3C;
    wire [15:0] _T_196;
    assign _T_196 = 16'h3333;
    wire [13:0] _T_197;
    SHR_UNSIGNED #(.width(16), .n(2)) u_shr_3629 (
        .y(_T_197),
        .in(_T_193)
    );
    wire [15:0] _T_198;
    wire [15:0] _WTEMP_498;
    PAD_UNSIGNED #(.width(14), .n(16)) u_pad_3630 (
        .y(_WTEMP_498),
        .in(_T_197)
    );
    BITWISEAND #(.width(16)) bitwiseand_3631 (
        .y(_T_198),
        .a(_WTEMP_498),
        .b(_T_196)
    );
    wire [13:0] _T_199;
    BITS #(.width(16), .high(13), .low(0)) bits_3632 (
        .y(_T_199),
        .in(_T_193)
    );
    wire [15:0] _T_200;
    SHL_UNSIGNED #(.width(14), .n(2)) u_shl_3633 (
        .y(_T_200),
        .in(_T_199)
    );
    wire [15:0] _T_201;
    assign _T_201 = 16'hCCCC;
    wire [15:0] _T_202;
    BITWISEAND #(.width(16)) bitwiseand_3634 (
        .y(_T_202),
        .a(_T_200),
        .b(_T_201)
    );
    wire [15:0] _T_203;
    BITWISEOR #(.width(16)) bitwiseor_3635 (
        .y(_T_203),
        .a(_T_198),
        .b(_T_202)
    );
    wire [14:0] _T_204;
    assign _T_204 = 15'h3333;
    wire [15:0] _T_205;
    assign _T_205 = 16'h6666;
    wire [15:0] _T_206;
    assign _T_206 = 16'h5555;
    wire [14:0] _T_207;
    SHR_UNSIGNED #(.width(16), .n(1)) u_shr_3636 (
        .y(_T_207),
        .in(_T_203)
    );
    wire [15:0] _T_208;
    wire [15:0] _WTEMP_499;
    PAD_UNSIGNED #(.width(15), .n(16)) u_pad_3637 (
        .y(_WTEMP_499),
        .in(_T_207)
    );
    BITWISEAND #(.width(16)) bitwiseand_3638 (
        .y(_T_208),
        .a(_WTEMP_499),
        .b(_T_206)
    );
    wire [14:0] _T_209;
    BITS #(.width(16), .high(14), .low(0)) bits_3639 (
        .y(_T_209),
        .in(_T_203)
    );
    wire [15:0] _T_210;
    SHL_UNSIGNED #(.width(15), .n(1)) u_shl_3640 (
        .y(_T_210),
        .in(_T_209)
    );
    wire [15:0] _T_211;
    assign _T_211 = 16'hAAAA;
    wire [15:0] _T_212;
    BITWISEAND #(.width(16)) bitwiseand_3641 (
        .y(_T_212),
        .a(_T_210),
        .b(_T_211)
    );
    wire [15:0] _T_213;
    BITWISEOR #(.width(16)) bitwiseor_3642 (
        .y(_T_213),
        .a(_T_208),
        .b(_T_212)
    );
    wire [3:0] _T_214;
    BITS #(.width(20), .high(19), .low(16)) bits_3643 (
        .y(_T_214),
        .in(_T_171)
    );
    wire [1:0] _T_215;
    BITS #(.width(4), .high(1), .low(0)) bits_3644 (
        .y(_T_215),
        .in(_T_214)
    );
    wire _T_216;
    BITS #(.width(2), .high(0), .low(0)) bits_3645 (
        .y(_T_216),
        .in(_T_215)
    );
    wire _T_217;
    BITS #(.width(2), .high(1), .low(1)) bits_3646 (
        .y(_T_217),
        .in(_T_215)
    );
    wire [1:0] _T_218;
    CAT #(.width_a(1), .width_b(1)) cat_3647 (
        .y(_T_218),
        .a(_T_216),
        .b(_T_217)
    );
    wire [1:0] _T_219;
    BITS #(.width(4), .high(3), .low(2)) bits_3648 (
        .y(_T_219),
        .in(_T_214)
    );
    wire _T_220;
    BITS #(.width(2), .high(0), .low(0)) bits_3649 (
        .y(_T_220),
        .in(_T_219)
    );
    wire _T_221;
    BITS #(.width(2), .high(1), .low(1)) bits_3650 (
        .y(_T_221),
        .in(_T_219)
    );
    wire [1:0] _T_222;
    CAT #(.width_a(1), .width_b(1)) cat_3651 (
        .y(_T_222),
        .a(_T_220),
        .b(_T_221)
    );
    wire [3:0] _T_223;
    CAT #(.width_a(2), .width_b(2)) cat_3652 (
        .y(_T_223),
        .a(_T_218),
        .b(_T_222)
    );
    wire [19:0] _T_224;
    CAT #(.width_a(16), .width_b(4)) cat_3653 (
        .y(_T_224),
        .a(_T_213),
        .b(_T_223)
    );
    wire [19:0] _T_226;
    wire [19:0] _WTEMP_500;
    PAD_UNSIGNED #(.width(1), .n(20)) u_pad_3654 (
        .y(_WTEMP_500),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(20)) u_mux_3655 (
        .y(_T_226),
        .sel(_T_167),
        .a(_T_224),
        .b(_WTEMP_500)
    );
    wire [52:0] CExtraMask;
    wire [52:0] _WTEMP_501;
    PAD_UNSIGNED #(.width(20), .n(53)) u_pad_3656 (
        .y(_WTEMP_501),
        .in(_T_226)
    );
    MUX_UNSIGNED #(.width(53)) u_mux_3657 (
        .y(CExtraMask),
        .sel(_T_100),
        .a(_T_166),
        .b(_WTEMP_501)
    );
    wire [52:0] _T_227;
    BITWISENOT #(.width(53)) bitwisenot_3658 (
        .y(_T_227),
        .in(sigC)
    );
    wire [52:0] negSigC;
    MUX_UNSIGNED #(.width(53)) u_mux_3659 (
        .y(negSigC),
        .sel(doSubMags),
        .a(_T_227),
        .b(sigC)
    );
    wire _T_228;
    BITS #(.width(1), .high(0), .low(0)) bits_3660 (
        .y(_T_228),
        .in(doSubMags)
    );
    wire [107:0] _T_231;
    MUX_UNSIGNED #(.width(108)) u_mux_3661 (
        .y(_T_231),
        .sel(_T_228),
        .a(108'hFFFFFFFFFFFFFFFFFFFFFFFFFFF),
        .b(108'h0)
    );
    wire [53:0] _T_232;
    CAT #(.width_a(1), .width_b(53)) cat_3662 (
        .y(_T_232),
        .a(doSubMags),
        .b(negSigC)
    );
    wire [161:0] _T_233;
    CAT #(.width_a(54), .width_b(108)) cat_3663 (
        .y(_T_233),
        .a(_T_232),
        .b(_T_231)
    );
    wire [161:0] _T_234;
    ASSINT #(.width(162)) assint_3664 (
        .y(_T_234),
        .in(_T_233)
    );
    wire [161:0] _T_235;
    DSHR_SIGNED #(.width_in(162), .width_n(8)) s_dshr_3665 (
        .y(_T_235),
        .in(_T_234),
        .n(CAlignDist)
    );
    wire [52:0] _T_236;
    BITWISEAND #(.width(53)) bitwiseand_3666 (
        .y(_T_236),
        .a(sigC),
        .b(CExtraMask)
    );
    wire _T_238;
    wire [52:0] _WTEMP_502;
    PAD_UNSIGNED #(.width(1), .n(53)) u_pad_3667 (
        .y(_WTEMP_502),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(53)) u_neq_3668 (
        .y(_T_238),
        .a(_T_236),
        .b(_WTEMP_502)
    );
    wire _T_239;
    BITWISEXOR #(.width(1)) bitwisexor_3669 (
        .y(_T_239),
        .a(_T_238),
        .b(doSubMags)
    );
    wire [161:0] _T_240;
    ASUINT #(.width(162)) asuint_3670 (
        .y(_T_240),
        .in(_T_235)
    );
    wire [162:0] _T_241;
    CAT #(.width_a(162), .width_b(1)) cat_3671 (
        .y(_T_241),
        .a(_T_240),
        .b(_T_239)
    );
    wire [161:0] alignedNegSigC;
    BITS #(.width(163), .high(161), .low(0)) bits_3672 (
        .y(alignedNegSigC),
        .in(_T_241)
    );
    wire [105:0] _T_242;
    BITS #(.width(162), .high(106), .low(1)) bits_3673 (
        .y(_T_242),
        .in(alignedNegSigC)
    );
    wire [2:0] _T_243;
    BITS #(.width(12), .high(11), .low(9)) bits_3674 (
        .y(_T_243),
        .in(expA)
    );
    wire _T_244;
    BITS #(.width(52), .high(51), .low(51)) bits_3675 (
        .y(_T_244),
        .in(fractA)
    );
    wire [2:0] _T_245;
    BITS #(.width(12), .high(11), .low(9)) bits_3676 (
        .y(_T_245),
        .in(expB)
    );
    wire _T_246;
    BITS #(.width(52), .high(51), .low(51)) bits_3677 (
        .y(_T_246),
        .in(fractB)
    );
    wire [2:0] _T_247;
    BITS #(.width(12), .high(11), .low(9)) bits_3678 (
        .y(_T_247),
        .in(expC)
    );
    wire _T_248;
    BITS #(.width(52), .high(51), .low(51)) bits_3679 (
        .y(_T_248),
        .in(fractC)
    );
    wire _T_249;
    BITS #(.width(162), .high(0), .low(0)) bits_3680 (
        .y(_T_249),
        .in(alignedNegSigC)
    );
    wire [54:0] _T_250;
    BITS #(.width(162), .high(161), .low(107)) bits_3681 (
        .y(_T_250),
        .in(alignedNegSigC)
    );
    assign io_mulAddA = sigA;
    assign io_mulAddB = sigB;
    assign io_mulAddC = _T_242;
    assign io_toPostMul_CAlignDist = CAlignDist;
    assign io_toPostMul_CAlignDist_0 = CAlignDist_0;
    assign io_toPostMul_bit0AlignedNegSigC = _T_249;
    assign io_toPostMul_highAlignedNegSigC = _T_250;
    assign io_toPostMul_highExpA = _T_243;
    assign io_toPostMul_highExpB = _T_245;
    assign io_toPostMul_highExpC = _T_247;
    assign io_toPostMul_isCDominant = isCDominant;
    assign io_toPostMul_isNaN_isQuietNaNA = _T_244;
    assign io_toPostMul_isNaN_isQuietNaNB = _T_246;
    assign io_toPostMul_isNaN_isQuietNaNC = _T_248;
    assign io_toPostMul_isZeroProd = isZeroProd;
    assign io_toPostMul_opSignC = opSignC;
    assign io_toPostMul_roundingMode = io_roundingMode;
    assign io_toPostMul_sExpSum = sExpSum;
    assign io_toPostMul_signProd = signProd;
endmodule //MulAddRecFN_preMul_1
module MulAddRecFN_postMul_1(
    input clock,
    input reset,
    input [2:0] io_fromPreMul_highExpA,
    input io_fromPreMul_isNaN_isQuietNaNA,
    input [2:0] io_fromPreMul_highExpB,
    input io_fromPreMul_isNaN_isQuietNaNB,
    input io_fromPreMul_signProd,
    input io_fromPreMul_isZeroProd,
    input io_fromPreMul_opSignC,
    input [2:0] io_fromPreMul_highExpC,
    input io_fromPreMul_isNaN_isQuietNaNC,
    input io_fromPreMul_isCDominant,
    input io_fromPreMul_CAlignDist_0,
    input [7:0] io_fromPreMul_CAlignDist,
    input io_fromPreMul_bit0AlignedNegSigC,
    input [54:0] io_fromPreMul_highAlignedNegSigC,
    input [13:0] io_fromPreMul_sExpSum,
    input [1:0] io_fromPreMul_roundingMode,
    input [106:0] io_mulAddResult,
    output [64:0] io_out,
    output [4:0] io_exceptionFlags
);
    wire isZeroA;
    wire [2:0] _WTEMP_503;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_3682 (
        .y(_WTEMP_503),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(3)) u_eq_3683 (
        .y(isZeroA),
        .a(io_fromPreMul_highExpA),
        .b(_WTEMP_503)
    );
    wire [1:0] _T_43;
    BITS #(.width(3), .high(2), .low(1)) bits_3684 (
        .y(_T_43),
        .in(io_fromPreMul_highExpA)
    );
    wire isSpecialA;
    EQ_UNSIGNED #(.width(2)) u_eq_3685 (
        .y(isSpecialA),
        .a(_T_43),
        .b(2'h3)
    );
    wire _T_45;
    BITS #(.width(3), .high(0), .low(0)) bits_3686 (
        .y(_T_45),
        .in(io_fromPreMul_highExpA)
    );
    wire _T_47;
    EQ_UNSIGNED #(.width(1)) u_eq_3687 (
        .y(_T_47),
        .a(_T_45),
        .b(1'h0)
    );
    wire isInfA;
    BITWISEAND #(.width(1)) bitwiseand_3688 (
        .y(isInfA),
        .a(isSpecialA),
        .b(_T_47)
    );
    wire _T_48;
    BITS #(.width(3), .high(0), .low(0)) bits_3689 (
        .y(_T_48),
        .in(io_fromPreMul_highExpA)
    );
    wire isNaNA;
    BITWISEAND #(.width(1)) bitwiseand_3690 (
        .y(isNaNA),
        .a(isSpecialA),
        .b(_T_48)
    );
    wire _T_50;
    EQ_UNSIGNED #(.width(1)) u_eq_3691 (
        .y(_T_50),
        .a(io_fromPreMul_isNaN_isQuietNaNA),
        .b(1'h0)
    );
    wire isSigNaNA;
    BITWISEAND #(.width(1)) bitwiseand_3692 (
        .y(isSigNaNA),
        .a(isNaNA),
        .b(_T_50)
    );
    wire isZeroB;
    wire [2:0] _WTEMP_504;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_3693 (
        .y(_WTEMP_504),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(3)) u_eq_3694 (
        .y(isZeroB),
        .a(io_fromPreMul_highExpB),
        .b(_WTEMP_504)
    );
    wire [1:0] _T_52;
    BITS #(.width(3), .high(2), .low(1)) bits_3695 (
        .y(_T_52),
        .in(io_fromPreMul_highExpB)
    );
    wire isSpecialB;
    EQ_UNSIGNED #(.width(2)) u_eq_3696 (
        .y(isSpecialB),
        .a(_T_52),
        .b(2'h3)
    );
    wire _T_54;
    BITS #(.width(3), .high(0), .low(0)) bits_3697 (
        .y(_T_54),
        .in(io_fromPreMul_highExpB)
    );
    wire _T_56;
    EQ_UNSIGNED #(.width(1)) u_eq_3698 (
        .y(_T_56),
        .a(_T_54),
        .b(1'h0)
    );
    wire isInfB;
    BITWISEAND #(.width(1)) bitwiseand_3699 (
        .y(isInfB),
        .a(isSpecialB),
        .b(_T_56)
    );
    wire _T_57;
    BITS #(.width(3), .high(0), .low(0)) bits_3700 (
        .y(_T_57),
        .in(io_fromPreMul_highExpB)
    );
    wire isNaNB;
    BITWISEAND #(.width(1)) bitwiseand_3701 (
        .y(isNaNB),
        .a(isSpecialB),
        .b(_T_57)
    );
    wire _T_59;
    EQ_UNSIGNED #(.width(1)) u_eq_3702 (
        .y(_T_59),
        .a(io_fromPreMul_isNaN_isQuietNaNB),
        .b(1'h0)
    );
    wire isSigNaNB;
    BITWISEAND #(.width(1)) bitwiseand_3703 (
        .y(isSigNaNB),
        .a(isNaNB),
        .b(_T_59)
    );
    wire isZeroC;
    wire [2:0] _WTEMP_505;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_3704 (
        .y(_WTEMP_505),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(3)) u_eq_3705 (
        .y(isZeroC),
        .a(io_fromPreMul_highExpC),
        .b(_WTEMP_505)
    );
    wire [1:0] _T_61;
    BITS #(.width(3), .high(2), .low(1)) bits_3706 (
        .y(_T_61),
        .in(io_fromPreMul_highExpC)
    );
    wire isSpecialC;
    EQ_UNSIGNED #(.width(2)) u_eq_3707 (
        .y(isSpecialC),
        .a(_T_61),
        .b(2'h3)
    );
    wire _T_63;
    BITS #(.width(3), .high(0), .low(0)) bits_3708 (
        .y(_T_63),
        .in(io_fromPreMul_highExpC)
    );
    wire _T_65;
    EQ_UNSIGNED #(.width(1)) u_eq_3709 (
        .y(_T_65),
        .a(_T_63),
        .b(1'h0)
    );
    wire isInfC;
    BITWISEAND #(.width(1)) bitwiseand_3710 (
        .y(isInfC),
        .a(isSpecialC),
        .b(_T_65)
    );
    wire _T_66;
    BITS #(.width(3), .high(0), .low(0)) bits_3711 (
        .y(_T_66),
        .in(io_fromPreMul_highExpC)
    );
    wire isNaNC;
    BITWISEAND #(.width(1)) bitwiseand_3712 (
        .y(isNaNC),
        .a(isSpecialC),
        .b(_T_66)
    );
    wire _T_68;
    EQ_UNSIGNED #(.width(1)) u_eq_3713 (
        .y(_T_68),
        .a(io_fromPreMul_isNaN_isQuietNaNC),
        .b(1'h0)
    );
    wire isSigNaNC;
    BITWISEAND #(.width(1)) bitwiseand_3714 (
        .y(isSigNaNC),
        .a(isNaNC),
        .b(_T_68)
    );
    wire roundingMode_nearest_even;
    EQ_UNSIGNED #(.width(2)) u_eq_3715 (
        .y(roundingMode_nearest_even),
        .a(io_fromPreMul_roundingMode),
        .b(2'h0)
    );
    wire roundingMode_minMag;
    EQ_UNSIGNED #(.width(2)) u_eq_3716 (
        .y(roundingMode_minMag),
        .a(io_fromPreMul_roundingMode),
        .b(2'h1)
    );
    wire roundingMode_min;
    EQ_UNSIGNED #(.width(2)) u_eq_3717 (
        .y(roundingMode_min),
        .a(io_fromPreMul_roundingMode),
        .b(2'h2)
    );
    wire roundingMode_max;
    EQ_UNSIGNED #(.width(2)) u_eq_3718 (
        .y(roundingMode_max),
        .a(io_fromPreMul_roundingMode),
        .b(2'h3)
    );
    wire signZeroNotEqOpSigns;
    MUX_UNSIGNED #(.width(1)) u_mux_3719 (
        .y(signZeroNotEqOpSigns),
        .sel(roundingMode_min),
        .a(1'h1),
        .b(1'h0)
    );
    wire doSubMags;
    BITWISEXOR #(.width(1)) bitwisexor_3720 (
        .y(doSubMags),
        .a(io_fromPreMul_signProd),
        .b(io_fromPreMul_opSignC)
    );
    wire _T_71;
    BITS #(.width(107), .high(106), .low(106)) bits_3721 (
        .y(_T_71),
        .in(io_mulAddResult)
    );
    wire [55:0] _T_73;
    wire [54:0] _WTEMP_506;
    PAD_UNSIGNED #(.width(1), .n(55)) u_pad_3722 (
        .y(_WTEMP_506),
        .in(1'h1)
    );
    ADD_UNSIGNED #(.width(55)) u_add_3723 (
        .y(_T_73),
        .a(io_fromPreMul_highAlignedNegSigC),
        .b(_WTEMP_506)
    );
    wire [54:0] _T_74;
    TAIL #(.width(56), .n(1)) tail_3724 (
        .y(_T_74),
        .in(_T_73)
    );
    wire [54:0] _T_75;
    MUX_UNSIGNED #(.width(55)) u_mux_3725 (
        .y(_T_75),
        .sel(_T_71),
        .a(_T_74),
        .b(io_fromPreMul_highAlignedNegSigC)
    );
    wire [105:0] _T_76;
    BITS #(.width(107), .high(105), .low(0)) bits_3726 (
        .y(_T_76),
        .in(io_mulAddResult)
    );
    wire [160:0] _T_77;
    CAT #(.width_a(55), .width_b(106)) cat_3727 (
        .y(_T_77),
        .a(_T_75),
        .b(_T_76)
    );
    wire [161:0] sigSum;
    CAT #(.width_a(161), .width_b(1)) cat_3728 (
        .y(sigSum),
        .a(_T_77),
        .b(io_fromPreMul_bit0AlignedNegSigC)
    );
    wire [107:0] _T_79;
    BITS #(.width(162), .high(108), .low(1)) bits_3729 (
        .y(_T_79),
        .in(sigSum)
    );
    wire [107:0] _T_80;
    BITWISEXOR #(.width(108)) bitwisexor_3730 (
        .y(_T_80),
        .a(108'h0),
        .b(_T_79)
    );
    wire [107:0] _T_81;
    BITWISEOR #(.width(108)) bitwiseor_3731 (
        .y(_T_81),
        .a(108'h0),
        .b(_T_79)
    );
    wire [108:0] _T_82;
    SHL_UNSIGNED #(.width(108), .n(1)) u_shl_3732 (
        .y(_T_82),
        .in(_T_81)
    );
    wire [108:0] _T_83;
    wire [108:0] _WTEMP_507;
    PAD_UNSIGNED #(.width(108), .n(109)) u_pad_3733 (
        .y(_WTEMP_507),
        .in(_T_80)
    );
    BITWISEXOR #(.width(109)) bitwisexor_3734 (
        .y(_T_83),
        .a(_WTEMP_507),
        .b(_T_82)
    );
    wire [107:0] _T_85;
    BITS #(.width(109), .high(107), .low(0)) bits_3735 (
        .y(_T_85),
        .in(_T_83)
    );
    wire [43:0] _T_86;
    BITS #(.width(108), .high(107), .low(64)) bits_3736 (
        .y(_T_86),
        .in(_T_85)
    );
    wire [63:0] _T_87;
    BITS #(.width(108), .high(63), .low(0)) bits_3737 (
        .y(_T_87),
        .in(_T_85)
    );
    wire _T_89;
    wire [43:0] _WTEMP_508;
    PAD_UNSIGNED #(.width(1), .n(44)) u_pad_3738 (
        .y(_WTEMP_508),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(44)) u_neq_3739 (
        .y(_T_89),
        .a(_T_86),
        .b(_WTEMP_508)
    );
    wire [11:0] _T_90;
    BITS #(.width(44), .high(43), .low(32)) bits_3740 (
        .y(_T_90),
        .in(_T_86)
    );
    wire [31:0] _T_91;
    BITS #(.width(44), .high(31), .low(0)) bits_3741 (
        .y(_T_91),
        .in(_T_86)
    );
    wire _T_93;
    wire [11:0] _WTEMP_509;
    PAD_UNSIGNED #(.width(1), .n(12)) u_pad_3742 (
        .y(_WTEMP_509),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(12)) u_neq_3743 (
        .y(_T_93),
        .a(_T_90),
        .b(_WTEMP_509)
    );
    wire [3:0] _T_94;
    BITS #(.width(12), .high(11), .low(8)) bits_3744 (
        .y(_T_94),
        .in(_T_90)
    );
    wire [7:0] _T_95;
    BITS #(.width(12), .high(7), .low(0)) bits_3745 (
        .y(_T_95),
        .in(_T_90)
    );
    wire _T_97;
    wire [3:0] _WTEMP_510;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_3746 (
        .y(_WTEMP_510),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_3747 (
        .y(_T_97),
        .a(_T_94),
        .b(_WTEMP_510)
    );
    wire _T_98;
    BITS #(.width(4), .high(3), .low(3)) bits_3748 (
        .y(_T_98),
        .in(_T_94)
    );
    wire _T_100;
    BITS #(.width(4), .high(2), .low(2)) bits_3749 (
        .y(_T_100),
        .in(_T_94)
    );
    wire _T_102;
    BITS #(.width(4), .high(1), .low(1)) bits_3750 (
        .y(_T_102),
        .in(_T_94)
    );
    wire [1:0] _T_103;
    wire [1:0] _WTEMP_511;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_3751 (
        .y(_WTEMP_511),
        .in(_T_102)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_3752 (
        .y(_T_103),
        .sel(_T_100),
        .a(2'h2),
        .b(_WTEMP_511)
    );
    wire [1:0] _T_104;
    MUX_UNSIGNED #(.width(2)) u_mux_3753 (
        .y(_T_104),
        .sel(_T_98),
        .a(2'h3),
        .b(_T_103)
    );
    wire [3:0] _T_105;
    BITS #(.width(8), .high(7), .low(4)) bits_3754 (
        .y(_T_105),
        .in(_T_95)
    );
    wire [3:0] _T_106;
    BITS #(.width(8), .high(3), .low(0)) bits_3755 (
        .y(_T_106),
        .in(_T_95)
    );
    wire _T_108;
    wire [3:0] _WTEMP_512;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_3756 (
        .y(_WTEMP_512),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_3757 (
        .y(_T_108),
        .a(_T_105),
        .b(_WTEMP_512)
    );
    wire _T_109;
    BITS #(.width(4), .high(3), .low(3)) bits_3758 (
        .y(_T_109),
        .in(_T_105)
    );
    wire _T_111;
    BITS #(.width(4), .high(2), .low(2)) bits_3759 (
        .y(_T_111),
        .in(_T_105)
    );
    wire _T_113;
    BITS #(.width(4), .high(1), .low(1)) bits_3760 (
        .y(_T_113),
        .in(_T_105)
    );
    wire [1:0] _T_114;
    wire [1:0] _WTEMP_513;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_3761 (
        .y(_WTEMP_513),
        .in(_T_113)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_3762 (
        .y(_T_114),
        .sel(_T_111),
        .a(2'h2),
        .b(_WTEMP_513)
    );
    wire [1:0] _T_115;
    MUX_UNSIGNED #(.width(2)) u_mux_3763 (
        .y(_T_115),
        .sel(_T_109),
        .a(2'h3),
        .b(_T_114)
    );
    wire _T_116;
    BITS #(.width(4), .high(3), .low(3)) bits_3764 (
        .y(_T_116),
        .in(_T_106)
    );
    wire _T_118;
    BITS #(.width(4), .high(2), .low(2)) bits_3765 (
        .y(_T_118),
        .in(_T_106)
    );
    wire _T_120;
    BITS #(.width(4), .high(1), .low(1)) bits_3766 (
        .y(_T_120),
        .in(_T_106)
    );
    wire [1:0] _T_121;
    wire [1:0] _WTEMP_514;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_3767 (
        .y(_WTEMP_514),
        .in(_T_120)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_3768 (
        .y(_T_121),
        .sel(_T_118),
        .a(2'h2),
        .b(_WTEMP_514)
    );
    wire [1:0] _T_122;
    MUX_UNSIGNED #(.width(2)) u_mux_3769 (
        .y(_T_122),
        .sel(_T_116),
        .a(2'h3),
        .b(_T_121)
    );
    wire [1:0] _T_123;
    MUX_UNSIGNED #(.width(2)) u_mux_3770 (
        .y(_T_123),
        .sel(_T_108),
        .a(_T_115),
        .b(_T_122)
    );
    wire [2:0] _T_124;
    CAT #(.width_a(1), .width_b(2)) cat_3771 (
        .y(_T_124),
        .a(_T_108),
        .b(_T_123)
    );
    wire [2:0] _T_125;
    wire [2:0] _WTEMP_515;
    PAD_UNSIGNED #(.width(2), .n(3)) u_pad_3772 (
        .y(_WTEMP_515),
        .in(_T_104)
    );
    MUX_UNSIGNED #(.width(3)) u_mux_3773 (
        .y(_T_125),
        .sel(_T_97),
        .a(_WTEMP_515),
        .b(_T_124)
    );
    wire [3:0] _T_126;
    CAT #(.width_a(1), .width_b(3)) cat_3774 (
        .y(_T_126),
        .a(_T_97),
        .b(_T_125)
    );
    wire [15:0] _T_127;
    BITS #(.width(32), .high(31), .low(16)) bits_3775 (
        .y(_T_127),
        .in(_T_91)
    );
    wire [15:0] _T_128;
    BITS #(.width(32), .high(15), .low(0)) bits_3776 (
        .y(_T_128),
        .in(_T_91)
    );
    wire _T_130;
    wire [15:0] _WTEMP_516;
    PAD_UNSIGNED #(.width(1), .n(16)) u_pad_3777 (
        .y(_WTEMP_516),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(16)) u_neq_3778 (
        .y(_T_130),
        .a(_T_127),
        .b(_WTEMP_516)
    );
    wire [7:0] _T_131;
    BITS #(.width(16), .high(15), .low(8)) bits_3779 (
        .y(_T_131),
        .in(_T_127)
    );
    wire [7:0] _T_132;
    BITS #(.width(16), .high(7), .low(0)) bits_3780 (
        .y(_T_132),
        .in(_T_127)
    );
    wire _T_134;
    wire [7:0] _WTEMP_517;
    PAD_UNSIGNED #(.width(1), .n(8)) u_pad_3781 (
        .y(_WTEMP_517),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(8)) u_neq_3782 (
        .y(_T_134),
        .a(_T_131),
        .b(_WTEMP_517)
    );
    wire [3:0] _T_135;
    BITS #(.width(8), .high(7), .low(4)) bits_3783 (
        .y(_T_135),
        .in(_T_131)
    );
    wire [3:0] _T_136;
    BITS #(.width(8), .high(3), .low(0)) bits_3784 (
        .y(_T_136),
        .in(_T_131)
    );
    wire _T_138;
    wire [3:0] _WTEMP_518;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_3785 (
        .y(_WTEMP_518),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_3786 (
        .y(_T_138),
        .a(_T_135),
        .b(_WTEMP_518)
    );
    wire _T_139;
    BITS #(.width(4), .high(3), .low(3)) bits_3787 (
        .y(_T_139),
        .in(_T_135)
    );
    wire _T_141;
    BITS #(.width(4), .high(2), .low(2)) bits_3788 (
        .y(_T_141),
        .in(_T_135)
    );
    wire _T_143;
    BITS #(.width(4), .high(1), .low(1)) bits_3789 (
        .y(_T_143),
        .in(_T_135)
    );
    wire [1:0] _T_144;
    wire [1:0] _WTEMP_519;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_3790 (
        .y(_WTEMP_519),
        .in(_T_143)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_3791 (
        .y(_T_144),
        .sel(_T_141),
        .a(2'h2),
        .b(_WTEMP_519)
    );
    wire [1:0] _T_145;
    MUX_UNSIGNED #(.width(2)) u_mux_3792 (
        .y(_T_145),
        .sel(_T_139),
        .a(2'h3),
        .b(_T_144)
    );
    wire _T_146;
    BITS #(.width(4), .high(3), .low(3)) bits_3793 (
        .y(_T_146),
        .in(_T_136)
    );
    wire _T_148;
    BITS #(.width(4), .high(2), .low(2)) bits_3794 (
        .y(_T_148),
        .in(_T_136)
    );
    wire _T_150;
    BITS #(.width(4), .high(1), .low(1)) bits_3795 (
        .y(_T_150),
        .in(_T_136)
    );
    wire [1:0] _T_151;
    wire [1:0] _WTEMP_520;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_3796 (
        .y(_WTEMP_520),
        .in(_T_150)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_3797 (
        .y(_T_151),
        .sel(_T_148),
        .a(2'h2),
        .b(_WTEMP_520)
    );
    wire [1:0] _T_152;
    MUX_UNSIGNED #(.width(2)) u_mux_3798 (
        .y(_T_152),
        .sel(_T_146),
        .a(2'h3),
        .b(_T_151)
    );
    wire [1:0] _T_153;
    MUX_UNSIGNED #(.width(2)) u_mux_3799 (
        .y(_T_153),
        .sel(_T_138),
        .a(_T_145),
        .b(_T_152)
    );
    wire [2:0] _T_154;
    CAT #(.width_a(1), .width_b(2)) cat_3800 (
        .y(_T_154),
        .a(_T_138),
        .b(_T_153)
    );
    wire [3:0] _T_155;
    BITS #(.width(8), .high(7), .low(4)) bits_3801 (
        .y(_T_155),
        .in(_T_132)
    );
    wire [3:0] _T_156;
    BITS #(.width(8), .high(3), .low(0)) bits_3802 (
        .y(_T_156),
        .in(_T_132)
    );
    wire _T_158;
    wire [3:0] _WTEMP_521;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_3803 (
        .y(_WTEMP_521),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_3804 (
        .y(_T_158),
        .a(_T_155),
        .b(_WTEMP_521)
    );
    wire _T_159;
    BITS #(.width(4), .high(3), .low(3)) bits_3805 (
        .y(_T_159),
        .in(_T_155)
    );
    wire _T_161;
    BITS #(.width(4), .high(2), .low(2)) bits_3806 (
        .y(_T_161),
        .in(_T_155)
    );
    wire _T_163;
    BITS #(.width(4), .high(1), .low(1)) bits_3807 (
        .y(_T_163),
        .in(_T_155)
    );
    wire [1:0] _T_164;
    wire [1:0] _WTEMP_522;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_3808 (
        .y(_WTEMP_522),
        .in(_T_163)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_3809 (
        .y(_T_164),
        .sel(_T_161),
        .a(2'h2),
        .b(_WTEMP_522)
    );
    wire [1:0] _T_165;
    MUX_UNSIGNED #(.width(2)) u_mux_3810 (
        .y(_T_165),
        .sel(_T_159),
        .a(2'h3),
        .b(_T_164)
    );
    wire _T_166;
    BITS #(.width(4), .high(3), .low(3)) bits_3811 (
        .y(_T_166),
        .in(_T_156)
    );
    wire _T_168;
    BITS #(.width(4), .high(2), .low(2)) bits_3812 (
        .y(_T_168),
        .in(_T_156)
    );
    wire _T_170;
    BITS #(.width(4), .high(1), .low(1)) bits_3813 (
        .y(_T_170),
        .in(_T_156)
    );
    wire [1:0] _T_171;
    wire [1:0] _WTEMP_523;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_3814 (
        .y(_WTEMP_523),
        .in(_T_170)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_3815 (
        .y(_T_171),
        .sel(_T_168),
        .a(2'h2),
        .b(_WTEMP_523)
    );
    wire [1:0] _T_172;
    MUX_UNSIGNED #(.width(2)) u_mux_3816 (
        .y(_T_172),
        .sel(_T_166),
        .a(2'h3),
        .b(_T_171)
    );
    wire [1:0] _T_173;
    MUX_UNSIGNED #(.width(2)) u_mux_3817 (
        .y(_T_173),
        .sel(_T_158),
        .a(_T_165),
        .b(_T_172)
    );
    wire [2:0] _T_174;
    CAT #(.width_a(1), .width_b(2)) cat_3818 (
        .y(_T_174),
        .a(_T_158),
        .b(_T_173)
    );
    wire [2:0] _T_175;
    MUX_UNSIGNED #(.width(3)) u_mux_3819 (
        .y(_T_175),
        .sel(_T_134),
        .a(_T_154),
        .b(_T_174)
    );
    wire [3:0] _T_176;
    CAT #(.width_a(1), .width_b(3)) cat_3820 (
        .y(_T_176),
        .a(_T_134),
        .b(_T_175)
    );
    wire [7:0] _T_177;
    BITS #(.width(16), .high(15), .low(8)) bits_3821 (
        .y(_T_177),
        .in(_T_128)
    );
    wire [7:0] _T_178;
    BITS #(.width(16), .high(7), .low(0)) bits_3822 (
        .y(_T_178),
        .in(_T_128)
    );
    wire _T_180;
    wire [7:0] _WTEMP_524;
    PAD_UNSIGNED #(.width(1), .n(8)) u_pad_3823 (
        .y(_WTEMP_524),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(8)) u_neq_3824 (
        .y(_T_180),
        .a(_T_177),
        .b(_WTEMP_524)
    );
    wire [3:0] _T_181;
    BITS #(.width(8), .high(7), .low(4)) bits_3825 (
        .y(_T_181),
        .in(_T_177)
    );
    wire [3:0] _T_182;
    BITS #(.width(8), .high(3), .low(0)) bits_3826 (
        .y(_T_182),
        .in(_T_177)
    );
    wire _T_184;
    wire [3:0] _WTEMP_525;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_3827 (
        .y(_WTEMP_525),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_3828 (
        .y(_T_184),
        .a(_T_181),
        .b(_WTEMP_525)
    );
    wire _T_185;
    BITS #(.width(4), .high(3), .low(3)) bits_3829 (
        .y(_T_185),
        .in(_T_181)
    );
    wire _T_187;
    BITS #(.width(4), .high(2), .low(2)) bits_3830 (
        .y(_T_187),
        .in(_T_181)
    );
    wire _T_189;
    BITS #(.width(4), .high(1), .low(1)) bits_3831 (
        .y(_T_189),
        .in(_T_181)
    );
    wire [1:0] _T_190;
    wire [1:0] _WTEMP_526;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_3832 (
        .y(_WTEMP_526),
        .in(_T_189)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_3833 (
        .y(_T_190),
        .sel(_T_187),
        .a(2'h2),
        .b(_WTEMP_526)
    );
    wire [1:0] _T_191;
    MUX_UNSIGNED #(.width(2)) u_mux_3834 (
        .y(_T_191),
        .sel(_T_185),
        .a(2'h3),
        .b(_T_190)
    );
    wire _T_192;
    BITS #(.width(4), .high(3), .low(3)) bits_3835 (
        .y(_T_192),
        .in(_T_182)
    );
    wire _T_194;
    BITS #(.width(4), .high(2), .low(2)) bits_3836 (
        .y(_T_194),
        .in(_T_182)
    );
    wire _T_196;
    BITS #(.width(4), .high(1), .low(1)) bits_3837 (
        .y(_T_196),
        .in(_T_182)
    );
    wire [1:0] _T_197;
    wire [1:0] _WTEMP_527;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_3838 (
        .y(_WTEMP_527),
        .in(_T_196)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_3839 (
        .y(_T_197),
        .sel(_T_194),
        .a(2'h2),
        .b(_WTEMP_527)
    );
    wire [1:0] _T_198;
    MUX_UNSIGNED #(.width(2)) u_mux_3840 (
        .y(_T_198),
        .sel(_T_192),
        .a(2'h3),
        .b(_T_197)
    );
    wire [1:0] _T_199;
    MUX_UNSIGNED #(.width(2)) u_mux_3841 (
        .y(_T_199),
        .sel(_T_184),
        .a(_T_191),
        .b(_T_198)
    );
    wire [2:0] _T_200;
    CAT #(.width_a(1), .width_b(2)) cat_3842 (
        .y(_T_200),
        .a(_T_184),
        .b(_T_199)
    );
    wire [3:0] _T_201;
    BITS #(.width(8), .high(7), .low(4)) bits_3843 (
        .y(_T_201),
        .in(_T_178)
    );
    wire [3:0] _T_202;
    BITS #(.width(8), .high(3), .low(0)) bits_3844 (
        .y(_T_202),
        .in(_T_178)
    );
    wire _T_204;
    wire [3:0] _WTEMP_528;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_3845 (
        .y(_WTEMP_528),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_3846 (
        .y(_T_204),
        .a(_T_201),
        .b(_WTEMP_528)
    );
    wire _T_205;
    BITS #(.width(4), .high(3), .low(3)) bits_3847 (
        .y(_T_205),
        .in(_T_201)
    );
    wire _T_207;
    BITS #(.width(4), .high(2), .low(2)) bits_3848 (
        .y(_T_207),
        .in(_T_201)
    );
    wire _T_209;
    BITS #(.width(4), .high(1), .low(1)) bits_3849 (
        .y(_T_209),
        .in(_T_201)
    );
    wire [1:0] _T_210;
    wire [1:0] _WTEMP_529;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_3850 (
        .y(_WTEMP_529),
        .in(_T_209)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_3851 (
        .y(_T_210),
        .sel(_T_207),
        .a(2'h2),
        .b(_WTEMP_529)
    );
    wire [1:0] _T_211;
    MUX_UNSIGNED #(.width(2)) u_mux_3852 (
        .y(_T_211),
        .sel(_T_205),
        .a(2'h3),
        .b(_T_210)
    );
    wire _T_212;
    BITS #(.width(4), .high(3), .low(3)) bits_3853 (
        .y(_T_212),
        .in(_T_202)
    );
    wire _T_214;
    BITS #(.width(4), .high(2), .low(2)) bits_3854 (
        .y(_T_214),
        .in(_T_202)
    );
    wire _T_216;
    BITS #(.width(4), .high(1), .low(1)) bits_3855 (
        .y(_T_216),
        .in(_T_202)
    );
    wire [1:0] _T_217;
    wire [1:0] _WTEMP_530;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_3856 (
        .y(_WTEMP_530),
        .in(_T_216)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_3857 (
        .y(_T_217),
        .sel(_T_214),
        .a(2'h2),
        .b(_WTEMP_530)
    );
    wire [1:0] _T_218;
    MUX_UNSIGNED #(.width(2)) u_mux_3858 (
        .y(_T_218),
        .sel(_T_212),
        .a(2'h3),
        .b(_T_217)
    );
    wire [1:0] _T_219;
    MUX_UNSIGNED #(.width(2)) u_mux_3859 (
        .y(_T_219),
        .sel(_T_204),
        .a(_T_211),
        .b(_T_218)
    );
    wire [2:0] _T_220;
    CAT #(.width_a(1), .width_b(2)) cat_3860 (
        .y(_T_220),
        .a(_T_204),
        .b(_T_219)
    );
    wire [2:0] _T_221;
    MUX_UNSIGNED #(.width(3)) u_mux_3861 (
        .y(_T_221),
        .sel(_T_180),
        .a(_T_200),
        .b(_T_220)
    );
    wire [3:0] _T_222;
    CAT #(.width_a(1), .width_b(3)) cat_3862 (
        .y(_T_222),
        .a(_T_180),
        .b(_T_221)
    );
    wire [3:0] _T_223;
    MUX_UNSIGNED #(.width(4)) u_mux_3863 (
        .y(_T_223),
        .sel(_T_130),
        .a(_T_176),
        .b(_T_222)
    );
    wire [4:0] _T_224;
    CAT #(.width_a(1), .width_b(4)) cat_3864 (
        .y(_T_224),
        .a(_T_130),
        .b(_T_223)
    );
    wire [4:0] _T_225;
    wire [4:0] _WTEMP_531;
    PAD_UNSIGNED #(.width(4), .n(5)) u_pad_3865 (
        .y(_WTEMP_531),
        .in(_T_126)
    );
    MUX_UNSIGNED #(.width(5)) u_mux_3866 (
        .y(_T_225),
        .sel(_T_93),
        .a(_WTEMP_531),
        .b(_T_224)
    );
    wire [5:0] _T_226;
    CAT #(.width_a(1), .width_b(5)) cat_3867 (
        .y(_T_226),
        .a(_T_93),
        .b(_T_225)
    );
    wire [31:0] _T_227;
    BITS #(.width(64), .high(63), .low(32)) bits_3868 (
        .y(_T_227),
        .in(_T_87)
    );
    wire [31:0] _T_228;
    BITS #(.width(64), .high(31), .low(0)) bits_3869 (
        .y(_T_228),
        .in(_T_87)
    );
    wire _T_230;
    wire [31:0] _WTEMP_532;
    PAD_UNSIGNED #(.width(1), .n(32)) u_pad_3870 (
        .y(_WTEMP_532),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(32)) u_neq_3871 (
        .y(_T_230),
        .a(_T_227),
        .b(_WTEMP_532)
    );
    wire [15:0] _T_231;
    BITS #(.width(32), .high(31), .low(16)) bits_3872 (
        .y(_T_231),
        .in(_T_227)
    );
    wire [15:0] _T_232;
    BITS #(.width(32), .high(15), .low(0)) bits_3873 (
        .y(_T_232),
        .in(_T_227)
    );
    wire _T_234;
    wire [15:0] _WTEMP_533;
    PAD_UNSIGNED #(.width(1), .n(16)) u_pad_3874 (
        .y(_WTEMP_533),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(16)) u_neq_3875 (
        .y(_T_234),
        .a(_T_231),
        .b(_WTEMP_533)
    );
    wire [7:0] _T_235;
    BITS #(.width(16), .high(15), .low(8)) bits_3876 (
        .y(_T_235),
        .in(_T_231)
    );
    wire [7:0] _T_236;
    BITS #(.width(16), .high(7), .low(0)) bits_3877 (
        .y(_T_236),
        .in(_T_231)
    );
    wire _T_238;
    wire [7:0] _WTEMP_534;
    PAD_UNSIGNED #(.width(1), .n(8)) u_pad_3878 (
        .y(_WTEMP_534),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(8)) u_neq_3879 (
        .y(_T_238),
        .a(_T_235),
        .b(_WTEMP_534)
    );
    wire [3:0] _T_239;
    BITS #(.width(8), .high(7), .low(4)) bits_3880 (
        .y(_T_239),
        .in(_T_235)
    );
    wire [3:0] _T_240;
    BITS #(.width(8), .high(3), .low(0)) bits_3881 (
        .y(_T_240),
        .in(_T_235)
    );
    wire _T_242;
    wire [3:0] _WTEMP_535;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_3882 (
        .y(_WTEMP_535),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_3883 (
        .y(_T_242),
        .a(_T_239),
        .b(_WTEMP_535)
    );
    wire _T_243;
    BITS #(.width(4), .high(3), .low(3)) bits_3884 (
        .y(_T_243),
        .in(_T_239)
    );
    wire _T_245;
    BITS #(.width(4), .high(2), .low(2)) bits_3885 (
        .y(_T_245),
        .in(_T_239)
    );
    wire _T_247;
    BITS #(.width(4), .high(1), .low(1)) bits_3886 (
        .y(_T_247),
        .in(_T_239)
    );
    wire [1:0] _T_248;
    wire [1:0] _WTEMP_536;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_3887 (
        .y(_WTEMP_536),
        .in(_T_247)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_3888 (
        .y(_T_248),
        .sel(_T_245),
        .a(2'h2),
        .b(_WTEMP_536)
    );
    wire [1:0] _T_249;
    MUX_UNSIGNED #(.width(2)) u_mux_3889 (
        .y(_T_249),
        .sel(_T_243),
        .a(2'h3),
        .b(_T_248)
    );
    wire _T_250;
    BITS #(.width(4), .high(3), .low(3)) bits_3890 (
        .y(_T_250),
        .in(_T_240)
    );
    wire _T_252;
    BITS #(.width(4), .high(2), .low(2)) bits_3891 (
        .y(_T_252),
        .in(_T_240)
    );
    wire _T_254;
    BITS #(.width(4), .high(1), .low(1)) bits_3892 (
        .y(_T_254),
        .in(_T_240)
    );
    wire [1:0] _T_255;
    wire [1:0] _WTEMP_537;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_3893 (
        .y(_WTEMP_537),
        .in(_T_254)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_3894 (
        .y(_T_255),
        .sel(_T_252),
        .a(2'h2),
        .b(_WTEMP_537)
    );
    wire [1:0] _T_256;
    MUX_UNSIGNED #(.width(2)) u_mux_3895 (
        .y(_T_256),
        .sel(_T_250),
        .a(2'h3),
        .b(_T_255)
    );
    wire [1:0] _T_257;
    MUX_UNSIGNED #(.width(2)) u_mux_3896 (
        .y(_T_257),
        .sel(_T_242),
        .a(_T_249),
        .b(_T_256)
    );
    wire [2:0] _T_258;
    CAT #(.width_a(1), .width_b(2)) cat_3897 (
        .y(_T_258),
        .a(_T_242),
        .b(_T_257)
    );
    wire [3:0] _T_259;
    BITS #(.width(8), .high(7), .low(4)) bits_3898 (
        .y(_T_259),
        .in(_T_236)
    );
    wire [3:0] _T_260;
    BITS #(.width(8), .high(3), .low(0)) bits_3899 (
        .y(_T_260),
        .in(_T_236)
    );
    wire _T_262;
    wire [3:0] _WTEMP_538;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_3900 (
        .y(_WTEMP_538),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_3901 (
        .y(_T_262),
        .a(_T_259),
        .b(_WTEMP_538)
    );
    wire _T_263;
    BITS #(.width(4), .high(3), .low(3)) bits_3902 (
        .y(_T_263),
        .in(_T_259)
    );
    wire _T_265;
    BITS #(.width(4), .high(2), .low(2)) bits_3903 (
        .y(_T_265),
        .in(_T_259)
    );
    wire _T_267;
    BITS #(.width(4), .high(1), .low(1)) bits_3904 (
        .y(_T_267),
        .in(_T_259)
    );
    wire [1:0] _T_268;
    wire [1:0] _WTEMP_539;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_3905 (
        .y(_WTEMP_539),
        .in(_T_267)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_3906 (
        .y(_T_268),
        .sel(_T_265),
        .a(2'h2),
        .b(_WTEMP_539)
    );
    wire [1:0] _T_269;
    MUX_UNSIGNED #(.width(2)) u_mux_3907 (
        .y(_T_269),
        .sel(_T_263),
        .a(2'h3),
        .b(_T_268)
    );
    wire _T_270;
    BITS #(.width(4), .high(3), .low(3)) bits_3908 (
        .y(_T_270),
        .in(_T_260)
    );
    wire _T_272;
    BITS #(.width(4), .high(2), .low(2)) bits_3909 (
        .y(_T_272),
        .in(_T_260)
    );
    wire _T_274;
    BITS #(.width(4), .high(1), .low(1)) bits_3910 (
        .y(_T_274),
        .in(_T_260)
    );
    wire [1:0] _T_275;
    wire [1:0] _WTEMP_540;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_3911 (
        .y(_WTEMP_540),
        .in(_T_274)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_3912 (
        .y(_T_275),
        .sel(_T_272),
        .a(2'h2),
        .b(_WTEMP_540)
    );
    wire [1:0] _T_276;
    MUX_UNSIGNED #(.width(2)) u_mux_3913 (
        .y(_T_276),
        .sel(_T_270),
        .a(2'h3),
        .b(_T_275)
    );
    wire [1:0] _T_277;
    MUX_UNSIGNED #(.width(2)) u_mux_3914 (
        .y(_T_277),
        .sel(_T_262),
        .a(_T_269),
        .b(_T_276)
    );
    wire [2:0] _T_278;
    CAT #(.width_a(1), .width_b(2)) cat_3915 (
        .y(_T_278),
        .a(_T_262),
        .b(_T_277)
    );
    wire [2:0] _T_279;
    MUX_UNSIGNED #(.width(3)) u_mux_3916 (
        .y(_T_279),
        .sel(_T_238),
        .a(_T_258),
        .b(_T_278)
    );
    wire [3:0] _T_280;
    CAT #(.width_a(1), .width_b(3)) cat_3917 (
        .y(_T_280),
        .a(_T_238),
        .b(_T_279)
    );
    wire [7:0] _T_281;
    BITS #(.width(16), .high(15), .low(8)) bits_3918 (
        .y(_T_281),
        .in(_T_232)
    );
    wire [7:0] _T_282;
    BITS #(.width(16), .high(7), .low(0)) bits_3919 (
        .y(_T_282),
        .in(_T_232)
    );
    wire _T_284;
    wire [7:0] _WTEMP_541;
    PAD_UNSIGNED #(.width(1), .n(8)) u_pad_3920 (
        .y(_WTEMP_541),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(8)) u_neq_3921 (
        .y(_T_284),
        .a(_T_281),
        .b(_WTEMP_541)
    );
    wire [3:0] _T_285;
    BITS #(.width(8), .high(7), .low(4)) bits_3922 (
        .y(_T_285),
        .in(_T_281)
    );
    wire [3:0] _T_286;
    BITS #(.width(8), .high(3), .low(0)) bits_3923 (
        .y(_T_286),
        .in(_T_281)
    );
    wire _T_288;
    wire [3:0] _WTEMP_542;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_3924 (
        .y(_WTEMP_542),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_3925 (
        .y(_T_288),
        .a(_T_285),
        .b(_WTEMP_542)
    );
    wire _T_289;
    BITS #(.width(4), .high(3), .low(3)) bits_3926 (
        .y(_T_289),
        .in(_T_285)
    );
    wire _T_291;
    BITS #(.width(4), .high(2), .low(2)) bits_3927 (
        .y(_T_291),
        .in(_T_285)
    );
    wire _T_293;
    BITS #(.width(4), .high(1), .low(1)) bits_3928 (
        .y(_T_293),
        .in(_T_285)
    );
    wire [1:0] _T_294;
    wire [1:0] _WTEMP_543;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_3929 (
        .y(_WTEMP_543),
        .in(_T_293)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_3930 (
        .y(_T_294),
        .sel(_T_291),
        .a(2'h2),
        .b(_WTEMP_543)
    );
    wire [1:0] _T_295;
    MUX_UNSIGNED #(.width(2)) u_mux_3931 (
        .y(_T_295),
        .sel(_T_289),
        .a(2'h3),
        .b(_T_294)
    );
    wire _T_296;
    BITS #(.width(4), .high(3), .low(3)) bits_3932 (
        .y(_T_296),
        .in(_T_286)
    );
    wire _T_298;
    BITS #(.width(4), .high(2), .low(2)) bits_3933 (
        .y(_T_298),
        .in(_T_286)
    );
    wire _T_300;
    BITS #(.width(4), .high(1), .low(1)) bits_3934 (
        .y(_T_300),
        .in(_T_286)
    );
    wire [1:0] _T_301;
    wire [1:0] _WTEMP_544;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_3935 (
        .y(_WTEMP_544),
        .in(_T_300)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_3936 (
        .y(_T_301),
        .sel(_T_298),
        .a(2'h2),
        .b(_WTEMP_544)
    );
    wire [1:0] _T_302;
    MUX_UNSIGNED #(.width(2)) u_mux_3937 (
        .y(_T_302),
        .sel(_T_296),
        .a(2'h3),
        .b(_T_301)
    );
    wire [1:0] _T_303;
    MUX_UNSIGNED #(.width(2)) u_mux_3938 (
        .y(_T_303),
        .sel(_T_288),
        .a(_T_295),
        .b(_T_302)
    );
    wire [2:0] _T_304;
    CAT #(.width_a(1), .width_b(2)) cat_3939 (
        .y(_T_304),
        .a(_T_288),
        .b(_T_303)
    );
    wire [3:0] _T_305;
    BITS #(.width(8), .high(7), .low(4)) bits_3940 (
        .y(_T_305),
        .in(_T_282)
    );
    wire [3:0] _T_306;
    BITS #(.width(8), .high(3), .low(0)) bits_3941 (
        .y(_T_306),
        .in(_T_282)
    );
    wire _T_308;
    wire [3:0] _WTEMP_545;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_3942 (
        .y(_WTEMP_545),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_3943 (
        .y(_T_308),
        .a(_T_305),
        .b(_WTEMP_545)
    );
    wire _T_309;
    BITS #(.width(4), .high(3), .low(3)) bits_3944 (
        .y(_T_309),
        .in(_T_305)
    );
    wire _T_311;
    BITS #(.width(4), .high(2), .low(2)) bits_3945 (
        .y(_T_311),
        .in(_T_305)
    );
    wire _T_313;
    BITS #(.width(4), .high(1), .low(1)) bits_3946 (
        .y(_T_313),
        .in(_T_305)
    );
    wire [1:0] _T_314;
    wire [1:0] _WTEMP_546;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_3947 (
        .y(_WTEMP_546),
        .in(_T_313)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_3948 (
        .y(_T_314),
        .sel(_T_311),
        .a(2'h2),
        .b(_WTEMP_546)
    );
    wire [1:0] _T_315;
    MUX_UNSIGNED #(.width(2)) u_mux_3949 (
        .y(_T_315),
        .sel(_T_309),
        .a(2'h3),
        .b(_T_314)
    );
    wire _T_316;
    BITS #(.width(4), .high(3), .low(3)) bits_3950 (
        .y(_T_316),
        .in(_T_306)
    );
    wire _T_318;
    BITS #(.width(4), .high(2), .low(2)) bits_3951 (
        .y(_T_318),
        .in(_T_306)
    );
    wire _T_320;
    BITS #(.width(4), .high(1), .low(1)) bits_3952 (
        .y(_T_320),
        .in(_T_306)
    );
    wire [1:0] _T_321;
    wire [1:0] _WTEMP_547;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_3953 (
        .y(_WTEMP_547),
        .in(_T_320)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_3954 (
        .y(_T_321),
        .sel(_T_318),
        .a(2'h2),
        .b(_WTEMP_547)
    );
    wire [1:0] _T_322;
    MUX_UNSIGNED #(.width(2)) u_mux_3955 (
        .y(_T_322),
        .sel(_T_316),
        .a(2'h3),
        .b(_T_321)
    );
    wire [1:0] _T_323;
    MUX_UNSIGNED #(.width(2)) u_mux_3956 (
        .y(_T_323),
        .sel(_T_308),
        .a(_T_315),
        .b(_T_322)
    );
    wire [2:0] _T_324;
    CAT #(.width_a(1), .width_b(2)) cat_3957 (
        .y(_T_324),
        .a(_T_308),
        .b(_T_323)
    );
    wire [2:0] _T_325;
    MUX_UNSIGNED #(.width(3)) u_mux_3958 (
        .y(_T_325),
        .sel(_T_284),
        .a(_T_304),
        .b(_T_324)
    );
    wire [3:0] _T_326;
    CAT #(.width_a(1), .width_b(3)) cat_3959 (
        .y(_T_326),
        .a(_T_284),
        .b(_T_325)
    );
    wire [3:0] _T_327;
    MUX_UNSIGNED #(.width(4)) u_mux_3960 (
        .y(_T_327),
        .sel(_T_234),
        .a(_T_280),
        .b(_T_326)
    );
    wire [4:0] _T_328;
    CAT #(.width_a(1), .width_b(4)) cat_3961 (
        .y(_T_328),
        .a(_T_234),
        .b(_T_327)
    );
    wire [15:0] _T_329;
    BITS #(.width(32), .high(31), .low(16)) bits_3962 (
        .y(_T_329),
        .in(_T_228)
    );
    wire [15:0] _T_330;
    BITS #(.width(32), .high(15), .low(0)) bits_3963 (
        .y(_T_330),
        .in(_T_228)
    );
    wire _T_332;
    wire [15:0] _WTEMP_548;
    PAD_UNSIGNED #(.width(1), .n(16)) u_pad_3964 (
        .y(_WTEMP_548),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(16)) u_neq_3965 (
        .y(_T_332),
        .a(_T_329),
        .b(_WTEMP_548)
    );
    wire [7:0] _T_333;
    BITS #(.width(16), .high(15), .low(8)) bits_3966 (
        .y(_T_333),
        .in(_T_329)
    );
    wire [7:0] _T_334;
    BITS #(.width(16), .high(7), .low(0)) bits_3967 (
        .y(_T_334),
        .in(_T_329)
    );
    wire _T_336;
    wire [7:0] _WTEMP_549;
    PAD_UNSIGNED #(.width(1), .n(8)) u_pad_3968 (
        .y(_WTEMP_549),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(8)) u_neq_3969 (
        .y(_T_336),
        .a(_T_333),
        .b(_WTEMP_549)
    );
    wire [3:0] _T_337;
    BITS #(.width(8), .high(7), .low(4)) bits_3970 (
        .y(_T_337),
        .in(_T_333)
    );
    wire [3:0] _T_338;
    BITS #(.width(8), .high(3), .low(0)) bits_3971 (
        .y(_T_338),
        .in(_T_333)
    );
    wire _T_340;
    wire [3:0] _WTEMP_550;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_3972 (
        .y(_WTEMP_550),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_3973 (
        .y(_T_340),
        .a(_T_337),
        .b(_WTEMP_550)
    );
    wire _T_341;
    BITS #(.width(4), .high(3), .low(3)) bits_3974 (
        .y(_T_341),
        .in(_T_337)
    );
    wire _T_343;
    BITS #(.width(4), .high(2), .low(2)) bits_3975 (
        .y(_T_343),
        .in(_T_337)
    );
    wire _T_345;
    BITS #(.width(4), .high(1), .low(1)) bits_3976 (
        .y(_T_345),
        .in(_T_337)
    );
    wire [1:0] _T_346;
    wire [1:0] _WTEMP_551;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_3977 (
        .y(_WTEMP_551),
        .in(_T_345)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_3978 (
        .y(_T_346),
        .sel(_T_343),
        .a(2'h2),
        .b(_WTEMP_551)
    );
    wire [1:0] _T_347;
    MUX_UNSIGNED #(.width(2)) u_mux_3979 (
        .y(_T_347),
        .sel(_T_341),
        .a(2'h3),
        .b(_T_346)
    );
    wire _T_348;
    BITS #(.width(4), .high(3), .low(3)) bits_3980 (
        .y(_T_348),
        .in(_T_338)
    );
    wire _T_350;
    BITS #(.width(4), .high(2), .low(2)) bits_3981 (
        .y(_T_350),
        .in(_T_338)
    );
    wire _T_352;
    BITS #(.width(4), .high(1), .low(1)) bits_3982 (
        .y(_T_352),
        .in(_T_338)
    );
    wire [1:0] _T_353;
    wire [1:0] _WTEMP_552;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_3983 (
        .y(_WTEMP_552),
        .in(_T_352)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_3984 (
        .y(_T_353),
        .sel(_T_350),
        .a(2'h2),
        .b(_WTEMP_552)
    );
    wire [1:0] _T_354;
    MUX_UNSIGNED #(.width(2)) u_mux_3985 (
        .y(_T_354),
        .sel(_T_348),
        .a(2'h3),
        .b(_T_353)
    );
    wire [1:0] _T_355;
    MUX_UNSIGNED #(.width(2)) u_mux_3986 (
        .y(_T_355),
        .sel(_T_340),
        .a(_T_347),
        .b(_T_354)
    );
    wire [2:0] _T_356;
    CAT #(.width_a(1), .width_b(2)) cat_3987 (
        .y(_T_356),
        .a(_T_340),
        .b(_T_355)
    );
    wire [3:0] _T_357;
    BITS #(.width(8), .high(7), .low(4)) bits_3988 (
        .y(_T_357),
        .in(_T_334)
    );
    wire [3:0] _T_358;
    BITS #(.width(8), .high(3), .low(0)) bits_3989 (
        .y(_T_358),
        .in(_T_334)
    );
    wire _T_360;
    wire [3:0] _WTEMP_553;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_3990 (
        .y(_WTEMP_553),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_3991 (
        .y(_T_360),
        .a(_T_357),
        .b(_WTEMP_553)
    );
    wire _T_361;
    BITS #(.width(4), .high(3), .low(3)) bits_3992 (
        .y(_T_361),
        .in(_T_357)
    );
    wire _T_363;
    BITS #(.width(4), .high(2), .low(2)) bits_3993 (
        .y(_T_363),
        .in(_T_357)
    );
    wire _T_365;
    BITS #(.width(4), .high(1), .low(1)) bits_3994 (
        .y(_T_365),
        .in(_T_357)
    );
    wire [1:0] _T_366;
    wire [1:0] _WTEMP_554;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_3995 (
        .y(_WTEMP_554),
        .in(_T_365)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_3996 (
        .y(_T_366),
        .sel(_T_363),
        .a(2'h2),
        .b(_WTEMP_554)
    );
    wire [1:0] _T_367;
    MUX_UNSIGNED #(.width(2)) u_mux_3997 (
        .y(_T_367),
        .sel(_T_361),
        .a(2'h3),
        .b(_T_366)
    );
    wire _T_368;
    BITS #(.width(4), .high(3), .low(3)) bits_3998 (
        .y(_T_368),
        .in(_T_358)
    );
    wire _T_370;
    BITS #(.width(4), .high(2), .low(2)) bits_3999 (
        .y(_T_370),
        .in(_T_358)
    );
    wire _T_372;
    BITS #(.width(4), .high(1), .low(1)) bits_4000 (
        .y(_T_372),
        .in(_T_358)
    );
    wire [1:0] _T_373;
    wire [1:0] _WTEMP_555;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_4001 (
        .y(_WTEMP_555),
        .in(_T_372)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_4002 (
        .y(_T_373),
        .sel(_T_370),
        .a(2'h2),
        .b(_WTEMP_555)
    );
    wire [1:0] _T_374;
    MUX_UNSIGNED #(.width(2)) u_mux_4003 (
        .y(_T_374),
        .sel(_T_368),
        .a(2'h3),
        .b(_T_373)
    );
    wire [1:0] _T_375;
    MUX_UNSIGNED #(.width(2)) u_mux_4004 (
        .y(_T_375),
        .sel(_T_360),
        .a(_T_367),
        .b(_T_374)
    );
    wire [2:0] _T_376;
    CAT #(.width_a(1), .width_b(2)) cat_4005 (
        .y(_T_376),
        .a(_T_360),
        .b(_T_375)
    );
    wire [2:0] _T_377;
    MUX_UNSIGNED #(.width(3)) u_mux_4006 (
        .y(_T_377),
        .sel(_T_336),
        .a(_T_356),
        .b(_T_376)
    );
    wire [3:0] _T_378;
    CAT #(.width_a(1), .width_b(3)) cat_4007 (
        .y(_T_378),
        .a(_T_336),
        .b(_T_377)
    );
    wire [7:0] _T_379;
    BITS #(.width(16), .high(15), .low(8)) bits_4008 (
        .y(_T_379),
        .in(_T_330)
    );
    wire [7:0] _T_380;
    BITS #(.width(16), .high(7), .low(0)) bits_4009 (
        .y(_T_380),
        .in(_T_330)
    );
    wire _T_382;
    wire [7:0] _WTEMP_556;
    PAD_UNSIGNED #(.width(1), .n(8)) u_pad_4010 (
        .y(_WTEMP_556),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(8)) u_neq_4011 (
        .y(_T_382),
        .a(_T_379),
        .b(_WTEMP_556)
    );
    wire [3:0] _T_383;
    BITS #(.width(8), .high(7), .low(4)) bits_4012 (
        .y(_T_383),
        .in(_T_379)
    );
    wire [3:0] _T_384;
    BITS #(.width(8), .high(3), .low(0)) bits_4013 (
        .y(_T_384),
        .in(_T_379)
    );
    wire _T_386;
    wire [3:0] _WTEMP_557;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_4014 (
        .y(_WTEMP_557),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_4015 (
        .y(_T_386),
        .a(_T_383),
        .b(_WTEMP_557)
    );
    wire _T_387;
    BITS #(.width(4), .high(3), .low(3)) bits_4016 (
        .y(_T_387),
        .in(_T_383)
    );
    wire _T_389;
    BITS #(.width(4), .high(2), .low(2)) bits_4017 (
        .y(_T_389),
        .in(_T_383)
    );
    wire _T_391;
    BITS #(.width(4), .high(1), .low(1)) bits_4018 (
        .y(_T_391),
        .in(_T_383)
    );
    wire [1:0] _T_392;
    wire [1:0] _WTEMP_558;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_4019 (
        .y(_WTEMP_558),
        .in(_T_391)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_4020 (
        .y(_T_392),
        .sel(_T_389),
        .a(2'h2),
        .b(_WTEMP_558)
    );
    wire [1:0] _T_393;
    MUX_UNSIGNED #(.width(2)) u_mux_4021 (
        .y(_T_393),
        .sel(_T_387),
        .a(2'h3),
        .b(_T_392)
    );
    wire _T_394;
    BITS #(.width(4), .high(3), .low(3)) bits_4022 (
        .y(_T_394),
        .in(_T_384)
    );
    wire _T_396;
    BITS #(.width(4), .high(2), .low(2)) bits_4023 (
        .y(_T_396),
        .in(_T_384)
    );
    wire _T_398;
    BITS #(.width(4), .high(1), .low(1)) bits_4024 (
        .y(_T_398),
        .in(_T_384)
    );
    wire [1:0] _T_399;
    wire [1:0] _WTEMP_559;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_4025 (
        .y(_WTEMP_559),
        .in(_T_398)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_4026 (
        .y(_T_399),
        .sel(_T_396),
        .a(2'h2),
        .b(_WTEMP_559)
    );
    wire [1:0] _T_400;
    MUX_UNSIGNED #(.width(2)) u_mux_4027 (
        .y(_T_400),
        .sel(_T_394),
        .a(2'h3),
        .b(_T_399)
    );
    wire [1:0] _T_401;
    MUX_UNSIGNED #(.width(2)) u_mux_4028 (
        .y(_T_401),
        .sel(_T_386),
        .a(_T_393),
        .b(_T_400)
    );
    wire [2:0] _T_402;
    CAT #(.width_a(1), .width_b(2)) cat_4029 (
        .y(_T_402),
        .a(_T_386),
        .b(_T_401)
    );
    wire [3:0] _T_403;
    BITS #(.width(8), .high(7), .low(4)) bits_4030 (
        .y(_T_403),
        .in(_T_380)
    );
    wire [3:0] _T_404;
    BITS #(.width(8), .high(3), .low(0)) bits_4031 (
        .y(_T_404),
        .in(_T_380)
    );
    wire _T_406;
    wire [3:0] _WTEMP_560;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_4032 (
        .y(_WTEMP_560),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_4033 (
        .y(_T_406),
        .a(_T_403),
        .b(_WTEMP_560)
    );
    wire _T_407;
    BITS #(.width(4), .high(3), .low(3)) bits_4034 (
        .y(_T_407),
        .in(_T_403)
    );
    wire _T_409;
    BITS #(.width(4), .high(2), .low(2)) bits_4035 (
        .y(_T_409),
        .in(_T_403)
    );
    wire _T_411;
    BITS #(.width(4), .high(1), .low(1)) bits_4036 (
        .y(_T_411),
        .in(_T_403)
    );
    wire [1:0] _T_412;
    wire [1:0] _WTEMP_561;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_4037 (
        .y(_WTEMP_561),
        .in(_T_411)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_4038 (
        .y(_T_412),
        .sel(_T_409),
        .a(2'h2),
        .b(_WTEMP_561)
    );
    wire [1:0] _T_413;
    MUX_UNSIGNED #(.width(2)) u_mux_4039 (
        .y(_T_413),
        .sel(_T_407),
        .a(2'h3),
        .b(_T_412)
    );
    wire _T_414;
    BITS #(.width(4), .high(3), .low(3)) bits_4040 (
        .y(_T_414),
        .in(_T_404)
    );
    wire _T_416;
    BITS #(.width(4), .high(2), .low(2)) bits_4041 (
        .y(_T_416),
        .in(_T_404)
    );
    wire _T_418;
    BITS #(.width(4), .high(1), .low(1)) bits_4042 (
        .y(_T_418),
        .in(_T_404)
    );
    wire [1:0] _T_419;
    wire [1:0] _WTEMP_562;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_4043 (
        .y(_WTEMP_562),
        .in(_T_418)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_4044 (
        .y(_T_419),
        .sel(_T_416),
        .a(2'h2),
        .b(_WTEMP_562)
    );
    wire [1:0] _T_420;
    MUX_UNSIGNED #(.width(2)) u_mux_4045 (
        .y(_T_420),
        .sel(_T_414),
        .a(2'h3),
        .b(_T_419)
    );
    wire [1:0] _T_421;
    MUX_UNSIGNED #(.width(2)) u_mux_4046 (
        .y(_T_421),
        .sel(_T_406),
        .a(_T_413),
        .b(_T_420)
    );
    wire [2:0] _T_422;
    CAT #(.width_a(1), .width_b(2)) cat_4047 (
        .y(_T_422),
        .a(_T_406),
        .b(_T_421)
    );
    wire [2:0] _T_423;
    MUX_UNSIGNED #(.width(3)) u_mux_4048 (
        .y(_T_423),
        .sel(_T_382),
        .a(_T_402),
        .b(_T_422)
    );
    wire [3:0] _T_424;
    CAT #(.width_a(1), .width_b(3)) cat_4049 (
        .y(_T_424),
        .a(_T_382),
        .b(_T_423)
    );
    wire [3:0] _T_425;
    MUX_UNSIGNED #(.width(4)) u_mux_4050 (
        .y(_T_425),
        .sel(_T_332),
        .a(_T_378),
        .b(_T_424)
    );
    wire [4:0] _T_426;
    CAT #(.width_a(1), .width_b(4)) cat_4051 (
        .y(_T_426),
        .a(_T_332),
        .b(_T_425)
    );
    wire [4:0] _T_427;
    MUX_UNSIGNED #(.width(5)) u_mux_4052 (
        .y(_T_427),
        .sel(_T_230),
        .a(_T_328),
        .b(_T_426)
    );
    wire [5:0] _T_428;
    CAT #(.width_a(1), .width_b(5)) cat_4053 (
        .y(_T_428),
        .a(_T_230),
        .b(_T_427)
    );
    wire [5:0] _T_429;
    MUX_UNSIGNED #(.width(6)) u_mux_4054 (
        .y(_T_429),
        .sel(_T_89),
        .a(_T_226),
        .b(_T_428)
    );
    wire [6:0] _T_430;
    CAT #(.width_a(1), .width_b(6)) cat_4055 (
        .y(_T_430),
        .a(_T_89),
        .b(_T_429)
    );
    wire [8:0] _T_431;
    wire [7:0] _WTEMP_563;
    PAD_UNSIGNED #(.width(7), .n(8)) u_pad_4056 (
        .y(_WTEMP_563),
        .in(_T_430)
    );
    SUB_UNSIGNED #(.width(8)) u_sub_4057 (
        .y(_T_431),
        .a(8'hA0),
        .b(_WTEMP_563)
    );
    wire [8:0] _T_432;
    ASUINT #(.width(9)) asuint_4058 (
        .y(_T_432),
        .in(_T_431)
    );
    wire [7:0] estNormNeg_dist;
    TAIL #(.width(9), .n(1)) tail_4059 (
        .y(estNormNeg_dist),
        .in(_T_432)
    );
    wire [31:0] _T_433;
    BITS #(.width(162), .high(75), .low(44)) bits_4060 (
        .y(_T_433),
        .in(sigSum)
    );
    wire _T_435;
    wire [31:0] _WTEMP_564;
    PAD_UNSIGNED #(.width(1), .n(32)) u_pad_4061 (
        .y(_WTEMP_564),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(32)) u_neq_4062 (
        .y(_T_435),
        .a(_T_433),
        .b(_WTEMP_564)
    );
    wire [43:0] _T_436;
    BITS #(.width(162), .high(43), .low(0)) bits_4063 (
        .y(_T_436),
        .in(sigSum)
    );
    wire _T_438;
    wire [43:0] _WTEMP_565;
    PAD_UNSIGNED #(.width(1), .n(44)) u_pad_4064 (
        .y(_WTEMP_565),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(44)) u_neq_4065 (
        .y(_T_438),
        .a(_T_436),
        .b(_WTEMP_565)
    );
    wire [1:0] firstReduceSigSum;
    CAT #(.width_a(1), .width_b(1)) cat_4066 (
        .y(firstReduceSigSum),
        .a(_T_435),
        .b(_T_438)
    );
    wire [161:0] complSigSum;
    BITWISENOT #(.width(162)) bitwisenot_4067 (
        .y(complSigSum),
        .in(sigSum)
    );
    wire [31:0] _T_439;
    BITS #(.width(162), .high(75), .low(44)) bits_4068 (
        .y(_T_439),
        .in(complSigSum)
    );
    wire _T_441;
    wire [31:0] _WTEMP_566;
    PAD_UNSIGNED #(.width(1), .n(32)) u_pad_4069 (
        .y(_WTEMP_566),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(32)) u_neq_4070 (
        .y(_T_441),
        .a(_T_439),
        .b(_WTEMP_566)
    );
    wire [43:0] _T_442;
    BITS #(.width(162), .high(43), .low(0)) bits_4071 (
        .y(_T_442),
        .in(complSigSum)
    );
    wire _T_444;
    wire [43:0] _WTEMP_567;
    PAD_UNSIGNED #(.width(1), .n(44)) u_pad_4072 (
        .y(_WTEMP_567),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(44)) u_neq_4073 (
        .y(_T_444),
        .a(_T_442),
        .b(_WTEMP_567)
    );
    wire [1:0] firstReduceComplSigSum;
    CAT #(.width_a(1), .width_b(1)) cat_4074 (
        .y(firstReduceComplSigSum),
        .a(_T_441),
        .b(_T_444)
    );
    wire _T_445;
    BITWISEOR #(.width(1)) bitwiseor_4075 (
        .y(_T_445),
        .a(io_fromPreMul_CAlignDist_0),
        .b(doSubMags)
    );
    wire [8:0] _T_447;
    wire [7:0] _WTEMP_568;
    PAD_UNSIGNED #(.width(1), .n(8)) u_pad_4076 (
        .y(_WTEMP_568),
        .in(1'h1)
    );
    SUB_UNSIGNED #(.width(8)) u_sub_4077 (
        .y(_T_447),
        .a(io_fromPreMul_CAlignDist),
        .b(_WTEMP_568)
    );
    wire [8:0] _T_448;
    ASUINT #(.width(9)) asuint_4078 (
        .y(_T_448),
        .in(_T_447)
    );
    wire [7:0] _T_449;
    TAIL #(.width(9), .n(1)) tail_4079 (
        .y(_T_449),
        .in(_T_448)
    );
    wire [5:0] _T_450;
    BITS #(.width(8), .high(5), .low(0)) bits_4080 (
        .y(_T_450),
        .in(_T_449)
    );
    wire [7:0] CDom_estNormDist;
    wire [7:0] _WTEMP_569;
    PAD_UNSIGNED #(.width(6), .n(8)) u_pad_4081 (
        .y(_WTEMP_569),
        .in(_T_450)
    );
    MUX_UNSIGNED #(.width(8)) u_mux_4082 (
        .y(CDom_estNormDist),
        .sel(_T_445),
        .a(io_fromPreMul_CAlignDist),
        .b(_WTEMP_569)
    );
    wire _T_452;
    EQ_UNSIGNED #(.width(1)) u_eq_4083 (
        .y(_T_452),
        .a(doSubMags),
        .b(1'h0)
    );
    wire _T_453;
    BITS #(.width(8), .high(5), .low(5)) bits_4084 (
        .y(_T_453),
        .in(CDom_estNormDist)
    );
    wire _T_455;
    EQ_UNSIGNED #(.width(1)) u_eq_4085 (
        .y(_T_455),
        .a(_T_453),
        .b(1'h0)
    );
    wire _T_456;
    BITWISEAND #(.width(1)) bitwiseand_4086 (
        .y(_T_456),
        .a(_T_452),
        .b(_T_455)
    );
    wire [85:0] _T_457;
    BITS #(.width(162), .high(161), .low(76)) bits_4087 (
        .y(_T_457),
        .in(sigSum)
    );
    wire _T_459;
    wire [1:0] _WTEMP_570;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_4088 (
        .y(_WTEMP_570),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(2)) u_neq_4089 (
        .y(_T_459),
        .a(firstReduceSigSum),
        .b(_WTEMP_570)
    );
    wire [86:0] _T_460;
    CAT #(.width_a(86), .width_b(1)) cat_4090 (
        .y(_T_460),
        .a(_T_457),
        .b(_T_459)
    );
    wire [86:0] _T_462;
    wire [86:0] _WTEMP_571;
    PAD_UNSIGNED #(.width(1), .n(87)) u_pad_4091 (
        .y(_WTEMP_571),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(87)) u_mux_4092 (
        .y(_T_462),
        .sel(_T_456),
        .a(_T_460),
        .b(_WTEMP_571)
    );
    wire _T_464;
    EQ_UNSIGNED #(.width(1)) u_eq_4093 (
        .y(_T_464),
        .a(doSubMags),
        .b(1'h0)
    );
    wire _T_465;
    BITS #(.width(8), .high(5), .low(5)) bits_4094 (
        .y(_T_465),
        .in(CDom_estNormDist)
    );
    wire _T_466;
    BITWISEAND #(.width(1)) bitwiseand_4095 (
        .y(_T_466),
        .a(_T_464),
        .b(_T_465)
    );
    wire [85:0] _T_467;
    BITS #(.width(162), .high(129), .low(44)) bits_4096 (
        .y(_T_467),
        .in(sigSum)
    );
    wire _T_468;
    BITS #(.width(2), .high(0), .low(0)) bits_4097 (
        .y(_T_468),
        .in(firstReduceSigSum)
    );
    wire [86:0] _T_469;
    CAT #(.width_a(86), .width_b(1)) cat_4098 (
        .y(_T_469),
        .a(_T_467),
        .b(_T_468)
    );
    wire [86:0] _T_471;
    wire [86:0] _WTEMP_572;
    PAD_UNSIGNED #(.width(1), .n(87)) u_pad_4099 (
        .y(_WTEMP_572),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(87)) u_mux_4100 (
        .y(_T_471),
        .sel(_T_466),
        .a(_T_469),
        .b(_WTEMP_572)
    );
    wire [86:0] _T_472;
    BITWISEOR #(.width(87)) bitwiseor_4101 (
        .y(_T_472),
        .a(_T_462),
        .b(_T_471)
    );
    wire _T_473;
    BITS #(.width(8), .high(5), .low(5)) bits_4102 (
        .y(_T_473),
        .in(CDom_estNormDist)
    );
    wire _T_475;
    EQ_UNSIGNED #(.width(1)) u_eq_4103 (
        .y(_T_475),
        .a(_T_473),
        .b(1'h0)
    );
    wire _T_476;
    BITWISEAND #(.width(1)) bitwiseand_4104 (
        .y(_T_476),
        .a(doSubMags),
        .b(_T_475)
    );
    wire [85:0] _T_477;
    BITS #(.width(162), .high(161), .low(76)) bits_4105 (
        .y(_T_477),
        .in(complSigSum)
    );
    wire _T_479;
    wire [1:0] _WTEMP_573;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_4106 (
        .y(_WTEMP_573),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(2)) u_neq_4107 (
        .y(_T_479),
        .a(firstReduceComplSigSum),
        .b(_WTEMP_573)
    );
    wire [86:0] _T_480;
    CAT #(.width_a(86), .width_b(1)) cat_4108 (
        .y(_T_480),
        .a(_T_477),
        .b(_T_479)
    );
    wire [86:0] _T_482;
    wire [86:0] _WTEMP_574;
    PAD_UNSIGNED #(.width(1), .n(87)) u_pad_4109 (
        .y(_WTEMP_574),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(87)) u_mux_4110 (
        .y(_T_482),
        .sel(_T_476),
        .a(_T_480),
        .b(_WTEMP_574)
    );
    wire [86:0] _T_483;
    BITWISEOR #(.width(87)) bitwiseor_4111 (
        .y(_T_483),
        .a(_T_472),
        .b(_T_482)
    );
    wire _T_484;
    BITS #(.width(8), .high(5), .low(5)) bits_4112 (
        .y(_T_484),
        .in(CDom_estNormDist)
    );
    wire _T_485;
    BITWISEAND #(.width(1)) bitwiseand_4113 (
        .y(_T_485),
        .a(doSubMags),
        .b(_T_484)
    );
    wire [85:0] _T_486;
    BITS #(.width(162), .high(129), .low(44)) bits_4114 (
        .y(_T_486),
        .in(complSigSum)
    );
    wire _T_487;
    BITS #(.width(2), .high(0), .low(0)) bits_4115 (
        .y(_T_487),
        .in(firstReduceComplSigSum)
    );
    wire [86:0] _T_488;
    CAT #(.width_a(86), .width_b(1)) cat_4116 (
        .y(_T_488),
        .a(_T_486),
        .b(_T_487)
    );
    wire [86:0] _T_490;
    wire [86:0] _WTEMP_575;
    PAD_UNSIGNED #(.width(1), .n(87)) u_pad_4117 (
        .y(_WTEMP_575),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(87)) u_mux_4118 (
        .y(_T_490),
        .sel(_T_485),
        .a(_T_488),
        .b(_WTEMP_575)
    );
    wire [86:0] CDom_firstNormAbsSigSum;
    BITWISEOR #(.width(87)) bitwiseor_4119 (
        .y(CDom_firstNormAbsSigSum),
        .a(_T_483),
        .b(_T_490)
    );
    wire [64:0] _T_491;
    BITS #(.width(162), .high(108), .low(44)) bits_4120 (
        .y(_T_491),
        .in(sigSum)
    );
    wire _T_492;
    BITS #(.width(2), .high(0), .low(0)) bits_4121 (
        .y(_T_492),
        .in(firstReduceComplSigSum)
    );
    wire _T_494;
    EQ_UNSIGNED #(.width(1)) u_eq_4122 (
        .y(_T_494),
        .a(_T_492),
        .b(1'h0)
    );
    wire _T_495;
    BITS #(.width(2), .high(0), .low(0)) bits_4123 (
        .y(_T_495),
        .in(firstReduceSigSum)
    );
    wire _T_496;
    MUX_UNSIGNED #(.width(1)) u_mux_4124 (
        .y(_T_496),
        .sel(doSubMags),
        .a(_T_494),
        .b(_T_495)
    );
    wire [65:0] _T_497;
    CAT #(.width_a(65), .width_b(1)) cat_4125 (
        .y(_T_497),
        .a(_T_491),
        .b(_T_496)
    );
    wire [96:0] _T_498;
    BITS #(.width(162), .high(97), .low(1)) bits_4126 (
        .y(_T_498),
        .in(sigSum)
    );
    wire _T_499;
    BITS #(.width(8), .high(4), .low(4)) bits_4127 (
        .y(_T_499),
        .in(estNormNeg_dist)
    );
    wire _T_500;
    BITS #(.width(162), .high(1), .low(1)) bits_4128 (
        .y(_T_500),
        .in(sigSum)
    );
    wire _T_501;
    BITS #(.width(1), .high(0), .low(0)) bits_4129 (
        .y(_T_501),
        .in(doSubMags)
    );
    wire [85:0] _T_504;
    MUX_UNSIGNED #(.width(86)) u_mux_4130 (
        .y(_T_504),
        .sel(_T_501),
        .a(86'h3FFFFFFFFFFFFFFFFFFFFF),
        .b(86'h0)
    );
    wire [86:0] _T_505;
    CAT #(.width_a(1), .width_b(86)) cat_4131 (
        .y(_T_505),
        .a(_T_500),
        .b(_T_504)
    );
    wire [86:0] _T_506;
    wire [86:0] _WTEMP_576;
    PAD_UNSIGNED #(.width(66), .n(87)) u_pad_4132 (
        .y(_WTEMP_576),
        .in(_T_497)
    );
    MUX_UNSIGNED #(.width(87)) u_mux_4133 (
        .y(_T_506),
        .sel(_T_499),
        .a(_WTEMP_576),
        .b(_T_505)
    );
    wire [85:0] _T_507;
    BITS #(.width(162), .high(97), .low(12)) bits_4134 (
        .y(_T_507),
        .in(sigSum)
    );
    wire [10:0] _T_508;
    BITS #(.width(162), .high(11), .low(1)) bits_4135 (
        .y(_T_508),
        .in(complSigSum)
    );
    wire _T_510;
    wire [10:0] _WTEMP_577;
    PAD_UNSIGNED #(.width(1), .n(11)) u_pad_4136 (
        .y(_WTEMP_577),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(11)) u_eq_4137 (
        .y(_T_510),
        .a(_T_508),
        .b(_WTEMP_577)
    );
    wire [10:0] _T_511;
    BITS #(.width(162), .high(11), .low(1)) bits_4138 (
        .y(_T_511),
        .in(sigSum)
    );
    wire _T_513;
    wire [10:0] _WTEMP_578;
    PAD_UNSIGNED #(.width(1), .n(11)) u_pad_4139 (
        .y(_WTEMP_578),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(11)) u_neq_4140 (
        .y(_T_513),
        .a(_T_511),
        .b(_WTEMP_578)
    );
    wire _T_514;
    MUX_UNSIGNED #(.width(1)) u_mux_4141 (
        .y(_T_514),
        .sel(doSubMags),
        .a(_T_510),
        .b(_T_513)
    );
    wire [86:0] _T_515;
    CAT #(.width_a(86), .width_b(1)) cat_4142 (
        .y(_T_515),
        .a(_T_507),
        .b(_T_514)
    );
    wire _T_516;
    BITS #(.width(8), .high(6), .low(6)) bits_4143 (
        .y(_T_516),
        .in(estNormNeg_dist)
    );
    wire _T_517;
    BITS #(.width(8), .high(5), .low(5)) bits_4144 (
        .y(_T_517),
        .in(estNormNeg_dist)
    );
    wire [64:0] _T_518;
    BITS #(.width(162), .high(65), .low(1)) bits_4145 (
        .y(_T_518),
        .in(sigSum)
    );
    wire _T_519;
    BITS #(.width(1), .high(0), .low(0)) bits_4146 (
        .y(_T_519),
        .in(doSubMags)
    );
    wire [21:0] _T_522;
    MUX_UNSIGNED #(.width(22)) u_mux_4147 (
        .y(_T_522),
        .sel(_T_519),
        .a(22'h3FFFFF),
        .b(22'h0)
    );
    wire [86:0] _T_523;
    CAT #(.width_a(65), .width_b(22)) cat_4148 (
        .y(_T_523),
        .a(_T_518),
        .b(_T_522)
    );
    wire [86:0] _T_524;
    MUX_UNSIGNED #(.width(87)) u_mux_4149 (
        .y(_T_524),
        .sel(_T_517),
        .a(_T_523),
        .b(_T_515)
    );
    wire _T_525;
    BITS #(.width(8), .high(5), .low(5)) bits_4150 (
        .y(_T_525),
        .in(estNormNeg_dist)
    );
    wire [32:0] _T_526;
    BITS #(.width(162), .high(33), .low(1)) bits_4151 (
        .y(_T_526),
        .in(sigSum)
    );
    wire _T_527;
    BITS #(.width(1), .high(0), .low(0)) bits_4152 (
        .y(_T_527),
        .in(doSubMags)
    );
    wire [53:0] _T_530;
    MUX_UNSIGNED #(.width(54)) u_mux_4153 (
        .y(_T_530),
        .sel(_T_527),
        .a(54'h3FFFFFFFFFFFFF),
        .b(54'h0)
    );
    wire [86:0] _T_531;
    CAT #(.width_a(33), .width_b(54)) cat_4154 (
        .y(_T_531),
        .a(_T_526),
        .b(_T_530)
    );
    wire [86:0] _T_532;
    MUX_UNSIGNED #(.width(87)) u_mux_4155 (
        .y(_T_532),
        .sel(_T_525),
        .a(_T_506),
        .b(_T_531)
    );
    wire [86:0] notCDom_pos_firstNormAbsSigSum;
    MUX_UNSIGNED #(.width(87)) u_mux_4156 (
        .y(notCDom_pos_firstNormAbsSigSum),
        .sel(_T_516),
        .a(_T_524),
        .b(_T_532)
    );
    wire [63:0] _T_533;
    BITS #(.width(162), .high(107), .low(44)) bits_4157 (
        .y(_T_533),
        .in(complSigSum)
    );
    wire _T_534;
    BITS #(.width(2), .high(0), .low(0)) bits_4158 (
        .y(_T_534),
        .in(firstReduceComplSigSum)
    );
    wire [64:0] _T_535;
    CAT #(.width_a(64), .width_b(1)) cat_4159 (
        .y(_T_535),
        .a(_T_533),
        .b(_T_534)
    );
    wire [96:0] _T_536;
    BITS #(.width(162), .high(97), .low(1)) bits_4160 (
        .y(_T_536),
        .in(complSigSum)
    );
    wire _T_537;
    BITS #(.width(8), .high(4), .low(4)) bits_4161 (
        .y(_T_537),
        .in(estNormNeg_dist)
    );
    wire [1:0] _T_538;
    BITS #(.width(162), .high(2), .low(1)) bits_4162 (
        .y(_T_538),
        .in(complSigSum)
    );
    wire [87:0] _T_539;
    SHL_UNSIGNED #(.width(2), .n(86)) u_shl_4163 (
        .y(_T_539),
        .in(_T_538)
    );
    wire [87:0] _T_540;
    wire [87:0] _WTEMP_579;
    PAD_UNSIGNED #(.width(65), .n(88)) u_pad_4164 (
        .y(_WTEMP_579),
        .in(_T_535)
    );
    MUX_UNSIGNED #(.width(88)) u_mux_4165 (
        .y(_T_540),
        .sel(_T_537),
        .a(_WTEMP_579),
        .b(_T_539)
    );
    wire [86:0] _T_541;
    BITS #(.width(162), .high(98), .low(12)) bits_4166 (
        .y(_T_541),
        .in(complSigSum)
    );
    wire [10:0] _T_542;
    BITS #(.width(162), .high(11), .low(1)) bits_4167 (
        .y(_T_542),
        .in(complSigSum)
    );
    wire _T_544;
    wire [10:0] _WTEMP_580;
    PAD_UNSIGNED #(.width(1), .n(11)) u_pad_4168 (
        .y(_WTEMP_580),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(11)) u_neq_4169 (
        .y(_T_544),
        .a(_T_542),
        .b(_WTEMP_580)
    );
    wire [87:0] _T_545;
    CAT #(.width_a(87), .width_b(1)) cat_4170 (
        .y(_T_545),
        .a(_T_541),
        .b(_T_544)
    );
    wire _T_546;
    BITS #(.width(8), .high(6), .low(6)) bits_4171 (
        .y(_T_546),
        .in(estNormNeg_dist)
    );
    wire _T_547;
    BITS #(.width(8), .high(5), .low(5)) bits_4172 (
        .y(_T_547),
        .in(estNormNeg_dist)
    );
    wire [65:0] _T_548;
    BITS #(.width(162), .high(66), .low(1)) bits_4173 (
        .y(_T_548),
        .in(complSigSum)
    );
    wire [87:0] _T_549;
    SHL_UNSIGNED #(.width(66), .n(22)) u_shl_4174 (
        .y(_T_549),
        .in(_T_548)
    );
    wire [87:0] _T_550;
    MUX_UNSIGNED #(.width(88)) u_mux_4175 (
        .y(_T_550),
        .sel(_T_547),
        .a(_T_549),
        .b(_T_545)
    );
    wire _T_551;
    BITS #(.width(8), .high(5), .low(5)) bits_4176 (
        .y(_T_551),
        .in(estNormNeg_dist)
    );
    wire [33:0] _T_552;
    BITS #(.width(162), .high(34), .low(1)) bits_4177 (
        .y(_T_552),
        .in(complSigSum)
    );
    wire [87:0] _T_553;
    SHL_UNSIGNED #(.width(34), .n(54)) u_shl_4178 (
        .y(_T_553),
        .in(_T_552)
    );
    wire [87:0] _T_554;
    MUX_UNSIGNED #(.width(88)) u_mux_4179 (
        .y(_T_554),
        .sel(_T_551),
        .a(_T_540),
        .b(_T_553)
    );
    wire [87:0] notCDom_neg_cFirstNormAbsSigSum;
    MUX_UNSIGNED #(.width(88)) u_mux_4180 (
        .y(notCDom_neg_cFirstNormAbsSigSum),
        .sel(_T_546),
        .a(_T_550),
        .b(_T_554)
    );
    wire notCDom_signSigSum;
    BITS #(.width(162), .high(109), .low(109)) bits_4181 (
        .y(notCDom_signSigSum),
        .in(sigSum)
    );
    wire _T_556;
    EQ_UNSIGNED #(.width(1)) u_eq_4182 (
        .y(_T_556),
        .a(isZeroC),
        .b(1'h0)
    );
    wire _T_557;
    BITWISEAND #(.width(1)) bitwiseand_4183 (
        .y(_T_557),
        .a(doSubMags),
        .b(_T_556)
    );
    wire doNegSignSum;
    MUX_UNSIGNED #(.width(1)) u_mux_4184 (
        .y(doNegSignSum),
        .sel(io_fromPreMul_isCDominant),
        .a(_T_557),
        .b(notCDom_signSigSum)
    );
    wire [7:0] _T_558;
    assign _T_558 = estNormNeg_dist;
    wire [7:0] estNormDist;
    MUX_UNSIGNED #(.width(8)) u_mux_4185 (
        .y(estNormDist),
        .sel(io_fromPreMul_isCDominant),
        .a(CDom_estNormDist),
        .b(_T_558)
    );
    wire [87:0] _T_559;
    wire [87:0] _WTEMP_581;
    PAD_UNSIGNED #(.width(87), .n(88)) u_pad_4186 (
        .y(_WTEMP_581),
        .in(CDom_firstNormAbsSigSum)
    );
    MUX_UNSIGNED #(.width(88)) u_mux_4187 (
        .y(_T_559),
        .sel(io_fromPreMul_isCDominant),
        .a(_WTEMP_581),
        .b(notCDom_neg_cFirstNormAbsSigSum)
    );
    wire [86:0] _T_560;
    MUX_UNSIGNED #(.width(87)) u_mux_4188 (
        .y(_T_560),
        .sel(io_fromPreMul_isCDominant),
        .a(CDom_firstNormAbsSigSum),
        .b(notCDom_pos_firstNormAbsSigSum)
    );
    wire [87:0] cFirstNormAbsSigSum;
    wire [87:0] _WTEMP_582;
    PAD_UNSIGNED #(.width(87), .n(88)) u_pad_4189 (
        .y(_WTEMP_582),
        .in(_T_560)
    );
    MUX_UNSIGNED #(.width(88)) u_mux_4190 (
        .y(cFirstNormAbsSigSum),
        .sel(notCDom_signSigSum),
        .a(_T_559),
        .b(_WTEMP_582)
    );
    wire _T_562;
    EQ_UNSIGNED #(.width(1)) u_eq_4191 (
        .y(_T_562),
        .a(io_fromPreMul_isCDominant),
        .b(1'h0)
    );
    wire _T_564;
    EQ_UNSIGNED #(.width(1)) u_eq_4192 (
        .y(_T_564),
        .a(notCDom_signSigSum),
        .b(1'h0)
    );
    wire _T_565;
    BITWISEAND #(.width(1)) bitwiseand_4193 (
        .y(_T_565),
        .a(_T_562),
        .b(_T_564)
    );
    wire doIncrSig;
    BITWISEAND #(.width(1)) bitwiseand_4194 (
        .y(doIncrSig),
        .a(_T_565),
        .b(doSubMags)
    );
    wire [4:0] estNormDist_5;
    BITS #(.width(8), .high(4), .low(0)) bits_4195 (
        .y(estNormDist_5),
        .in(estNormDist)
    );
    wire [4:0] normTo2ShiftDist;
    BITWISENOT #(.width(5)) bitwisenot_4196 (
        .y(normTo2ShiftDist),
        .in(estNormDist_5)
    );
    wire [32:0] _T_567;
    DSHR_SIGNED #(.width_in(33), .width_n(5)) s_dshr_4197 (
        .y(_T_567),
        .in(-33'sh100000000),
        .n(normTo2ShiftDist)
    );
    wire [30:0] _T_568;
    BITS #(.width(33), .high(31), .low(1)) bits_4198 (
        .y(_T_568),
        .in(_T_567)
    );
    wire [15:0] _T_569;
    BITS #(.width(31), .high(15), .low(0)) bits_4199 (
        .y(_T_569),
        .in(_T_568)
    );
    wire [15:0] _T_572;
    assign _T_572 = 16'hFF00;
    wire [15:0] _T_573;
    assign _T_573 = 16'hFF;
    wire [7:0] _T_574;
    SHR_UNSIGNED #(.width(16), .n(8)) u_shr_4200 (
        .y(_T_574),
        .in(_T_569)
    );
    wire [15:0] _T_575;
    wire [15:0] _WTEMP_583;
    PAD_UNSIGNED #(.width(8), .n(16)) u_pad_4201 (
        .y(_WTEMP_583),
        .in(_T_574)
    );
    BITWISEAND #(.width(16)) bitwiseand_4202 (
        .y(_T_575),
        .a(_WTEMP_583),
        .b(_T_573)
    );
    wire [7:0] _T_576;
    BITS #(.width(16), .high(7), .low(0)) bits_4203 (
        .y(_T_576),
        .in(_T_569)
    );
    wire [15:0] _T_577;
    SHL_UNSIGNED #(.width(8), .n(8)) u_shl_4204 (
        .y(_T_577),
        .in(_T_576)
    );
    wire [15:0] _T_578;
    assign _T_578 = 16'hFF00;
    wire [15:0] _T_579;
    BITWISEAND #(.width(16)) bitwiseand_4205 (
        .y(_T_579),
        .a(_T_577),
        .b(_T_578)
    );
    wire [15:0] _T_580;
    BITWISEOR #(.width(16)) bitwiseor_4206 (
        .y(_T_580),
        .a(_T_575),
        .b(_T_579)
    );
    wire [11:0] _T_581;
    assign _T_581 = 12'hFF;
    wire [15:0] _T_582;
    assign _T_582 = 16'hFF0;
    wire [15:0] _T_583;
    assign _T_583 = 16'hF0F;
    wire [11:0] _T_584;
    SHR_UNSIGNED #(.width(16), .n(4)) u_shr_4207 (
        .y(_T_584),
        .in(_T_580)
    );
    wire [15:0] _T_585;
    wire [15:0] _WTEMP_584;
    PAD_UNSIGNED #(.width(12), .n(16)) u_pad_4208 (
        .y(_WTEMP_584),
        .in(_T_584)
    );
    BITWISEAND #(.width(16)) bitwiseand_4209 (
        .y(_T_585),
        .a(_WTEMP_584),
        .b(_T_583)
    );
    wire [11:0] _T_586;
    BITS #(.width(16), .high(11), .low(0)) bits_4210 (
        .y(_T_586),
        .in(_T_580)
    );
    wire [15:0] _T_587;
    SHL_UNSIGNED #(.width(12), .n(4)) u_shl_4211 (
        .y(_T_587),
        .in(_T_586)
    );
    wire [15:0] _T_588;
    assign _T_588 = 16'hF0F0;
    wire [15:0] _T_589;
    BITWISEAND #(.width(16)) bitwiseand_4212 (
        .y(_T_589),
        .a(_T_587),
        .b(_T_588)
    );
    wire [15:0] _T_590;
    BITWISEOR #(.width(16)) bitwiseor_4213 (
        .y(_T_590),
        .a(_T_585),
        .b(_T_589)
    );
    wire [13:0] _T_591;
    assign _T_591 = 14'hF0F;
    wire [15:0] _T_592;
    assign _T_592 = 16'h3C3C;
    wire [15:0] _T_593;
    assign _T_593 = 16'h3333;
    wire [13:0] _T_594;
    SHR_UNSIGNED #(.width(16), .n(2)) u_shr_4214 (
        .y(_T_594),
        .in(_T_590)
    );
    wire [15:0] _T_595;
    wire [15:0] _WTEMP_585;
    PAD_UNSIGNED #(.width(14), .n(16)) u_pad_4215 (
        .y(_WTEMP_585),
        .in(_T_594)
    );
    BITWISEAND #(.width(16)) bitwiseand_4216 (
        .y(_T_595),
        .a(_WTEMP_585),
        .b(_T_593)
    );
    wire [13:0] _T_596;
    BITS #(.width(16), .high(13), .low(0)) bits_4217 (
        .y(_T_596),
        .in(_T_590)
    );
    wire [15:0] _T_597;
    SHL_UNSIGNED #(.width(14), .n(2)) u_shl_4218 (
        .y(_T_597),
        .in(_T_596)
    );
    wire [15:0] _T_598;
    assign _T_598 = 16'hCCCC;
    wire [15:0] _T_599;
    BITWISEAND #(.width(16)) bitwiseand_4219 (
        .y(_T_599),
        .a(_T_597),
        .b(_T_598)
    );
    wire [15:0] _T_600;
    BITWISEOR #(.width(16)) bitwiseor_4220 (
        .y(_T_600),
        .a(_T_595),
        .b(_T_599)
    );
    wire [14:0] _T_601;
    assign _T_601 = 15'h3333;
    wire [15:0] _T_602;
    assign _T_602 = 16'h6666;
    wire [15:0] _T_603;
    assign _T_603 = 16'h5555;
    wire [14:0] _T_604;
    SHR_UNSIGNED #(.width(16), .n(1)) u_shr_4221 (
        .y(_T_604),
        .in(_T_600)
    );
    wire [15:0] _T_605;
    wire [15:0] _WTEMP_586;
    PAD_UNSIGNED #(.width(15), .n(16)) u_pad_4222 (
        .y(_WTEMP_586),
        .in(_T_604)
    );
    BITWISEAND #(.width(16)) bitwiseand_4223 (
        .y(_T_605),
        .a(_WTEMP_586),
        .b(_T_603)
    );
    wire [14:0] _T_606;
    BITS #(.width(16), .high(14), .low(0)) bits_4224 (
        .y(_T_606),
        .in(_T_600)
    );
    wire [15:0] _T_607;
    SHL_UNSIGNED #(.width(15), .n(1)) u_shl_4225 (
        .y(_T_607),
        .in(_T_606)
    );
    wire [15:0] _T_608;
    assign _T_608 = 16'hAAAA;
    wire [15:0] _T_609;
    BITWISEAND #(.width(16)) bitwiseand_4226 (
        .y(_T_609),
        .a(_T_607),
        .b(_T_608)
    );
    wire [15:0] _T_610;
    BITWISEOR #(.width(16)) bitwiseor_4227 (
        .y(_T_610),
        .a(_T_605),
        .b(_T_609)
    );
    wire [14:0] _T_611;
    BITS #(.width(31), .high(30), .low(16)) bits_4228 (
        .y(_T_611),
        .in(_T_568)
    );
    wire [7:0] _T_612;
    BITS #(.width(15), .high(7), .low(0)) bits_4229 (
        .y(_T_612),
        .in(_T_611)
    );
    wire [7:0] _T_615;
    assign _T_615 = 8'hF0;
    wire [7:0] _T_616;
    assign _T_616 = 8'hF;
    wire [3:0] _T_617;
    SHR_UNSIGNED #(.width(8), .n(4)) u_shr_4230 (
        .y(_T_617),
        .in(_T_612)
    );
    wire [7:0] _T_618;
    wire [7:0] _WTEMP_587;
    PAD_UNSIGNED #(.width(4), .n(8)) u_pad_4231 (
        .y(_WTEMP_587),
        .in(_T_617)
    );
    BITWISEAND #(.width(8)) bitwiseand_4232 (
        .y(_T_618),
        .a(_WTEMP_587),
        .b(_T_616)
    );
    wire [3:0] _T_619;
    BITS #(.width(8), .high(3), .low(0)) bits_4233 (
        .y(_T_619),
        .in(_T_612)
    );
    wire [7:0] _T_620;
    SHL_UNSIGNED #(.width(4), .n(4)) u_shl_4234 (
        .y(_T_620),
        .in(_T_619)
    );
    wire [7:0] _T_621;
    assign _T_621 = 8'hF0;
    wire [7:0] _T_622;
    BITWISEAND #(.width(8)) bitwiseand_4235 (
        .y(_T_622),
        .a(_T_620),
        .b(_T_621)
    );
    wire [7:0] _T_623;
    BITWISEOR #(.width(8)) bitwiseor_4236 (
        .y(_T_623),
        .a(_T_618),
        .b(_T_622)
    );
    wire [5:0] _T_624;
    assign _T_624 = 6'hF;
    wire [7:0] _T_625;
    assign _T_625 = 8'h3C;
    wire [7:0] _T_626;
    assign _T_626 = 8'h33;
    wire [5:0] _T_627;
    SHR_UNSIGNED #(.width(8), .n(2)) u_shr_4237 (
        .y(_T_627),
        .in(_T_623)
    );
    wire [7:0] _T_628;
    wire [7:0] _WTEMP_588;
    PAD_UNSIGNED #(.width(6), .n(8)) u_pad_4238 (
        .y(_WTEMP_588),
        .in(_T_627)
    );
    BITWISEAND #(.width(8)) bitwiseand_4239 (
        .y(_T_628),
        .a(_WTEMP_588),
        .b(_T_626)
    );
    wire [5:0] _T_629;
    BITS #(.width(8), .high(5), .low(0)) bits_4240 (
        .y(_T_629),
        .in(_T_623)
    );
    wire [7:0] _T_630;
    SHL_UNSIGNED #(.width(6), .n(2)) u_shl_4241 (
        .y(_T_630),
        .in(_T_629)
    );
    wire [7:0] _T_631;
    assign _T_631 = 8'hCC;
    wire [7:0] _T_632;
    BITWISEAND #(.width(8)) bitwiseand_4242 (
        .y(_T_632),
        .a(_T_630),
        .b(_T_631)
    );
    wire [7:0] _T_633;
    BITWISEOR #(.width(8)) bitwiseor_4243 (
        .y(_T_633),
        .a(_T_628),
        .b(_T_632)
    );
    wire [6:0] _T_634;
    assign _T_634 = 7'h33;
    wire [7:0] _T_635;
    assign _T_635 = 8'h66;
    wire [7:0] _T_636;
    assign _T_636 = 8'h55;
    wire [6:0] _T_637;
    SHR_UNSIGNED #(.width(8), .n(1)) u_shr_4244 (
        .y(_T_637),
        .in(_T_633)
    );
    wire [7:0] _T_638;
    wire [7:0] _WTEMP_589;
    PAD_UNSIGNED #(.width(7), .n(8)) u_pad_4245 (
        .y(_WTEMP_589),
        .in(_T_637)
    );
    BITWISEAND #(.width(8)) bitwiseand_4246 (
        .y(_T_638),
        .a(_WTEMP_589),
        .b(_T_636)
    );
    wire [6:0] _T_639;
    BITS #(.width(8), .high(6), .low(0)) bits_4247 (
        .y(_T_639),
        .in(_T_633)
    );
    wire [7:0] _T_640;
    SHL_UNSIGNED #(.width(7), .n(1)) u_shl_4248 (
        .y(_T_640),
        .in(_T_639)
    );
    wire [7:0] _T_641;
    assign _T_641 = 8'hAA;
    wire [7:0] _T_642;
    BITWISEAND #(.width(8)) bitwiseand_4249 (
        .y(_T_642),
        .a(_T_640),
        .b(_T_641)
    );
    wire [7:0] _T_643;
    BITWISEOR #(.width(8)) bitwiseor_4250 (
        .y(_T_643),
        .a(_T_638),
        .b(_T_642)
    );
    wire [6:0] _T_644;
    BITS #(.width(15), .high(14), .low(8)) bits_4251 (
        .y(_T_644),
        .in(_T_611)
    );
    wire [3:0] _T_645;
    BITS #(.width(7), .high(3), .low(0)) bits_4252 (
        .y(_T_645),
        .in(_T_644)
    );
    wire [1:0] _T_646;
    BITS #(.width(4), .high(1), .low(0)) bits_4253 (
        .y(_T_646),
        .in(_T_645)
    );
    wire _T_647;
    BITS #(.width(2), .high(0), .low(0)) bits_4254 (
        .y(_T_647),
        .in(_T_646)
    );
    wire _T_648;
    BITS #(.width(2), .high(1), .low(1)) bits_4255 (
        .y(_T_648),
        .in(_T_646)
    );
    wire [1:0] _T_649;
    CAT #(.width_a(1), .width_b(1)) cat_4256 (
        .y(_T_649),
        .a(_T_647),
        .b(_T_648)
    );
    wire [1:0] _T_650;
    BITS #(.width(4), .high(3), .low(2)) bits_4257 (
        .y(_T_650),
        .in(_T_645)
    );
    wire _T_651;
    BITS #(.width(2), .high(0), .low(0)) bits_4258 (
        .y(_T_651),
        .in(_T_650)
    );
    wire _T_652;
    BITS #(.width(2), .high(1), .low(1)) bits_4259 (
        .y(_T_652),
        .in(_T_650)
    );
    wire [1:0] _T_653;
    CAT #(.width_a(1), .width_b(1)) cat_4260 (
        .y(_T_653),
        .a(_T_651),
        .b(_T_652)
    );
    wire [3:0] _T_654;
    CAT #(.width_a(2), .width_b(2)) cat_4261 (
        .y(_T_654),
        .a(_T_649),
        .b(_T_653)
    );
    wire [2:0] _T_655;
    BITS #(.width(7), .high(6), .low(4)) bits_4262 (
        .y(_T_655),
        .in(_T_644)
    );
    wire [1:0] _T_656;
    BITS #(.width(3), .high(1), .low(0)) bits_4263 (
        .y(_T_656),
        .in(_T_655)
    );
    wire _T_657;
    BITS #(.width(2), .high(0), .low(0)) bits_4264 (
        .y(_T_657),
        .in(_T_656)
    );
    wire _T_658;
    BITS #(.width(2), .high(1), .low(1)) bits_4265 (
        .y(_T_658),
        .in(_T_656)
    );
    wire [1:0] _T_659;
    CAT #(.width_a(1), .width_b(1)) cat_4266 (
        .y(_T_659),
        .a(_T_657),
        .b(_T_658)
    );
    wire _T_660;
    BITS #(.width(3), .high(2), .low(2)) bits_4267 (
        .y(_T_660),
        .in(_T_655)
    );
    wire [2:0] _T_661;
    CAT #(.width_a(2), .width_b(1)) cat_4268 (
        .y(_T_661),
        .a(_T_659),
        .b(_T_660)
    );
    wire [6:0] _T_662;
    CAT #(.width_a(4), .width_b(3)) cat_4269 (
        .y(_T_662),
        .a(_T_654),
        .b(_T_661)
    );
    wire [14:0] _T_663;
    CAT #(.width_a(8), .width_b(7)) cat_4270 (
        .y(_T_663),
        .a(_T_643),
        .b(_T_662)
    );
    wire [30:0] _T_664;
    CAT #(.width_a(16), .width_b(15)) cat_4271 (
        .y(_T_664),
        .a(_T_610),
        .b(_T_663)
    );
    wire [31:0] absSigSumExtraMask;
    CAT #(.width_a(31), .width_b(1)) cat_4272 (
        .y(absSigSumExtraMask),
        .a(_T_664),
        .b(1'h1)
    );
    wire [86:0] _T_666;
    BITS #(.width(88), .high(87), .low(1)) bits_4273 (
        .y(_T_666),
        .in(cFirstNormAbsSigSum)
    );
    wire [86:0] _T_667;
    DSHR_UNSIGNED #(.width_in(87), .width_n(5)) u_dshr_4274 (
        .y(_T_667),
        .in(_T_666),
        .n(normTo2ShiftDist)
    );
    wire [31:0] _T_668;
    BITS #(.width(88), .high(31), .low(0)) bits_4275 (
        .y(_T_668),
        .in(cFirstNormAbsSigSum)
    );
    wire [31:0] _T_669;
    BITWISENOT #(.width(32)) bitwisenot_4276 (
        .y(_T_669),
        .in(_T_668)
    );
    wire [31:0] _T_670;
    BITWISEAND #(.width(32)) bitwiseand_4277 (
        .y(_T_670),
        .a(_T_669),
        .b(absSigSumExtraMask)
    );
    wire _T_672;
    wire [31:0] _WTEMP_590;
    PAD_UNSIGNED #(.width(1), .n(32)) u_pad_4278 (
        .y(_WTEMP_590),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(32)) u_eq_4279 (
        .y(_T_672),
        .a(_T_670),
        .b(_WTEMP_590)
    );
    wire [31:0] _T_673;
    BITS #(.width(88), .high(31), .low(0)) bits_4280 (
        .y(_T_673),
        .in(cFirstNormAbsSigSum)
    );
    wire [31:0] _T_674;
    BITWISEAND #(.width(32)) bitwiseand_4281 (
        .y(_T_674),
        .a(_T_673),
        .b(absSigSumExtraMask)
    );
    wire _T_676;
    wire [31:0] _WTEMP_591;
    PAD_UNSIGNED #(.width(1), .n(32)) u_pad_4282 (
        .y(_WTEMP_591),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(32)) u_neq_4283 (
        .y(_T_676),
        .a(_T_674),
        .b(_WTEMP_591)
    );
    wire _T_677;
    MUX_UNSIGNED #(.width(1)) u_mux_4284 (
        .y(_T_677),
        .sel(doIncrSig),
        .a(_T_672),
        .b(_T_676)
    );
    wire [87:0] _T_678;
    CAT #(.width_a(87), .width_b(1)) cat_4285 (
        .y(_T_678),
        .a(_T_667),
        .b(_T_677)
    );
    wire [56:0] sigX3;
    BITS #(.width(88), .high(56), .low(0)) bits_4286 (
        .y(sigX3),
        .in(_T_678)
    );
    wire [1:0] _T_679;
    BITS #(.width(57), .high(56), .low(55)) bits_4287 (
        .y(_T_679),
        .in(sigX3)
    );
    wire sigX3Shift1;
    wire [1:0] _WTEMP_592;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_4288 (
        .y(_WTEMP_592),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(2)) u_eq_4289 (
        .y(sigX3Shift1),
        .a(_T_679),
        .b(_WTEMP_592)
    );
    wire [14:0] _T_681;
    wire [13:0] _WTEMP_593;
    PAD_UNSIGNED #(.width(8), .n(14)) u_pad_4290 (
        .y(_WTEMP_593),
        .in(estNormDist)
    );
    SUB_UNSIGNED #(.width(14)) u_sub_4291 (
        .y(_T_681),
        .a(io_fromPreMul_sExpSum),
        .b(_WTEMP_593)
    );
    wire [14:0] _T_682;
    ASUINT #(.width(15)) asuint_4292 (
        .y(_T_682),
        .in(_T_681)
    );
    wire [13:0] sExpX3;
    TAIL #(.width(15), .n(1)) tail_4293 (
        .y(sExpX3),
        .in(_T_682)
    );
    wire [2:0] _T_683;
    BITS #(.width(57), .high(56), .low(54)) bits_4294 (
        .y(_T_683),
        .in(sigX3)
    );
    wire isZeroY;
    wire [2:0] _WTEMP_594;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_4295 (
        .y(_WTEMP_594),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(3)) u_eq_4296 (
        .y(isZeroY),
        .a(_T_683),
        .b(_WTEMP_594)
    );
    wire _T_685;
    BITWISEXOR #(.width(1)) bitwisexor_4297 (
        .y(_T_685),
        .a(io_fromPreMul_signProd),
        .b(doNegSignSum)
    );
    wire signY;
    MUX_UNSIGNED #(.width(1)) u_mux_4298 (
        .y(signY),
        .sel(isZeroY),
        .a(signZeroNotEqOpSigns),
        .b(_T_685)
    );
    wire [12:0] sExpX3_13;
    BITS #(.width(14), .high(12), .low(0)) bits_4299 (
        .y(sExpX3_13),
        .in(sExpX3)
    );
    wire _T_686;
    BITS #(.width(14), .high(13), .low(13)) bits_4300 (
        .y(_T_686),
        .in(sExpX3)
    );
    wire _T_687;
    BITS #(.width(1), .high(0), .low(0)) bits_4301 (
        .y(_T_687),
        .in(_T_686)
    );
    wire [55:0] _T_690;
    MUX_UNSIGNED #(.width(56)) u_mux_4302 (
        .y(_T_690),
        .sel(_T_687),
        .a(56'hFFFFFFFFFFFFFF),
        .b(56'h0)
    );
    wire [12:0] _T_691;
    BITWISENOT #(.width(13)) bitwisenot_4303 (
        .y(_T_691),
        .in(sExpX3_13)
    );
    wire _T_692;
    BITS #(.width(13), .high(12), .low(12)) bits_4304 (
        .y(_T_692),
        .in(_T_691)
    );
    wire [11:0] _T_693;
    BITS #(.width(13), .high(11), .low(0)) bits_4305 (
        .y(_T_693),
        .in(_T_691)
    );
    wire _T_694;
    BITS #(.width(12), .high(11), .low(11)) bits_4306 (
        .y(_T_694),
        .in(_T_693)
    );
    wire [10:0] _T_695;
    BITS #(.width(12), .high(10), .low(0)) bits_4307 (
        .y(_T_695),
        .in(_T_693)
    );
    wire _T_696;
    BITS #(.width(11), .high(10), .low(10)) bits_4308 (
        .y(_T_696),
        .in(_T_695)
    );
    wire [9:0] _T_697;
    BITS #(.width(11), .high(9), .low(0)) bits_4309 (
        .y(_T_697),
        .in(_T_695)
    );
    wire _T_698;
    BITS #(.width(10), .high(9), .low(9)) bits_4310 (
        .y(_T_698),
        .in(_T_697)
    );
    wire [8:0] _T_699;
    BITS #(.width(10), .high(8), .low(0)) bits_4311 (
        .y(_T_699),
        .in(_T_697)
    );
    wire _T_701;
    BITS #(.width(9), .high(8), .low(8)) bits_4312 (
        .y(_T_701),
        .in(_T_699)
    );
    wire [7:0] _T_702;
    BITS #(.width(9), .high(7), .low(0)) bits_4313 (
        .y(_T_702),
        .in(_T_699)
    );
    wire _T_704;
    BITS #(.width(8), .high(7), .low(7)) bits_4314 (
        .y(_T_704),
        .in(_T_702)
    );
    wire [6:0] _T_705;
    BITS #(.width(8), .high(6), .low(0)) bits_4315 (
        .y(_T_705),
        .in(_T_702)
    );
    wire _T_707;
    BITS #(.width(7), .high(6), .low(6)) bits_4316 (
        .y(_T_707),
        .in(_T_705)
    );
    wire [5:0] _T_708;
    BITS #(.width(7), .high(5), .low(0)) bits_4317 (
        .y(_T_708),
        .in(_T_705)
    );
    wire [64:0] _T_711;
    DSHR_SIGNED #(.width_in(65), .width_n(6)) s_dshr_4318 (
        .y(_T_711),
        .in(-65'sh10000000000000000),
        .n(_T_708)
    );
    wire [49:0] _T_712;
    BITS #(.width(65), .high(63), .low(14)) bits_4319 (
        .y(_T_712),
        .in(_T_711)
    );
    wire [31:0] _T_713;
    BITS #(.width(50), .high(31), .low(0)) bits_4320 (
        .y(_T_713),
        .in(_T_712)
    );
    wire [31:0] _T_716;
    assign _T_716 = 32'hFFFF0000;
    wire [31:0] _T_717;
    assign _T_717 = 32'hFFFF;
    wire [15:0] _T_718;
    SHR_UNSIGNED #(.width(32), .n(16)) u_shr_4321 (
        .y(_T_718),
        .in(_T_713)
    );
    wire [31:0] _T_719;
    wire [31:0] _WTEMP_595;
    PAD_UNSIGNED #(.width(16), .n(32)) u_pad_4322 (
        .y(_WTEMP_595),
        .in(_T_718)
    );
    BITWISEAND #(.width(32)) bitwiseand_4323 (
        .y(_T_719),
        .a(_WTEMP_595),
        .b(_T_717)
    );
    wire [15:0] _T_720;
    BITS #(.width(32), .high(15), .low(0)) bits_4324 (
        .y(_T_720),
        .in(_T_713)
    );
    wire [31:0] _T_721;
    SHL_UNSIGNED #(.width(16), .n(16)) u_shl_4325 (
        .y(_T_721),
        .in(_T_720)
    );
    wire [31:0] _T_722;
    assign _T_722 = 32'hFFFF0000;
    wire [31:0] _T_723;
    BITWISEAND #(.width(32)) bitwiseand_4326 (
        .y(_T_723),
        .a(_T_721),
        .b(_T_722)
    );
    wire [31:0] _T_724;
    BITWISEOR #(.width(32)) bitwiseor_4327 (
        .y(_T_724),
        .a(_T_719),
        .b(_T_723)
    );
    wire [23:0] _T_725;
    assign _T_725 = 24'hFFFF;
    wire [31:0] _T_726;
    assign _T_726 = 32'hFFFF00;
    wire [31:0] _T_727;
    assign _T_727 = 32'hFF00FF;
    wire [23:0] _T_728;
    SHR_UNSIGNED #(.width(32), .n(8)) u_shr_4328 (
        .y(_T_728),
        .in(_T_724)
    );
    wire [31:0] _T_729;
    wire [31:0] _WTEMP_596;
    PAD_UNSIGNED #(.width(24), .n(32)) u_pad_4329 (
        .y(_WTEMP_596),
        .in(_T_728)
    );
    BITWISEAND #(.width(32)) bitwiseand_4330 (
        .y(_T_729),
        .a(_WTEMP_596),
        .b(_T_727)
    );
    wire [23:0] _T_730;
    BITS #(.width(32), .high(23), .low(0)) bits_4331 (
        .y(_T_730),
        .in(_T_724)
    );
    wire [31:0] _T_731;
    SHL_UNSIGNED #(.width(24), .n(8)) u_shl_4332 (
        .y(_T_731),
        .in(_T_730)
    );
    wire [31:0] _T_732;
    assign _T_732 = 32'hFF00FF00;
    wire [31:0] _T_733;
    BITWISEAND #(.width(32)) bitwiseand_4333 (
        .y(_T_733),
        .a(_T_731),
        .b(_T_732)
    );
    wire [31:0] _T_734;
    BITWISEOR #(.width(32)) bitwiseor_4334 (
        .y(_T_734),
        .a(_T_729),
        .b(_T_733)
    );
    wire [27:0] _T_735;
    assign _T_735 = 28'hFF00FF;
    wire [31:0] _T_736;
    assign _T_736 = 32'hFF00FF0;
    wire [31:0] _T_737;
    assign _T_737 = 32'hF0F0F0F;
    wire [27:0] _T_738;
    SHR_UNSIGNED #(.width(32), .n(4)) u_shr_4335 (
        .y(_T_738),
        .in(_T_734)
    );
    wire [31:0] _T_739;
    wire [31:0] _WTEMP_597;
    PAD_UNSIGNED #(.width(28), .n(32)) u_pad_4336 (
        .y(_WTEMP_597),
        .in(_T_738)
    );
    BITWISEAND #(.width(32)) bitwiseand_4337 (
        .y(_T_739),
        .a(_WTEMP_597),
        .b(_T_737)
    );
    wire [27:0] _T_740;
    BITS #(.width(32), .high(27), .low(0)) bits_4338 (
        .y(_T_740),
        .in(_T_734)
    );
    wire [31:0] _T_741;
    SHL_UNSIGNED #(.width(28), .n(4)) u_shl_4339 (
        .y(_T_741),
        .in(_T_740)
    );
    wire [31:0] _T_742;
    assign _T_742 = 32'hF0F0F0F0;
    wire [31:0] _T_743;
    BITWISEAND #(.width(32)) bitwiseand_4340 (
        .y(_T_743),
        .a(_T_741),
        .b(_T_742)
    );
    wire [31:0] _T_744;
    BITWISEOR #(.width(32)) bitwiseor_4341 (
        .y(_T_744),
        .a(_T_739),
        .b(_T_743)
    );
    wire [29:0] _T_745;
    assign _T_745 = 30'hF0F0F0F;
    wire [31:0] _T_746;
    assign _T_746 = 32'h3C3C3C3C;
    wire [31:0] _T_747;
    assign _T_747 = 32'h33333333;
    wire [29:0] _T_748;
    SHR_UNSIGNED #(.width(32), .n(2)) u_shr_4342 (
        .y(_T_748),
        .in(_T_744)
    );
    wire [31:0] _T_749;
    wire [31:0] _WTEMP_598;
    PAD_UNSIGNED #(.width(30), .n(32)) u_pad_4343 (
        .y(_WTEMP_598),
        .in(_T_748)
    );
    BITWISEAND #(.width(32)) bitwiseand_4344 (
        .y(_T_749),
        .a(_WTEMP_598),
        .b(_T_747)
    );
    wire [29:0] _T_750;
    BITS #(.width(32), .high(29), .low(0)) bits_4345 (
        .y(_T_750),
        .in(_T_744)
    );
    wire [31:0] _T_751;
    SHL_UNSIGNED #(.width(30), .n(2)) u_shl_4346 (
        .y(_T_751),
        .in(_T_750)
    );
    wire [31:0] _T_752;
    assign _T_752 = 32'hCCCCCCCC;
    wire [31:0] _T_753;
    BITWISEAND #(.width(32)) bitwiseand_4347 (
        .y(_T_753),
        .a(_T_751),
        .b(_T_752)
    );
    wire [31:0] _T_754;
    BITWISEOR #(.width(32)) bitwiseor_4348 (
        .y(_T_754),
        .a(_T_749),
        .b(_T_753)
    );
    wire [30:0] _T_755;
    assign _T_755 = 31'h33333333;
    wire [31:0] _T_756;
    assign _T_756 = 32'h66666666;
    wire [31:0] _T_757;
    assign _T_757 = 32'h55555555;
    wire [30:0] _T_758;
    SHR_UNSIGNED #(.width(32), .n(1)) u_shr_4349 (
        .y(_T_758),
        .in(_T_754)
    );
    wire [31:0] _T_759;
    wire [31:0] _WTEMP_599;
    PAD_UNSIGNED #(.width(31), .n(32)) u_pad_4350 (
        .y(_WTEMP_599),
        .in(_T_758)
    );
    BITWISEAND #(.width(32)) bitwiseand_4351 (
        .y(_T_759),
        .a(_WTEMP_599),
        .b(_T_757)
    );
    wire [30:0] _T_760;
    BITS #(.width(32), .high(30), .low(0)) bits_4352 (
        .y(_T_760),
        .in(_T_754)
    );
    wire [31:0] _T_761;
    SHL_UNSIGNED #(.width(31), .n(1)) u_shl_4353 (
        .y(_T_761),
        .in(_T_760)
    );
    wire [31:0] _T_762;
    assign _T_762 = 32'hAAAAAAAA;
    wire [31:0] _T_763;
    BITWISEAND #(.width(32)) bitwiseand_4354 (
        .y(_T_763),
        .a(_T_761),
        .b(_T_762)
    );
    wire [31:0] _T_764;
    BITWISEOR #(.width(32)) bitwiseor_4355 (
        .y(_T_764),
        .a(_T_759),
        .b(_T_763)
    );
    wire [17:0] _T_765;
    BITS #(.width(50), .high(49), .low(32)) bits_4356 (
        .y(_T_765),
        .in(_T_712)
    );
    wire [15:0] _T_766;
    BITS #(.width(18), .high(15), .low(0)) bits_4357 (
        .y(_T_766),
        .in(_T_765)
    );
    wire [15:0] _T_769;
    assign _T_769 = 16'hFF00;
    wire [15:0] _T_770;
    assign _T_770 = 16'hFF;
    wire [7:0] _T_771;
    SHR_UNSIGNED #(.width(16), .n(8)) u_shr_4358 (
        .y(_T_771),
        .in(_T_766)
    );
    wire [15:0] _T_772;
    wire [15:0] _WTEMP_600;
    PAD_UNSIGNED #(.width(8), .n(16)) u_pad_4359 (
        .y(_WTEMP_600),
        .in(_T_771)
    );
    BITWISEAND #(.width(16)) bitwiseand_4360 (
        .y(_T_772),
        .a(_WTEMP_600),
        .b(_T_770)
    );
    wire [7:0] _T_773;
    BITS #(.width(16), .high(7), .low(0)) bits_4361 (
        .y(_T_773),
        .in(_T_766)
    );
    wire [15:0] _T_774;
    SHL_UNSIGNED #(.width(8), .n(8)) u_shl_4362 (
        .y(_T_774),
        .in(_T_773)
    );
    wire [15:0] _T_775;
    assign _T_775 = 16'hFF00;
    wire [15:0] _T_776;
    BITWISEAND #(.width(16)) bitwiseand_4363 (
        .y(_T_776),
        .a(_T_774),
        .b(_T_775)
    );
    wire [15:0] _T_777;
    BITWISEOR #(.width(16)) bitwiseor_4364 (
        .y(_T_777),
        .a(_T_772),
        .b(_T_776)
    );
    wire [11:0] _T_778;
    assign _T_778 = 12'hFF;
    wire [15:0] _T_779;
    assign _T_779 = 16'hFF0;
    wire [15:0] _T_780;
    assign _T_780 = 16'hF0F;
    wire [11:0] _T_781;
    SHR_UNSIGNED #(.width(16), .n(4)) u_shr_4365 (
        .y(_T_781),
        .in(_T_777)
    );
    wire [15:0] _T_782;
    wire [15:0] _WTEMP_601;
    PAD_UNSIGNED #(.width(12), .n(16)) u_pad_4366 (
        .y(_WTEMP_601),
        .in(_T_781)
    );
    BITWISEAND #(.width(16)) bitwiseand_4367 (
        .y(_T_782),
        .a(_WTEMP_601),
        .b(_T_780)
    );
    wire [11:0] _T_783;
    BITS #(.width(16), .high(11), .low(0)) bits_4368 (
        .y(_T_783),
        .in(_T_777)
    );
    wire [15:0] _T_784;
    SHL_UNSIGNED #(.width(12), .n(4)) u_shl_4369 (
        .y(_T_784),
        .in(_T_783)
    );
    wire [15:0] _T_785;
    assign _T_785 = 16'hF0F0;
    wire [15:0] _T_786;
    BITWISEAND #(.width(16)) bitwiseand_4370 (
        .y(_T_786),
        .a(_T_784),
        .b(_T_785)
    );
    wire [15:0] _T_787;
    BITWISEOR #(.width(16)) bitwiseor_4371 (
        .y(_T_787),
        .a(_T_782),
        .b(_T_786)
    );
    wire [13:0] _T_788;
    assign _T_788 = 14'hF0F;
    wire [15:0] _T_789;
    assign _T_789 = 16'h3C3C;
    wire [15:0] _T_790;
    assign _T_790 = 16'h3333;
    wire [13:0] _T_791;
    SHR_UNSIGNED #(.width(16), .n(2)) u_shr_4372 (
        .y(_T_791),
        .in(_T_787)
    );
    wire [15:0] _T_792;
    wire [15:0] _WTEMP_602;
    PAD_UNSIGNED #(.width(14), .n(16)) u_pad_4373 (
        .y(_WTEMP_602),
        .in(_T_791)
    );
    BITWISEAND #(.width(16)) bitwiseand_4374 (
        .y(_T_792),
        .a(_WTEMP_602),
        .b(_T_790)
    );
    wire [13:0] _T_793;
    BITS #(.width(16), .high(13), .low(0)) bits_4375 (
        .y(_T_793),
        .in(_T_787)
    );
    wire [15:0] _T_794;
    SHL_UNSIGNED #(.width(14), .n(2)) u_shl_4376 (
        .y(_T_794),
        .in(_T_793)
    );
    wire [15:0] _T_795;
    assign _T_795 = 16'hCCCC;
    wire [15:0] _T_796;
    BITWISEAND #(.width(16)) bitwiseand_4377 (
        .y(_T_796),
        .a(_T_794),
        .b(_T_795)
    );
    wire [15:0] _T_797;
    BITWISEOR #(.width(16)) bitwiseor_4378 (
        .y(_T_797),
        .a(_T_792),
        .b(_T_796)
    );
    wire [14:0] _T_798;
    assign _T_798 = 15'h3333;
    wire [15:0] _T_799;
    assign _T_799 = 16'h6666;
    wire [15:0] _T_800;
    assign _T_800 = 16'h5555;
    wire [14:0] _T_801;
    SHR_UNSIGNED #(.width(16), .n(1)) u_shr_4379 (
        .y(_T_801),
        .in(_T_797)
    );
    wire [15:0] _T_802;
    wire [15:0] _WTEMP_603;
    PAD_UNSIGNED #(.width(15), .n(16)) u_pad_4380 (
        .y(_WTEMP_603),
        .in(_T_801)
    );
    BITWISEAND #(.width(16)) bitwiseand_4381 (
        .y(_T_802),
        .a(_WTEMP_603),
        .b(_T_800)
    );
    wire [14:0] _T_803;
    BITS #(.width(16), .high(14), .low(0)) bits_4382 (
        .y(_T_803),
        .in(_T_797)
    );
    wire [15:0] _T_804;
    SHL_UNSIGNED #(.width(15), .n(1)) u_shl_4383 (
        .y(_T_804),
        .in(_T_803)
    );
    wire [15:0] _T_805;
    assign _T_805 = 16'hAAAA;
    wire [15:0] _T_806;
    BITWISEAND #(.width(16)) bitwiseand_4384 (
        .y(_T_806),
        .a(_T_804),
        .b(_T_805)
    );
    wire [15:0] _T_807;
    BITWISEOR #(.width(16)) bitwiseor_4385 (
        .y(_T_807),
        .a(_T_802),
        .b(_T_806)
    );
    wire [1:0] _T_808;
    BITS #(.width(18), .high(17), .low(16)) bits_4386 (
        .y(_T_808),
        .in(_T_765)
    );
    wire _T_809;
    BITS #(.width(2), .high(0), .low(0)) bits_4387 (
        .y(_T_809),
        .in(_T_808)
    );
    wire _T_810;
    BITS #(.width(2), .high(1), .low(1)) bits_4388 (
        .y(_T_810),
        .in(_T_808)
    );
    wire [1:0] _T_811;
    CAT #(.width_a(1), .width_b(1)) cat_4389 (
        .y(_T_811),
        .a(_T_809),
        .b(_T_810)
    );
    wire [17:0] _T_812;
    CAT #(.width_a(16), .width_b(2)) cat_4390 (
        .y(_T_812),
        .a(_T_807),
        .b(_T_811)
    );
    wire [49:0] _T_813;
    CAT #(.width_a(32), .width_b(18)) cat_4391 (
        .y(_T_813),
        .a(_T_764),
        .b(_T_812)
    );
    wire [49:0] _T_814;
    BITWISENOT #(.width(50)) bitwisenot_4392 (
        .y(_T_814),
        .in(_T_813)
    );
    wire [49:0] _T_815;
    wire [49:0] _WTEMP_604;
    PAD_UNSIGNED #(.width(1), .n(50)) u_pad_4393 (
        .y(_WTEMP_604),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(50)) u_mux_4394 (
        .y(_T_815),
        .sel(_T_707),
        .a(_WTEMP_604),
        .b(_T_814)
    );
    wire [49:0] _T_816;
    BITWISENOT #(.width(50)) bitwisenot_4395 (
        .y(_T_816),
        .in(_T_815)
    );
    wire [49:0] _T_817;
    BITWISENOT #(.width(50)) bitwisenot_4396 (
        .y(_T_817),
        .in(_T_816)
    );
    wire [49:0] _T_818;
    wire [49:0] _WTEMP_605;
    PAD_UNSIGNED #(.width(1), .n(50)) u_pad_4397 (
        .y(_WTEMP_605),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(50)) u_mux_4398 (
        .y(_T_818),
        .sel(_T_704),
        .a(_WTEMP_605),
        .b(_T_817)
    );
    wire [49:0] _T_819;
    BITWISENOT #(.width(50)) bitwisenot_4399 (
        .y(_T_819),
        .in(_T_818)
    );
    wire [49:0] _T_820;
    BITWISENOT #(.width(50)) bitwisenot_4400 (
        .y(_T_820),
        .in(_T_819)
    );
    wire [49:0] _T_821;
    wire [49:0] _WTEMP_606;
    PAD_UNSIGNED #(.width(1), .n(50)) u_pad_4401 (
        .y(_WTEMP_606),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(50)) u_mux_4402 (
        .y(_T_821),
        .sel(_T_701),
        .a(_WTEMP_606),
        .b(_T_820)
    );
    wire [49:0] _T_822;
    BITWISENOT #(.width(50)) bitwisenot_4403 (
        .y(_T_822),
        .in(_T_821)
    );
    wire [49:0] _T_823;
    BITWISENOT #(.width(50)) bitwisenot_4404 (
        .y(_T_823),
        .in(_T_822)
    );
    wire [49:0] _T_824;
    wire [49:0] _WTEMP_607;
    PAD_UNSIGNED #(.width(1), .n(50)) u_pad_4405 (
        .y(_WTEMP_607),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(50)) u_mux_4406 (
        .y(_T_824),
        .sel(_T_698),
        .a(_WTEMP_607),
        .b(_T_823)
    );
    wire [49:0] _T_825;
    BITWISENOT #(.width(50)) bitwisenot_4407 (
        .y(_T_825),
        .in(_T_824)
    );
    wire [53:0] _T_827;
    CAT #(.width_a(50), .width_b(4)) cat_4408 (
        .y(_T_827),
        .a(_T_825),
        .b(4'hF)
    );
    wire _T_828;
    BITS #(.width(10), .high(9), .low(9)) bits_4409 (
        .y(_T_828),
        .in(_T_697)
    );
    wire [8:0] _T_829;
    BITS #(.width(10), .high(8), .low(0)) bits_4410 (
        .y(_T_829),
        .in(_T_697)
    );
    wire _T_830;
    BITS #(.width(9), .high(8), .low(8)) bits_4411 (
        .y(_T_830),
        .in(_T_829)
    );
    wire [7:0] _T_831;
    BITS #(.width(9), .high(7), .low(0)) bits_4412 (
        .y(_T_831),
        .in(_T_829)
    );
    wire _T_832;
    BITS #(.width(8), .high(7), .low(7)) bits_4413 (
        .y(_T_832),
        .in(_T_831)
    );
    wire [6:0] _T_833;
    BITS #(.width(8), .high(6), .low(0)) bits_4414 (
        .y(_T_833),
        .in(_T_831)
    );
    wire _T_834;
    BITS #(.width(7), .high(6), .low(6)) bits_4415 (
        .y(_T_834),
        .in(_T_833)
    );
    wire [5:0] _T_835;
    BITS #(.width(7), .high(5), .low(0)) bits_4416 (
        .y(_T_835),
        .in(_T_833)
    );
    wire [64:0] _T_837;
    DSHR_SIGNED #(.width_in(65), .width_n(6)) s_dshr_4417 (
        .y(_T_837),
        .in(-65'sh10000000000000000),
        .n(_T_835)
    );
    wire [3:0] _T_838;
    BITS #(.width(65), .high(3), .low(0)) bits_4418 (
        .y(_T_838),
        .in(_T_837)
    );
    wire [1:0] _T_839;
    BITS #(.width(4), .high(1), .low(0)) bits_4419 (
        .y(_T_839),
        .in(_T_838)
    );
    wire _T_840;
    BITS #(.width(2), .high(0), .low(0)) bits_4420 (
        .y(_T_840),
        .in(_T_839)
    );
    wire _T_841;
    BITS #(.width(2), .high(1), .low(1)) bits_4421 (
        .y(_T_841),
        .in(_T_839)
    );
    wire [1:0] _T_842;
    CAT #(.width_a(1), .width_b(1)) cat_4422 (
        .y(_T_842),
        .a(_T_840),
        .b(_T_841)
    );
    wire [1:0] _T_843;
    BITS #(.width(4), .high(3), .low(2)) bits_4423 (
        .y(_T_843),
        .in(_T_838)
    );
    wire _T_844;
    BITS #(.width(2), .high(0), .low(0)) bits_4424 (
        .y(_T_844),
        .in(_T_843)
    );
    wire _T_845;
    BITS #(.width(2), .high(1), .low(1)) bits_4425 (
        .y(_T_845),
        .in(_T_843)
    );
    wire [1:0] _T_846;
    CAT #(.width_a(1), .width_b(1)) cat_4426 (
        .y(_T_846),
        .a(_T_844),
        .b(_T_845)
    );
    wire [3:0] _T_847;
    CAT #(.width_a(2), .width_b(2)) cat_4427 (
        .y(_T_847),
        .a(_T_842),
        .b(_T_846)
    );
    wire [3:0] _T_849;
    wire [3:0] _WTEMP_608;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_4428 (
        .y(_WTEMP_608),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(4)) u_mux_4429 (
        .y(_T_849),
        .sel(_T_834),
        .a(_T_847),
        .b(_WTEMP_608)
    );
    wire [3:0] _T_851;
    wire [3:0] _WTEMP_609;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_4430 (
        .y(_WTEMP_609),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(4)) u_mux_4431 (
        .y(_T_851),
        .sel(_T_832),
        .a(_T_849),
        .b(_WTEMP_609)
    );
    wire [3:0] _T_853;
    wire [3:0] _WTEMP_610;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_4432 (
        .y(_WTEMP_610),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(4)) u_mux_4433 (
        .y(_T_853),
        .sel(_T_830),
        .a(_T_851),
        .b(_WTEMP_610)
    );
    wire [3:0] _T_855;
    wire [3:0] _WTEMP_611;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_4434 (
        .y(_WTEMP_611),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(4)) u_mux_4435 (
        .y(_T_855),
        .sel(_T_828),
        .a(_T_853),
        .b(_WTEMP_611)
    );
    wire [53:0] _T_856;
    wire [53:0] _WTEMP_612;
    PAD_UNSIGNED #(.width(4), .n(54)) u_pad_4436 (
        .y(_WTEMP_612),
        .in(_T_855)
    );
    MUX_UNSIGNED #(.width(54)) u_mux_4437 (
        .y(_T_856),
        .sel(_T_696),
        .a(_T_827),
        .b(_WTEMP_612)
    );
    wire [53:0] _T_858;
    wire [53:0] _WTEMP_613;
    PAD_UNSIGNED #(.width(1), .n(54)) u_pad_4438 (
        .y(_WTEMP_613),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(54)) u_mux_4439 (
        .y(_T_858),
        .sel(_T_694),
        .a(_T_856),
        .b(_WTEMP_613)
    );
    wire [53:0] _T_860;
    wire [53:0] _WTEMP_614;
    PAD_UNSIGNED #(.width(1), .n(54)) u_pad_4440 (
        .y(_WTEMP_614),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(54)) u_mux_4441 (
        .y(_T_860),
        .sel(_T_692),
        .a(_T_858),
        .b(_WTEMP_614)
    );
    wire _T_861;
    BITS #(.width(57), .high(55), .low(55)) bits_4442 (
        .y(_T_861),
        .in(sigX3)
    );
    wire [53:0] _T_862;
    wire [53:0] _WTEMP_615;
    PAD_UNSIGNED #(.width(1), .n(54)) u_pad_4443 (
        .y(_WTEMP_615),
        .in(_T_861)
    );
    BITWISEOR #(.width(54)) bitwiseor_4444 (
        .y(_T_862),
        .a(_T_860),
        .b(_WTEMP_615)
    );
    wire [55:0] _T_864;
    CAT #(.width_a(54), .width_b(2)) cat_4445 (
        .y(_T_864),
        .a(_T_862),
        .b(2'h3)
    );
    wire [55:0] roundMask;
    BITWISEOR #(.width(56)) bitwiseor_4446 (
        .y(roundMask),
        .a(_T_690),
        .b(_T_864)
    );
    wire [54:0] _T_865;
    SHR_UNSIGNED #(.width(56), .n(1)) u_shr_4447 (
        .y(_T_865),
        .in(roundMask)
    );
    wire [54:0] _T_866;
    BITWISENOT #(.width(55)) bitwisenot_4448 (
        .y(_T_866),
        .in(_T_865)
    );
    wire [55:0] roundPosMask;
    wire [55:0] _WTEMP_616;
    PAD_UNSIGNED #(.width(55), .n(56)) u_pad_4449 (
        .y(_WTEMP_616),
        .in(_T_866)
    );
    BITWISEAND #(.width(56)) bitwiseand_4450 (
        .y(roundPosMask),
        .a(_WTEMP_616),
        .b(roundMask)
    );
    wire [56:0] _T_867;
    wire [56:0] _WTEMP_617;
    PAD_UNSIGNED #(.width(56), .n(57)) u_pad_4451 (
        .y(_WTEMP_617),
        .in(roundPosMask)
    );
    BITWISEAND #(.width(57)) bitwiseand_4452 (
        .y(_T_867),
        .a(sigX3),
        .b(_WTEMP_617)
    );
    wire roundPosBit;
    wire [56:0] _WTEMP_618;
    PAD_UNSIGNED #(.width(1), .n(57)) u_pad_4453 (
        .y(_WTEMP_618),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(57)) u_neq_4454 (
        .y(roundPosBit),
        .a(_T_867),
        .b(_WTEMP_618)
    );
    wire [54:0] _T_869;
    SHR_UNSIGNED #(.width(56), .n(1)) u_shr_4455 (
        .y(_T_869),
        .in(roundMask)
    );
    wire [56:0] _T_870;
    wire [56:0] _WTEMP_619;
    PAD_UNSIGNED #(.width(55), .n(57)) u_pad_4456 (
        .y(_WTEMP_619),
        .in(_T_869)
    );
    BITWISEAND #(.width(57)) bitwiseand_4457 (
        .y(_T_870),
        .a(sigX3),
        .b(_WTEMP_619)
    );
    wire anyRoundExtra;
    wire [56:0] _WTEMP_620;
    PAD_UNSIGNED #(.width(1), .n(57)) u_pad_4458 (
        .y(_WTEMP_620),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(57)) u_neq_4459 (
        .y(anyRoundExtra),
        .a(_T_870),
        .b(_WTEMP_620)
    );
    wire [56:0] _T_872;
    BITWISENOT #(.width(57)) bitwisenot_4460 (
        .y(_T_872),
        .in(sigX3)
    );
    wire [54:0] _T_873;
    SHR_UNSIGNED #(.width(56), .n(1)) u_shr_4461 (
        .y(_T_873),
        .in(roundMask)
    );
    wire [56:0] _T_874;
    wire [56:0] _WTEMP_621;
    PAD_UNSIGNED #(.width(55), .n(57)) u_pad_4462 (
        .y(_WTEMP_621),
        .in(_T_873)
    );
    BITWISEAND #(.width(57)) bitwiseand_4463 (
        .y(_T_874),
        .a(_T_872),
        .b(_WTEMP_621)
    );
    wire allRoundExtra;
    wire [56:0] _WTEMP_622;
    PAD_UNSIGNED #(.width(1), .n(57)) u_pad_4464 (
        .y(_WTEMP_622),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(57)) u_eq_4465 (
        .y(allRoundExtra),
        .a(_T_874),
        .b(_WTEMP_622)
    );
    wire anyRound;
    BITWISEOR #(.width(1)) bitwiseor_4466 (
        .y(anyRound),
        .a(roundPosBit),
        .b(anyRoundExtra)
    );
    wire allRound;
    BITWISEAND #(.width(1)) bitwiseand_4467 (
        .y(allRound),
        .a(roundPosBit),
        .b(allRoundExtra)
    );
    wire roundDirectUp;
    MUX_UNSIGNED #(.width(1)) u_mux_4468 (
        .y(roundDirectUp),
        .sel(signY),
        .a(roundingMode_min),
        .b(roundingMode_max)
    );
    wire _T_877;
    EQ_UNSIGNED #(.width(1)) u_eq_4469 (
        .y(_T_877),
        .a(doIncrSig),
        .b(1'h0)
    );
    wire _T_878;
    BITWISEAND #(.width(1)) bitwiseand_4470 (
        .y(_T_878),
        .a(_T_877),
        .b(roundingMode_nearest_even)
    );
    wire _T_879;
    BITWISEAND #(.width(1)) bitwiseand_4471 (
        .y(_T_879),
        .a(_T_878),
        .b(roundPosBit)
    );
    wire _T_880;
    BITWISEAND #(.width(1)) bitwiseand_4472 (
        .y(_T_880),
        .a(_T_879),
        .b(anyRoundExtra)
    );
    wire _T_882;
    EQ_UNSIGNED #(.width(1)) u_eq_4473 (
        .y(_T_882),
        .a(doIncrSig),
        .b(1'h0)
    );
    wire _T_883;
    BITWISEAND #(.width(1)) bitwiseand_4474 (
        .y(_T_883),
        .a(_T_882),
        .b(roundDirectUp)
    );
    wire _T_884;
    BITWISEAND #(.width(1)) bitwiseand_4475 (
        .y(_T_884),
        .a(_T_883),
        .b(anyRound)
    );
    wire _T_885;
    BITWISEOR #(.width(1)) bitwiseor_4476 (
        .y(_T_885),
        .a(_T_880),
        .b(_T_884)
    );
    wire _T_886;
    BITWISEAND #(.width(1)) bitwiseand_4477 (
        .y(_T_886),
        .a(doIncrSig),
        .b(allRound)
    );
    wire _T_887;
    BITWISEOR #(.width(1)) bitwiseor_4478 (
        .y(_T_887),
        .a(_T_885),
        .b(_T_886)
    );
    wire _T_888;
    BITWISEAND #(.width(1)) bitwiseand_4479 (
        .y(_T_888),
        .a(doIncrSig),
        .b(roundingMode_nearest_even)
    );
    wire _T_889;
    BITWISEAND #(.width(1)) bitwiseand_4480 (
        .y(_T_889),
        .a(_T_888),
        .b(roundPosBit)
    );
    wire _T_890;
    BITWISEOR #(.width(1)) bitwiseor_4481 (
        .y(_T_890),
        .a(_T_887),
        .b(_T_889)
    );
    wire _T_891;
    BITWISEAND #(.width(1)) bitwiseand_4482 (
        .y(_T_891),
        .a(doIncrSig),
        .b(roundDirectUp)
    );
    wire _T_893;
    BITWISEAND #(.width(1)) bitwiseand_4483 (
        .y(_T_893),
        .a(_T_891),
        .b(1'h1)
    );
    wire roundUp;
    BITWISEOR #(.width(1)) bitwiseor_4484 (
        .y(roundUp),
        .a(_T_890),
        .b(_T_893)
    );
    wire _T_895;
    EQ_UNSIGNED #(.width(1)) u_eq_4485 (
        .y(_T_895),
        .a(roundPosBit),
        .b(1'h0)
    );
    wire _T_896;
    BITWISEAND #(.width(1)) bitwiseand_4486 (
        .y(_T_896),
        .a(roundingMode_nearest_even),
        .b(_T_895)
    );
    wire _T_897;
    BITWISEAND #(.width(1)) bitwiseand_4487 (
        .y(_T_897),
        .a(_T_896),
        .b(allRoundExtra)
    );
    wire _T_898;
    BITWISEAND #(.width(1)) bitwiseand_4488 (
        .y(_T_898),
        .a(roundingMode_nearest_even),
        .b(roundPosBit)
    );
    wire _T_900;
    EQ_UNSIGNED #(.width(1)) u_eq_4489 (
        .y(_T_900),
        .a(anyRoundExtra),
        .b(1'h0)
    );
    wire _T_901;
    BITWISEAND #(.width(1)) bitwiseand_4490 (
        .y(_T_901),
        .a(_T_898),
        .b(_T_900)
    );
    wire roundEven;
    MUX_UNSIGNED #(.width(1)) u_mux_4491 (
        .y(roundEven),
        .sel(doIncrSig),
        .a(_T_897),
        .b(_T_901)
    );
    wire _T_903;
    EQ_UNSIGNED #(.width(1)) u_eq_4492 (
        .y(_T_903),
        .a(allRound),
        .b(1'h0)
    );
    wire inexactY;
    MUX_UNSIGNED #(.width(1)) u_mux_4493 (
        .y(inexactY),
        .sel(doIncrSig),
        .a(_T_903),
        .b(anyRound)
    );
    wire [56:0] _T_904;
    wire [56:0] _WTEMP_623;
    PAD_UNSIGNED #(.width(56), .n(57)) u_pad_4494 (
        .y(_WTEMP_623),
        .in(roundMask)
    );
    BITWISEOR #(.width(57)) bitwiseor_4495 (
        .y(_T_904),
        .a(sigX3),
        .b(_WTEMP_623)
    );
    wire [54:0] _T_905;
    SHR_UNSIGNED #(.width(57), .n(2)) u_shr_4496 (
        .y(_T_905),
        .in(_T_904)
    );
    wire [55:0] _T_907;
    wire [54:0] _WTEMP_624;
    PAD_UNSIGNED #(.width(1), .n(55)) u_pad_4497 (
        .y(_WTEMP_624),
        .in(1'h1)
    );
    ADD_UNSIGNED #(.width(55)) u_add_4498 (
        .y(_T_907),
        .a(_T_905),
        .b(_WTEMP_624)
    );
    wire [54:0] _T_908;
    TAIL #(.width(56), .n(1)) tail_4499 (
        .y(_T_908),
        .in(_T_907)
    );
    wire [54:0] roundUp_sigY3;
    BITS #(.width(55), .high(54), .low(0)) bits_4500 (
        .y(roundUp_sigY3),
        .in(_T_908)
    );
    wire _T_910;
    EQ_UNSIGNED #(.width(1)) u_eq_4501 (
        .y(_T_910),
        .a(roundUp),
        .b(1'h0)
    );
    wire _T_912;
    EQ_UNSIGNED #(.width(1)) u_eq_4502 (
        .y(_T_912),
        .a(roundEven),
        .b(1'h0)
    );
    wire _T_913;
    BITWISEAND #(.width(1)) bitwiseand_4503 (
        .y(_T_913),
        .a(_T_910),
        .b(_T_912)
    );
    wire [55:0] _T_914;
    BITWISENOT #(.width(56)) bitwisenot_4504 (
        .y(_T_914),
        .in(roundMask)
    );
    wire [56:0] _T_915;
    wire [56:0] _WTEMP_625;
    PAD_UNSIGNED #(.width(56), .n(57)) u_pad_4505 (
        .y(_WTEMP_625),
        .in(_T_914)
    );
    BITWISEAND #(.width(57)) bitwiseand_4506 (
        .y(_T_915),
        .a(sigX3),
        .b(_WTEMP_625)
    );
    wire [54:0] _T_916;
    SHR_UNSIGNED #(.width(57), .n(2)) u_shr_4507 (
        .y(_T_916),
        .in(_T_915)
    );
    wire [54:0] _T_918;
    wire [54:0] _WTEMP_626;
    PAD_UNSIGNED #(.width(1), .n(55)) u_pad_4508 (
        .y(_WTEMP_626),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(55)) u_mux_4509 (
        .y(_T_918),
        .sel(_T_913),
        .a(_T_916),
        .b(_WTEMP_626)
    );
    wire [54:0] _T_920;
    wire [54:0] _WTEMP_627;
    PAD_UNSIGNED #(.width(1), .n(55)) u_pad_4510 (
        .y(_WTEMP_627),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(55)) u_mux_4511 (
        .y(_T_920),
        .sel(roundUp),
        .a(roundUp_sigY3),
        .b(_WTEMP_627)
    );
    wire [54:0] _T_921;
    BITWISEOR #(.width(55)) bitwiseor_4512 (
        .y(_T_921),
        .a(_T_918),
        .b(_T_920)
    );
    wire [54:0] _T_922;
    SHR_UNSIGNED #(.width(56), .n(1)) u_shr_4513 (
        .y(_T_922),
        .in(roundMask)
    );
    wire [54:0] _T_923;
    BITWISENOT #(.width(55)) bitwisenot_4514 (
        .y(_T_923),
        .in(_T_922)
    );
    wire [54:0] _T_924;
    BITWISEAND #(.width(55)) bitwiseand_4515 (
        .y(_T_924),
        .a(roundUp_sigY3),
        .b(_T_923)
    );
    wire [54:0] _T_926;
    wire [54:0] _WTEMP_628;
    PAD_UNSIGNED #(.width(1), .n(55)) u_pad_4516 (
        .y(_WTEMP_628),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(55)) u_mux_4517 (
        .y(_T_926),
        .sel(roundEven),
        .a(_T_924),
        .b(_WTEMP_628)
    );
    wire [54:0] sigY3;
    BITWISEOR #(.width(55)) bitwiseor_4518 (
        .y(sigY3),
        .a(_T_921),
        .b(_T_926)
    );
    wire _T_927;
    BITS #(.width(55), .high(54), .low(54)) bits_4519 (
        .y(_T_927),
        .in(sigY3)
    );
    wire [14:0] _T_929;
    wire [13:0] _WTEMP_629;
    PAD_UNSIGNED #(.width(1), .n(14)) u_pad_4520 (
        .y(_WTEMP_629),
        .in(1'h1)
    );
    ADD_UNSIGNED #(.width(14)) u_add_4521 (
        .y(_T_929),
        .a(sExpX3),
        .b(_WTEMP_629)
    );
    wire [13:0] _T_930;
    TAIL #(.width(15), .n(1)) tail_4522 (
        .y(_T_930),
        .in(_T_929)
    );
    wire [13:0] _T_932;
    wire [13:0] _WTEMP_630;
    PAD_UNSIGNED #(.width(1), .n(14)) u_pad_4523 (
        .y(_WTEMP_630),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(14)) u_mux_4524 (
        .y(_T_932),
        .sel(_T_927),
        .a(_T_930),
        .b(_WTEMP_630)
    );
    wire _T_933;
    BITS #(.width(55), .high(53), .low(53)) bits_4525 (
        .y(_T_933),
        .in(sigY3)
    );
    wire [13:0] _T_935;
    wire [13:0] _WTEMP_631;
    PAD_UNSIGNED #(.width(1), .n(14)) u_pad_4526 (
        .y(_WTEMP_631),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(14)) u_mux_4527 (
        .y(_T_935),
        .sel(_T_933),
        .a(sExpX3),
        .b(_WTEMP_631)
    );
    wire [13:0] _T_936;
    BITWISEOR #(.width(14)) bitwiseor_4528 (
        .y(_T_936),
        .a(_T_932),
        .b(_T_935)
    );
    wire [1:0] _T_937;
    BITS #(.width(55), .high(54), .low(53)) bits_4529 (
        .y(_T_937),
        .in(sigY3)
    );
    wire _T_939;
    wire [1:0] _WTEMP_632;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_4530 (
        .y(_WTEMP_632),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(2)) u_eq_4531 (
        .y(_T_939),
        .a(_T_937),
        .b(_WTEMP_632)
    );
    wire [14:0] _T_941;
    wire [13:0] _WTEMP_633;
    PAD_UNSIGNED #(.width(1), .n(14)) u_pad_4532 (
        .y(_WTEMP_633),
        .in(1'h1)
    );
    SUB_UNSIGNED #(.width(14)) u_sub_4533 (
        .y(_T_941),
        .a(sExpX3),
        .b(_WTEMP_633)
    );
    wire [14:0] _T_942;
    ASUINT #(.width(15)) asuint_4534 (
        .y(_T_942),
        .in(_T_941)
    );
    wire [13:0] _T_943;
    TAIL #(.width(15), .n(1)) tail_4535 (
        .y(_T_943),
        .in(_T_942)
    );
    wire [13:0] _T_945;
    wire [13:0] _WTEMP_634;
    PAD_UNSIGNED #(.width(1), .n(14)) u_pad_4536 (
        .y(_WTEMP_634),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(14)) u_mux_4537 (
        .y(_T_945),
        .sel(_T_939),
        .a(_T_943),
        .b(_WTEMP_634)
    );
    wire [13:0] sExpY;
    BITWISEOR #(.width(14)) bitwiseor_4538 (
        .y(sExpY),
        .a(_T_936),
        .b(_T_945)
    );
    wire [11:0] expY;
    BITS #(.width(14), .high(11), .low(0)) bits_4539 (
        .y(expY),
        .in(sExpY)
    );
    wire [51:0] _T_946;
    BITS #(.width(55), .high(51), .low(0)) bits_4540 (
        .y(_T_946),
        .in(sigY3)
    );
    wire [51:0] _T_947;
    BITS #(.width(55), .high(52), .low(1)) bits_4541 (
        .y(_T_947),
        .in(sigY3)
    );
    wire [51:0] fractY;
    MUX_UNSIGNED #(.width(52)) u_mux_4542 (
        .y(fractY),
        .sel(sigX3Shift1),
        .a(_T_946),
        .b(_T_947)
    );
    wire [2:0] _T_948;
    BITS #(.width(14), .high(12), .low(10)) bits_4543 (
        .y(_T_948),
        .in(sExpY)
    );
    wire overflowY;
    wire [2:0] _WTEMP_635;
    PAD_UNSIGNED #(.width(2), .n(3)) u_pad_4544 (
        .y(_WTEMP_635),
        .in(2'h3)
    );
    EQ_UNSIGNED #(.width(3)) u_eq_4545 (
        .y(overflowY),
        .a(_T_948),
        .b(_WTEMP_635)
    );
    wire _T_951;
    EQ_UNSIGNED #(.width(1)) u_eq_4546 (
        .y(_T_951),
        .a(isZeroY),
        .b(1'h0)
    );
    wire _T_952;
    BITS #(.width(14), .high(12), .low(12)) bits_4547 (
        .y(_T_952),
        .in(sExpY)
    );
    wire [11:0] _T_953;
    BITS #(.width(14), .high(11), .low(0)) bits_4548 (
        .y(_T_953),
        .in(sExpY)
    );
    wire _T_955;
    wire [11:0] _WTEMP_636;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_4549 (
        .y(_WTEMP_636),
        .in(10'h3CE)
    );
    LT_UNSIGNED #(.width(12)) u_lt_4550 (
        .y(_T_955),
        .a(_T_953),
        .b(_WTEMP_636)
    );
    wire _T_956;
    BITWISEOR #(.width(1)) bitwiseor_4551 (
        .y(_T_956),
        .a(_T_952),
        .b(_T_955)
    );
    wire totalUnderflowY;
    BITWISEAND #(.width(1)) bitwiseand_4552 (
        .y(totalUnderflowY),
        .a(_T_951),
        .b(_T_956)
    );
    wire _T_957;
    BITS #(.width(14), .high(13), .low(13)) bits_4553 (
        .y(_T_957),
        .in(sExpX3)
    );
    wire [10:0] _T_960;
    MUX_UNSIGNED #(.width(11)) u_mux_4554 (
        .y(_T_960),
        .sel(sigX3Shift1),
        .a(11'h402),
        .b(11'h401)
    );
    wire _T_961;
    wire [12:0] _WTEMP_637;
    PAD_UNSIGNED #(.width(11), .n(13)) u_pad_4555 (
        .y(_WTEMP_637),
        .in(_T_960)
    );
    LEQ_UNSIGNED #(.width(13)) u_leq_4556 (
        .y(_T_961),
        .a(sExpX3_13),
        .b(_WTEMP_637)
    );
    wire _T_962;
    BITWISEOR #(.width(1)) bitwiseor_4557 (
        .y(_T_962),
        .a(_T_957),
        .b(_T_961)
    );
    wire underflowY;
    BITWISEAND #(.width(1)) bitwiseand_4558 (
        .y(underflowY),
        .a(inexactY),
        .b(_T_962)
    );
    wire _T_963;
    BITWISEAND #(.width(1)) bitwiseand_4559 (
        .y(_T_963),
        .a(roundingMode_min),
        .b(signY)
    );
    wire _T_965;
    EQ_UNSIGNED #(.width(1)) u_eq_4560 (
        .y(_T_965),
        .a(signY),
        .b(1'h0)
    );
    wire _T_966;
    BITWISEAND #(.width(1)) bitwiseand_4561 (
        .y(_T_966),
        .a(roundingMode_max),
        .b(_T_965)
    );
    wire roundMagUp;
    BITWISEOR #(.width(1)) bitwiseor_4562 (
        .y(roundMagUp),
        .a(_T_963),
        .b(_T_966)
    );
    wire overflowY_roundMagUp;
    BITWISEOR #(.width(1)) bitwiseor_4563 (
        .y(overflowY_roundMagUp),
        .a(roundingMode_nearest_even),
        .b(roundMagUp)
    );
    wire mulSpecial;
    BITWISEOR #(.width(1)) bitwiseor_4564 (
        .y(mulSpecial),
        .a(isSpecialA),
        .b(isSpecialB)
    );
    wire addSpecial;
    BITWISEOR #(.width(1)) bitwiseor_4565 (
        .y(addSpecial),
        .a(mulSpecial),
        .b(isSpecialC)
    );
    wire notSpecial_addZeros;
    BITWISEAND #(.width(1)) bitwiseand_4566 (
        .y(notSpecial_addZeros),
        .a(io_fromPreMul_isZeroProd),
        .b(isZeroC)
    );
    wire _T_968;
    EQ_UNSIGNED #(.width(1)) u_eq_4567 (
        .y(_T_968),
        .a(addSpecial),
        .b(1'h0)
    );
    wire _T_970;
    EQ_UNSIGNED #(.width(1)) u_eq_4568 (
        .y(_T_970),
        .a(notSpecial_addZeros),
        .b(1'h0)
    );
    wire commonCase;
    BITWISEAND #(.width(1)) bitwiseand_4569 (
        .y(commonCase),
        .a(_T_968),
        .b(_T_970)
    );
    wire _T_971;
    BITWISEAND #(.width(1)) bitwiseand_4570 (
        .y(_T_971),
        .a(isInfA),
        .b(isZeroB)
    );
    wire _T_972;
    BITWISEAND #(.width(1)) bitwiseand_4571 (
        .y(_T_972),
        .a(isZeroA),
        .b(isInfB)
    );
    wire _T_973;
    BITWISEOR #(.width(1)) bitwiseor_4572 (
        .y(_T_973),
        .a(_T_971),
        .b(_T_972)
    );
    wire _T_975;
    EQ_UNSIGNED #(.width(1)) u_eq_4573 (
        .y(_T_975),
        .a(isNaNA),
        .b(1'h0)
    );
    wire _T_977;
    EQ_UNSIGNED #(.width(1)) u_eq_4574 (
        .y(_T_977),
        .a(isNaNB),
        .b(1'h0)
    );
    wire _T_978;
    BITWISEAND #(.width(1)) bitwiseand_4575 (
        .y(_T_978),
        .a(_T_975),
        .b(_T_977)
    );
    wire _T_979;
    BITWISEOR #(.width(1)) bitwiseor_4576 (
        .y(_T_979),
        .a(isInfA),
        .b(isInfB)
    );
    wire _T_980;
    BITWISEAND #(.width(1)) bitwiseand_4577 (
        .y(_T_980),
        .a(_T_978),
        .b(_T_979)
    );
    wire _T_981;
    BITWISEAND #(.width(1)) bitwiseand_4578 (
        .y(_T_981),
        .a(_T_980),
        .b(isInfC)
    );
    wire _T_982;
    BITWISEAND #(.width(1)) bitwiseand_4579 (
        .y(_T_982),
        .a(_T_981),
        .b(doSubMags)
    );
    wire notSigNaN_invalid;
    BITWISEOR #(.width(1)) bitwiseor_4580 (
        .y(notSigNaN_invalid),
        .a(_T_973),
        .b(_T_982)
    );
    wire _T_983;
    BITWISEOR #(.width(1)) bitwiseor_4581 (
        .y(_T_983),
        .a(isSigNaNA),
        .b(isSigNaNB)
    );
    wire _T_984;
    BITWISEOR #(.width(1)) bitwiseor_4582 (
        .y(_T_984),
        .a(_T_983),
        .b(isSigNaNC)
    );
    wire invalid;
    BITWISEOR #(.width(1)) bitwiseor_4583 (
        .y(invalid),
        .a(_T_984),
        .b(notSigNaN_invalid)
    );
    wire overflow;
    BITWISEAND #(.width(1)) bitwiseand_4584 (
        .y(overflow),
        .a(commonCase),
        .b(overflowY)
    );
    wire underflow;
    BITWISEAND #(.width(1)) bitwiseand_4585 (
        .y(underflow),
        .a(commonCase),
        .b(underflowY)
    );
    wire _T_985;
    BITWISEAND #(.width(1)) bitwiseand_4586 (
        .y(_T_985),
        .a(commonCase),
        .b(inexactY)
    );
    wire inexact;
    BITWISEOR #(.width(1)) bitwiseor_4587 (
        .y(inexact),
        .a(overflow),
        .b(_T_985)
    );
    wire _T_986;
    BITWISEOR #(.width(1)) bitwiseor_4588 (
        .y(_T_986),
        .a(notSpecial_addZeros),
        .b(isZeroY)
    );
    wire notSpecial_isZeroOut;
    BITWISEOR #(.width(1)) bitwiseor_4589 (
        .y(notSpecial_isZeroOut),
        .a(_T_986),
        .b(totalUnderflowY)
    );
    wire _T_987;
    BITWISEAND #(.width(1)) bitwiseand_4590 (
        .y(_T_987),
        .a(commonCase),
        .b(totalUnderflowY)
    );
    wire pegMinFiniteMagOut;
    BITWISEAND #(.width(1)) bitwiseand_4591 (
        .y(pegMinFiniteMagOut),
        .a(_T_987),
        .b(roundMagUp)
    );
    wire _T_989;
    EQ_UNSIGNED #(.width(1)) u_eq_4592 (
        .y(_T_989),
        .a(overflowY_roundMagUp),
        .b(1'h0)
    );
    wire pegMaxFiniteMagOut;
    BITWISEAND #(.width(1)) bitwiseand_4593 (
        .y(pegMaxFiniteMagOut),
        .a(overflow),
        .b(_T_989)
    );
    wire _T_990;
    BITWISEOR #(.width(1)) bitwiseor_4594 (
        .y(_T_990),
        .a(isInfA),
        .b(isInfB)
    );
    wire _T_991;
    BITWISEOR #(.width(1)) bitwiseor_4595 (
        .y(_T_991),
        .a(_T_990),
        .b(isInfC)
    );
    wire _T_992;
    BITWISEAND #(.width(1)) bitwiseand_4596 (
        .y(_T_992),
        .a(overflow),
        .b(overflowY_roundMagUp)
    );
    wire notNaN_isInfOut;
    BITWISEOR #(.width(1)) bitwiseor_4597 (
        .y(notNaN_isInfOut),
        .a(_T_991),
        .b(_T_992)
    );
    wire _T_993;
    BITWISEOR #(.width(1)) bitwiseor_4598 (
        .y(_T_993),
        .a(isNaNA),
        .b(isNaNB)
    );
    wire _T_994;
    BITWISEOR #(.width(1)) bitwiseor_4599 (
        .y(_T_994),
        .a(_T_993),
        .b(isNaNC)
    );
    wire isNaNOut;
    BITWISEOR #(.width(1)) bitwiseor_4600 (
        .y(isNaNOut),
        .a(_T_994),
        .b(notSigNaN_invalid)
    );
    wire _T_996;
    EQ_UNSIGNED #(.width(1)) u_eq_4601 (
        .y(_T_996),
        .a(doSubMags),
        .b(1'h0)
    );
    wire _T_997;
    BITWISEAND #(.width(1)) bitwiseand_4602 (
        .y(_T_997),
        .a(_T_996),
        .b(io_fromPreMul_opSignC)
    );
    wire _T_999;
    EQ_UNSIGNED #(.width(1)) u_eq_4603 (
        .y(_T_999),
        .a(isSpecialC),
        .b(1'h0)
    );
    wire _T_1000;
    BITWISEAND #(.width(1)) bitwiseand_4604 (
        .y(_T_1000),
        .a(mulSpecial),
        .b(_T_999)
    );
    wire _T_1001;
    BITWISEAND #(.width(1)) bitwiseand_4605 (
        .y(_T_1001),
        .a(_T_1000),
        .b(io_fromPreMul_signProd)
    );
    wire _T_1002;
    BITWISEOR #(.width(1)) bitwiseor_4606 (
        .y(_T_1002),
        .a(_T_997),
        .b(_T_1001)
    );
    wire _T_1004;
    EQ_UNSIGNED #(.width(1)) u_eq_4607 (
        .y(_T_1004),
        .a(mulSpecial),
        .b(1'h0)
    );
    wire _T_1005;
    BITWISEAND #(.width(1)) bitwiseand_4608 (
        .y(_T_1005),
        .a(_T_1004),
        .b(isSpecialC)
    );
    wire _T_1006;
    BITWISEAND #(.width(1)) bitwiseand_4609 (
        .y(_T_1006),
        .a(_T_1005),
        .b(io_fromPreMul_opSignC)
    );
    wire _T_1007;
    BITWISEOR #(.width(1)) bitwiseor_4610 (
        .y(_T_1007),
        .a(_T_1002),
        .b(_T_1006)
    );
    wire _T_1009;
    EQ_UNSIGNED #(.width(1)) u_eq_4611 (
        .y(_T_1009),
        .a(mulSpecial),
        .b(1'h0)
    );
    wire _T_1010;
    BITWISEAND #(.width(1)) bitwiseand_4612 (
        .y(_T_1010),
        .a(_T_1009),
        .b(notSpecial_addZeros)
    );
    wire _T_1011;
    BITWISEAND #(.width(1)) bitwiseand_4613 (
        .y(_T_1011),
        .a(_T_1010),
        .b(doSubMags)
    );
    wire _T_1012;
    BITWISEAND #(.width(1)) bitwiseand_4614 (
        .y(_T_1012),
        .a(_T_1011),
        .b(signZeroNotEqOpSigns)
    );
    wire uncommonCaseSignOut;
    BITWISEOR #(.width(1)) bitwiseor_4615 (
        .y(uncommonCaseSignOut),
        .a(_T_1007),
        .b(_T_1012)
    );
    wire _T_1014;
    EQ_UNSIGNED #(.width(1)) u_eq_4616 (
        .y(_T_1014),
        .a(isNaNOut),
        .b(1'h0)
    );
    wire _T_1015;
    BITWISEAND #(.width(1)) bitwiseand_4617 (
        .y(_T_1015),
        .a(_T_1014),
        .b(uncommonCaseSignOut)
    );
    wire _T_1016;
    BITWISEAND #(.width(1)) bitwiseand_4618 (
        .y(_T_1016),
        .a(commonCase),
        .b(signY)
    );
    wire signOut;
    BITWISEOR #(.width(1)) bitwiseor_4619 (
        .y(signOut),
        .a(_T_1015),
        .b(_T_1016)
    );
    wire [11:0] _T_1019;
    MUX_UNSIGNED #(.width(12)) u_mux_4620 (
        .y(_T_1019),
        .sel(notSpecial_isZeroOut),
        .a(12'hE00),
        .b(12'h0)
    );
    wire [11:0] _T_1020;
    BITWISENOT #(.width(12)) bitwisenot_4621 (
        .y(_T_1020),
        .in(_T_1019)
    );
    wire [11:0] _T_1021;
    BITWISEAND #(.width(12)) bitwiseand_4622 (
        .y(_T_1021),
        .a(expY),
        .b(_T_1020)
    );
    wire [11:0] _T_1023;
    assign _T_1023 = 12'hC31;
    wire [11:0] _T_1025;
    MUX_UNSIGNED #(.width(12)) u_mux_4623 (
        .y(_T_1025),
        .sel(pegMinFiniteMagOut),
        .a(_T_1023),
        .b(12'h0)
    );
    wire [11:0] _T_1026;
    BITWISENOT #(.width(12)) bitwisenot_4624 (
        .y(_T_1026),
        .in(_T_1025)
    );
    wire [11:0] _T_1027;
    BITWISEAND #(.width(12)) bitwiseand_4625 (
        .y(_T_1027),
        .a(_T_1021),
        .b(_T_1026)
    );
    wire [11:0] _T_1030;
    MUX_UNSIGNED #(.width(12)) u_mux_4626 (
        .y(_T_1030),
        .sel(pegMaxFiniteMagOut),
        .a(12'h400),
        .b(12'h0)
    );
    wire [11:0] _T_1031;
    BITWISENOT #(.width(12)) bitwisenot_4627 (
        .y(_T_1031),
        .in(_T_1030)
    );
    wire [11:0] _T_1032;
    BITWISEAND #(.width(12)) bitwiseand_4628 (
        .y(_T_1032),
        .a(_T_1027),
        .b(_T_1031)
    );
    wire [11:0] _T_1035;
    wire [11:0] _WTEMP_638;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_4629 (
        .y(_WTEMP_638),
        .in(10'h200)
    );
    MUX_UNSIGNED #(.width(12)) u_mux_4630 (
        .y(_T_1035),
        .sel(notNaN_isInfOut),
        .a(_WTEMP_638),
        .b(12'h0)
    );
    wire [11:0] _T_1036;
    BITWISENOT #(.width(12)) bitwisenot_4631 (
        .y(_T_1036),
        .in(_T_1035)
    );
    wire [11:0] _T_1037;
    BITWISEAND #(.width(12)) bitwiseand_4632 (
        .y(_T_1037),
        .a(_T_1032),
        .b(_T_1036)
    );
    wire [11:0] _T_1040;
    wire [11:0] _WTEMP_639;
    PAD_UNSIGNED #(.width(10), .n(12)) u_pad_4633 (
        .y(_WTEMP_639),
        .in(10'h3CE)
    );
    MUX_UNSIGNED #(.width(12)) u_mux_4634 (
        .y(_T_1040),
        .sel(pegMinFiniteMagOut),
        .a(_WTEMP_639),
        .b(12'h0)
    );
    wire [11:0] _T_1041;
    BITWISEOR #(.width(12)) bitwiseor_4635 (
        .y(_T_1041),
        .a(_T_1037),
        .b(_T_1040)
    );
    wire [11:0] _T_1044;
    MUX_UNSIGNED #(.width(12)) u_mux_4636 (
        .y(_T_1044),
        .sel(pegMaxFiniteMagOut),
        .a(12'hBFF),
        .b(12'h0)
    );
    wire [11:0] _T_1045;
    BITWISEOR #(.width(12)) bitwiseor_4637 (
        .y(_T_1045),
        .a(_T_1041),
        .b(_T_1044)
    );
    wire [11:0] _T_1048;
    MUX_UNSIGNED #(.width(12)) u_mux_4638 (
        .y(_T_1048),
        .sel(notNaN_isInfOut),
        .a(12'hC00),
        .b(12'h0)
    );
    wire [11:0] _T_1049;
    BITWISEOR #(.width(12)) bitwiseor_4639 (
        .y(_T_1049),
        .a(_T_1045),
        .b(_T_1048)
    );
    wire [11:0] _T_1052;
    MUX_UNSIGNED #(.width(12)) u_mux_4640 (
        .y(_T_1052),
        .sel(isNaNOut),
        .a(12'hE00),
        .b(12'h0)
    );
    wire [11:0] expOut;
    BITWISEOR #(.width(12)) bitwiseor_4641 (
        .y(expOut),
        .a(_T_1049),
        .b(_T_1052)
    );
    wire _T_1053;
    BITWISEAND #(.width(1)) bitwiseand_4642 (
        .y(_T_1053),
        .a(totalUnderflowY),
        .b(roundMagUp)
    );
    wire _T_1054;
    BITWISEOR #(.width(1)) bitwiseor_4643 (
        .y(_T_1054),
        .a(_T_1053),
        .b(isNaNOut)
    );
    wire [51:0] _T_1056;
    assign _T_1056 = 52'h8000000000000;
    wire [51:0] _T_1058;
    wire [51:0] _WTEMP_640;
    PAD_UNSIGNED #(.width(1), .n(52)) u_pad_4644 (
        .y(_WTEMP_640),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(52)) u_mux_4645 (
        .y(_T_1058),
        .sel(isNaNOut),
        .a(_T_1056),
        .b(_WTEMP_640)
    );
    wire [51:0] _T_1059;
    MUX_UNSIGNED #(.width(52)) u_mux_4646 (
        .y(_T_1059),
        .sel(_T_1054),
        .a(_T_1058),
        .b(fractY)
    );
    wire _T_1060;
    BITS #(.width(1), .high(0), .low(0)) bits_4647 (
        .y(_T_1060),
        .in(pegMaxFiniteMagOut)
    );
    wire [51:0] _T_1063;
    MUX_UNSIGNED #(.width(52)) u_mux_4648 (
        .y(_T_1063),
        .sel(_T_1060),
        .a(52'hFFFFFFFFFFFFF),
        .b(52'h0)
    );
    wire [51:0] fractOut;
    BITWISEOR #(.width(52)) bitwiseor_4649 (
        .y(fractOut),
        .a(_T_1059),
        .b(_T_1063)
    );
    wire [12:0] _T_1064;
    CAT #(.width_a(1), .width_b(12)) cat_4650 (
        .y(_T_1064),
        .a(signOut),
        .b(expOut)
    );
    wire [64:0] _T_1065;
    CAT #(.width_a(13), .width_b(52)) cat_4651 (
        .y(_T_1065),
        .a(_T_1064),
        .b(fractOut)
    );
    wire [1:0] _T_1067;
    CAT #(.width_a(1), .width_b(1)) cat_4652 (
        .y(_T_1067),
        .a(underflow),
        .b(inexact)
    );
    wire [1:0] _T_1068;
    CAT #(.width_a(1), .width_b(1)) cat_4653 (
        .y(_T_1068),
        .a(invalid),
        .b(1'h0)
    );
    wire [2:0] _T_1069;
    CAT #(.width_a(2), .width_b(1)) cat_4654 (
        .y(_T_1069),
        .a(_T_1068),
        .b(overflow)
    );
    wire [4:0] _T_1070;
    CAT #(.width_a(3), .width_b(2)) cat_4655 (
        .y(_T_1070),
        .a(_T_1069),
        .b(_T_1067)
    );
    assign io_exceptionFlags = _T_1070;
    assign io_out = _T_1065;
endmodule //MulAddRecFN_postMul_1
module DivSqrtRecF64(
    input clock,
    input reset,
    output io_inReady_div,
    output io_inReady_sqrt,
    input io_inValid,
    input io_sqrtOp,
    input [64:0] io_a,
    input [64:0] io_b,
    input [1:0] io_roundingMode,
    output io_outValid_div,
    output io_outValid_sqrt,
    output [64:0] io_out,
    output [4:0] io_exceptionFlags
);
    wire _ds__clock;
    wire _ds__reset;
    wire _ds__io_inReady_div;
    wire _ds__io_inReady_sqrt;
    wire _ds__io_inValid;
    wire _ds__io_sqrtOp;
    wire [64:0] _ds__io_a;
    wire [64:0] _ds__io_b;
    wire [1:0] _ds__io_roundingMode;
    wire _ds__io_outValid_div;
    wire _ds__io_outValid_sqrt;
    wire [64:0] _ds__io_out;
    wire [4:0] _ds__io_exceptionFlags;
    wire [3:0] _ds__io_usingMulAdd;
    wire _ds__io_latchMulAddA_0;
    wire [53:0] _ds__io_mulAddA_0;
    wire _ds__io_latchMulAddB_0;
    wire [53:0] _ds__io_mulAddB_0;
    wire [104:0] _ds__io_mulAddC_2;
    wire [104:0] _ds__io_mulAddResult_3;
    DivSqrtRecF64_mulAddZ31 ds (
        .clock(_ds__clock),
        .reset(_ds__reset),
        .io_inReady_div(_ds__io_inReady_div),
        .io_inReady_sqrt(_ds__io_inReady_sqrt),
        .io_inValid(_ds__io_inValid),
        .io_sqrtOp(_ds__io_sqrtOp),
        .io_a(_ds__io_a),
        .io_b(_ds__io_b),
        .io_roundingMode(_ds__io_roundingMode),
        .io_outValid_div(_ds__io_outValid_div),
        .io_outValid_sqrt(_ds__io_outValid_sqrt),
        .io_out(_ds__io_out),
        .io_exceptionFlags(_ds__io_exceptionFlags),
        .io_usingMulAdd(_ds__io_usingMulAdd),
        .io_latchMulAddA_0(_ds__io_latchMulAddA_0),
        .io_mulAddA_0(_ds__io_mulAddA_0),
        .io_latchMulAddB_0(_ds__io_latchMulAddB_0),
        .io_mulAddB_0(_ds__io_mulAddB_0),
        .io_mulAddC_2(_ds__io_mulAddC_2),
        .io_mulAddResult_3(_ds__io_mulAddResult_3)
    );
    wire _mul__clock;
    wire _mul__reset;
    wire _mul__io_val_s0;
    wire _mul__io_latch_a_s0;
    wire [53:0] _mul__io_a_s0;
    wire _mul__io_latch_b_s0;
    wire [53:0] _mul__io_b_s0;
    wire [104:0] _mul__io_c_s2;
    wire [104:0] _mul__io_result_s3;
    Mul54 mul (
        .clock(_mul__clock),
        .reset(_mul__reset),
        .io_val_s0(_mul__io_val_s0),
        .io_latch_a_s0(_mul__io_latch_a_s0),
        .io_a_s0(_mul__io_a_s0),
        .io_latch_b_s0(_mul__io_latch_b_s0),
        .io_b_s0(_mul__io_b_s0),
        .io_c_s2(_mul__io_c_s2),
        .io_result_s3(_mul__io_result_s3)
    );
    wire _T_24;
    BITS #(.width(4), .high(0), .low(0)) bits_6279 (
        .y(_T_24),
        .in(_ds__io_usingMulAdd)
    );
    assign _ds__clock = clock;
    assign _ds__io_a = io_a;
    assign _ds__io_b = io_b;
    assign _ds__io_inValid = io_inValid;
    assign _ds__io_mulAddResult_3 = _mul__io_result_s3;
    assign _ds__io_roundingMode = io_roundingMode;
    assign _ds__io_sqrtOp = io_sqrtOp;
    assign _ds__reset = reset;
    assign io_exceptionFlags = _ds__io_exceptionFlags;
    assign io_inReady_div = _ds__io_inReady_div;
    assign io_inReady_sqrt = _ds__io_inReady_sqrt;
    assign io_out = _ds__io_out;
    assign io_outValid_div = _ds__io_outValid_div;
    assign io_outValid_sqrt = _ds__io_outValid_sqrt;
    assign _mul__clock = clock;
    assign _mul__io_a_s0 = _ds__io_mulAddA_0;
    assign _mul__io_b_s0 = _ds__io_mulAddB_0;
    assign _mul__io_c_s2 = _ds__io_mulAddC_2;
    assign _mul__io_latch_a_s0 = _ds__io_latchMulAddA_0;
    assign _mul__io_latch_b_s0 = _ds__io_latchMulAddB_0;
    assign _mul__io_val_s0 = _T_24;
    assign _mul__reset = reset;
endmodule //DivSqrtRecF64
module DivSqrtRecF64_mulAddZ31(
    input clock,
    input reset,
    output io_inReady_div,
    output io_inReady_sqrt,
    input io_inValid,
    input io_sqrtOp,
    input [64:0] io_a,
    input [64:0] io_b,
    input [1:0] io_roundingMode,
    output io_outValid_div,
    output io_outValid_sqrt,
    output [64:0] io_out,
    output [4:0] io_exceptionFlags,
    output [3:0] io_usingMulAdd,
    output io_latchMulAddA_0,
    output [53:0] io_mulAddA_0,
    output io_latchMulAddB_0,
    output [53:0] io_mulAddB_0,
    output [104:0] io_mulAddC_2,
    input [104:0] io_mulAddResult_3
);
    wire _valid_PA__q;
    wire _valid_PA__d;
    DFF_POSCLK #(.width(1)) valid_PA (
        .q(_valid_PA__q),
        .d(_valid_PA__d),
        .clk(clock)
    );
    wire _WTEMP_691;
    MUX_UNSIGNED #(.width(1)) u_mux_4932 (
        .y(_valid_PA__d),
        .sel(reset),
        .a(1'h0),
        .b(_WTEMP_691)
    );
    wire _sqrtOp_PA__q;
    wire _sqrtOp_PA__d;
    DFF_POSCLK #(.width(1)) sqrtOp_PA (
        .q(_sqrtOp_PA__q),
        .d(_sqrtOp_PA__d),
        .clk(clock)
    );
    wire _sign_PA__q;
    wire _sign_PA__d;
    DFF_POSCLK #(.width(1)) sign_PA (
        .q(_sign_PA__q),
        .d(_sign_PA__d),
        .clk(clock)
    );
    wire [2:0] _specialCodeB_PA__q;
    wire [2:0] _specialCodeB_PA__d;
    DFF_POSCLK #(.width(3)) specialCodeB_PA (
        .q(_specialCodeB_PA__q),
        .d(_specialCodeB_PA__d),
        .clk(clock)
    );
    wire _fractB_51_PA__q;
    wire _fractB_51_PA__d;
    DFF_POSCLK #(.width(1)) fractB_51_PA (
        .q(_fractB_51_PA__q),
        .d(_fractB_51_PA__d),
        .clk(clock)
    );
    wire [1:0] _roundingMode_PA__q;
    wire [1:0] _roundingMode_PA__d;
    DFF_POSCLK #(.width(2)) roundingMode_PA (
        .q(_roundingMode_PA__q),
        .d(_roundingMode_PA__d),
        .clk(clock)
    );
    wire [2:0] _specialCodeA_PA__q;
    wire [2:0] _specialCodeA_PA__d;
    DFF_POSCLK #(.width(3)) specialCodeA_PA (
        .q(_specialCodeA_PA__q),
        .d(_specialCodeA_PA__d),
        .clk(clock)
    );
    wire _fractA_51_PA__q;
    wire _fractA_51_PA__d;
    DFF_POSCLK #(.width(1)) fractA_51_PA (
        .q(_fractA_51_PA__q),
        .d(_fractA_51_PA__d),
        .clk(clock)
    );
    wire [13:0] _exp_PA__q;
    wire [13:0] _exp_PA__d;
    DFF_POSCLK #(.width(14)) exp_PA (
        .q(_exp_PA__q),
        .d(_exp_PA__d),
        .clk(clock)
    );
    wire [50:0] _fractB_other_PA__q;
    wire [50:0] _fractB_other_PA__d;
    DFF_POSCLK #(.width(51)) fractB_other_PA (
        .q(_fractB_other_PA__q),
        .d(_fractB_other_PA__d),
        .clk(clock)
    );
    wire [50:0] _fractA_other_PA__q;
    wire [50:0] _fractA_other_PA__d;
    DFF_POSCLK #(.width(51)) fractA_other_PA (
        .q(_fractA_other_PA__q),
        .d(_fractA_other_PA__d),
        .clk(clock)
    );
    wire _valid_PB__q;
    wire _valid_PB__d;
    DFF_POSCLK #(.width(1)) valid_PB (
        .q(_valid_PB__q),
        .d(_valid_PB__d),
        .clk(clock)
    );
    wire _WTEMP_692;
    MUX_UNSIGNED #(.width(1)) u_mux_4933 (
        .y(_valid_PB__d),
        .sel(reset),
        .a(1'h0),
        .b(_WTEMP_692)
    );
    wire _sqrtOp_PB__q;
    wire _sqrtOp_PB__d;
    DFF_POSCLK #(.width(1)) sqrtOp_PB (
        .q(_sqrtOp_PB__q),
        .d(_sqrtOp_PB__d),
        .clk(clock)
    );
    wire _sign_PB__q;
    wire _sign_PB__d;
    DFF_POSCLK #(.width(1)) sign_PB (
        .q(_sign_PB__q),
        .d(_sign_PB__d),
        .clk(clock)
    );
    wire [2:0] _specialCodeA_PB__q;
    wire [2:0] _specialCodeA_PB__d;
    DFF_POSCLK #(.width(3)) specialCodeA_PB (
        .q(_specialCodeA_PB__q),
        .d(_specialCodeA_PB__d),
        .clk(clock)
    );
    wire _fractA_51_PB__q;
    wire _fractA_51_PB__d;
    DFF_POSCLK #(.width(1)) fractA_51_PB (
        .q(_fractA_51_PB__q),
        .d(_fractA_51_PB__d),
        .clk(clock)
    );
    wire [2:0] _specialCodeB_PB__q;
    wire [2:0] _specialCodeB_PB__d;
    DFF_POSCLK #(.width(3)) specialCodeB_PB (
        .q(_specialCodeB_PB__q),
        .d(_specialCodeB_PB__d),
        .clk(clock)
    );
    wire _fractB_51_PB__q;
    wire _fractB_51_PB__d;
    DFF_POSCLK #(.width(1)) fractB_51_PB (
        .q(_fractB_51_PB__q),
        .d(_fractB_51_PB__d),
        .clk(clock)
    );
    wire [1:0] _roundingMode_PB__q;
    wire [1:0] _roundingMode_PB__d;
    DFF_POSCLK #(.width(2)) roundingMode_PB (
        .q(_roundingMode_PB__q),
        .d(_roundingMode_PB__d),
        .clk(clock)
    );
    wire [13:0] _exp_PB__q;
    wire [13:0] _exp_PB__d;
    DFF_POSCLK #(.width(14)) exp_PB (
        .q(_exp_PB__q),
        .d(_exp_PB__d),
        .clk(clock)
    );
    wire _fractA_0_PB__q;
    wire _fractA_0_PB__d;
    DFF_POSCLK #(.width(1)) fractA_0_PB (
        .q(_fractA_0_PB__q),
        .d(_fractA_0_PB__d),
        .clk(clock)
    );
    wire [50:0] _fractB_other_PB__q;
    wire [50:0] _fractB_other_PB__d;
    DFF_POSCLK #(.width(51)) fractB_other_PB (
        .q(_fractB_other_PB__q),
        .d(_fractB_other_PB__d),
        .clk(clock)
    );
    wire _valid_PC__q;
    wire _valid_PC__d;
    DFF_POSCLK #(.width(1)) valid_PC (
        .q(_valid_PC__q),
        .d(_valid_PC__d),
        .clk(clock)
    );
    wire _WTEMP_693;
    MUX_UNSIGNED #(.width(1)) u_mux_4934 (
        .y(_valid_PC__d),
        .sel(reset),
        .a(1'h0),
        .b(_WTEMP_693)
    );
    wire _sqrtOp_PC__q;
    wire _sqrtOp_PC__d;
    DFF_POSCLK #(.width(1)) sqrtOp_PC (
        .q(_sqrtOp_PC__q),
        .d(_sqrtOp_PC__d),
        .clk(clock)
    );
    wire _sign_PC__q;
    wire _sign_PC__d;
    DFF_POSCLK #(.width(1)) sign_PC (
        .q(_sign_PC__q),
        .d(_sign_PC__d),
        .clk(clock)
    );
    wire [2:0] _specialCodeA_PC__q;
    wire [2:0] _specialCodeA_PC__d;
    DFF_POSCLK #(.width(3)) specialCodeA_PC (
        .q(_specialCodeA_PC__q),
        .d(_specialCodeA_PC__d),
        .clk(clock)
    );
    wire _fractA_51_PC__q;
    wire _fractA_51_PC__d;
    DFF_POSCLK #(.width(1)) fractA_51_PC (
        .q(_fractA_51_PC__q),
        .d(_fractA_51_PC__d),
        .clk(clock)
    );
    wire [2:0] _specialCodeB_PC__q;
    wire [2:0] _specialCodeB_PC__d;
    DFF_POSCLK #(.width(3)) specialCodeB_PC (
        .q(_specialCodeB_PC__q),
        .d(_specialCodeB_PC__d),
        .clk(clock)
    );
    wire _fractB_51_PC__q;
    wire _fractB_51_PC__d;
    DFF_POSCLK #(.width(1)) fractB_51_PC (
        .q(_fractB_51_PC__q),
        .d(_fractB_51_PC__d),
        .clk(clock)
    );
    wire [1:0] _roundingMode_PC__q;
    wire [1:0] _roundingMode_PC__d;
    DFF_POSCLK #(.width(2)) roundingMode_PC (
        .q(_roundingMode_PC__q),
        .d(_roundingMode_PC__d),
        .clk(clock)
    );
    wire [13:0] _exp_PC__q;
    wire [13:0] _exp_PC__d;
    DFF_POSCLK #(.width(14)) exp_PC (
        .q(_exp_PC__q),
        .d(_exp_PC__d),
        .clk(clock)
    );
    wire _fractA_0_PC__q;
    wire _fractA_0_PC__d;
    DFF_POSCLK #(.width(1)) fractA_0_PC (
        .q(_fractA_0_PC__q),
        .d(_fractA_0_PC__d),
        .clk(clock)
    );
    wire [50:0] _fractB_other_PC__q;
    wire [50:0] _fractB_other_PC__d;
    DFF_POSCLK #(.width(51)) fractB_other_PC (
        .q(_fractB_other_PC__q),
        .d(_fractB_other_PC__d),
        .clk(clock)
    );
    wire [2:0] _cycleNum_A__q;
    wire [2:0] _cycleNum_A__d;
    DFF_POSCLK #(.width(3)) cycleNum_A (
        .q(_cycleNum_A__q),
        .d(_cycleNum_A__d),
        .clk(clock)
    );
    wire [2:0] _WTEMP_694;
    MUX_UNSIGNED #(.width(3)) u_mux_4935 (
        .y(_cycleNum_A__d),
        .sel(reset),
        .a(3'h0),
        .b(_WTEMP_694)
    );
    wire [3:0] _cycleNum_B__q;
    wire [3:0] _cycleNum_B__d;
    DFF_POSCLK #(.width(4)) cycleNum_B (
        .q(_cycleNum_B__q),
        .d(_cycleNum_B__d),
        .clk(clock)
    );
    wire [3:0] _WTEMP_695;
    MUX_UNSIGNED #(.width(4)) u_mux_4936 (
        .y(_cycleNum_B__d),
        .sel(reset),
        .a(4'h0),
        .b(_WTEMP_695)
    );
    wire [2:0] _cycleNum_C__q;
    wire [2:0] _cycleNum_C__d;
    DFF_POSCLK #(.width(3)) cycleNum_C (
        .q(_cycleNum_C__q),
        .d(_cycleNum_C__d),
        .clk(clock)
    );
    wire [2:0] _WTEMP_696;
    MUX_UNSIGNED #(.width(3)) u_mux_4937 (
        .y(_cycleNum_C__d),
        .sel(reset),
        .a(3'h0),
        .b(_WTEMP_696)
    );
    wire [2:0] _cycleNum_E__q;
    wire [2:0] _cycleNum_E__d;
    DFF_POSCLK #(.width(3)) cycleNum_E (
        .q(_cycleNum_E__q),
        .d(_cycleNum_E__d),
        .clk(clock)
    );
    wire [2:0] _WTEMP_697;
    MUX_UNSIGNED #(.width(3)) u_mux_4938 (
        .y(_cycleNum_E__d),
        .sel(reset),
        .a(3'h0),
        .b(_WTEMP_697)
    );
    wire [8:0] _fractR0_A__q;
    wire [8:0] _fractR0_A__d;
    DFF_POSCLK #(.width(9)) fractR0_A (
        .q(_fractR0_A__q),
        .d(_fractR0_A__d),
        .clk(clock)
    );
    wire [9:0] _hiSqrR0_A_sqrt__q;
    wire [9:0] _hiSqrR0_A_sqrt__d;
    DFF_POSCLK #(.width(10)) hiSqrR0_A_sqrt (
        .q(_hiSqrR0_A_sqrt__q),
        .d(_hiSqrR0_A_sqrt__d),
        .clk(clock)
    );
    wire [20:0] _partNegSigma0_A__q;
    wire [20:0] _partNegSigma0_A__d;
    DFF_POSCLK #(.width(21)) partNegSigma0_A (
        .q(_partNegSigma0_A__q),
        .d(_partNegSigma0_A__d),
        .clk(clock)
    );
    wire [8:0] _nextMulAdd9A_A__q;
    wire [8:0] _nextMulAdd9A_A__d;
    DFF_POSCLK #(.width(9)) nextMulAdd9A_A (
        .q(_nextMulAdd9A_A__q),
        .d(_nextMulAdd9A_A__d),
        .clk(clock)
    );
    wire [8:0] _nextMulAdd9B_A__q;
    wire [8:0] _nextMulAdd9B_A__d;
    DFF_POSCLK #(.width(9)) nextMulAdd9B_A (
        .q(_nextMulAdd9B_A__q),
        .d(_nextMulAdd9B_A__d),
        .clk(clock)
    );
    wire [16:0] _ER1_B_sqrt__q;
    wire [16:0] _ER1_B_sqrt__d;
    DFF_POSCLK #(.width(17)) ER1_B_sqrt (
        .q(_ER1_B_sqrt__q),
        .d(_ER1_B_sqrt__d),
        .clk(clock)
    );
    wire [31:0] _ESqrR1_B_sqrt__q;
    wire [31:0] _ESqrR1_B_sqrt__d;
    DFF_POSCLK #(.width(32)) ESqrR1_B_sqrt (
        .q(_ESqrR1_B_sqrt__q),
        .d(_ESqrR1_B_sqrt__d),
        .clk(clock)
    );
    wire [57:0] _sigX1_B__q;
    wire [57:0] _sigX1_B__d;
    DFF_POSCLK #(.width(58)) sigX1_B (
        .q(_sigX1_B__q),
        .d(_sigX1_B__d),
        .clk(clock)
    );
    wire [32:0] _sqrSigma1_C__q;
    wire [32:0] _sqrSigma1_C__d;
    DFF_POSCLK #(.width(33)) sqrSigma1_C (
        .q(_sqrSigma1_C__q),
        .d(_sqrSigma1_C__d),
        .clk(clock)
    );
    wire [57:0] _sigXN_C__q;
    wire [57:0] _sigXN_C__d;
    DFF_POSCLK #(.width(58)) sigXN_C (
        .q(_sigXN_C__q),
        .d(_sigXN_C__d),
        .clk(clock)
    );
    wire [30:0] _u_C_sqrt__q;
    wire [30:0] _u_C_sqrt__d;
    DFF_POSCLK #(.width(31)) u_C_sqrt (
        .q(_u_C_sqrt__q),
        .d(_u_C_sqrt__d),
        .clk(clock)
    );
    wire _E_E_div__q;
    wire _E_E_div__d;
    DFF_POSCLK #(.width(1)) E_E_div (
        .q(_E_E_div__q),
        .d(_E_E_div__d),
        .clk(clock)
    );
    wire [52:0] _sigT_E__q;
    wire [52:0] _sigT_E__d;
    DFF_POSCLK #(.width(53)) sigT_E (
        .q(_sigT_E__q),
        .d(_sigT_E__d),
        .clk(clock)
    );
    wire _extraT_E__q;
    wire _extraT_E__d;
    DFF_POSCLK #(.width(1)) extraT_E (
        .q(_extraT_E__q),
        .d(_extraT_E__d),
        .clk(clock)
    );
    wire _isNegRemT_E__q;
    wire _isNegRemT_E__d;
    DFF_POSCLK #(.width(1)) isNegRemT_E (
        .q(_isNegRemT_E__q),
        .d(_isNegRemT_E__d),
        .clk(clock)
    );
    wire _isZeroRemT_E__q;
    wire _isZeroRemT_E__d;
    DFF_POSCLK #(.width(1)) isZeroRemT_E (
        .q(_isZeroRemT_E__q),
        .d(_isZeroRemT_E__d),
        .clk(clock)
    );
    wire ready_PA;
    wire ready_PB;
    wire ready_PC;
    wire leaving_PA;
    wire leaving_PB;
    wire leaving_PC;
    wire cyc_B10_sqrt;
    wire cyc_B9_sqrt;
    wire cyc_B8_sqrt;
    wire cyc_B7_sqrt;
    wire cyc_B6;
    wire cyc_B5;
    wire cyc_B4;
    wire cyc_B3;
    wire cyc_B2;
    wire cyc_B1;
    wire cyc_B6_div;
    wire cyc_B5_div;
    wire cyc_B4_div;
    wire cyc_B3_div;
    wire cyc_B2_div;
    wire cyc_B1_div;
    wire cyc_B6_sqrt;
    wire cyc_B5_sqrt;
    wire cyc_B4_sqrt;
    wire cyc_B3_sqrt;
    wire cyc_B2_sqrt;
    wire cyc_B1_sqrt;
    wire cyc_C5;
    wire cyc_C4;
    wire cyc_C3;
    wire cyc_C2;
    wire cyc_C1;
    wire cyc_E4;
    wire cyc_E3;
    wire cyc_E2;
    wire cyc_E1;
    wire [45:0] zSigma1_B4;
    wire [57:0] sigXNU_B3_CX;
    wire [53:0] zComplSigT_C1_sqrt;
    wire [53:0] zComplSigT_C1;
    wire _T_133;
    EQ_UNSIGNED #(.width(1)) u_eq_4939 (
        .y(_T_133),
        .a(cyc_B7_sqrt),
        .b(1'h0)
    );
    wire _T_134;
    BITWISEAND #(.width(1)) bitwiseand_4940 (
        .y(_T_134),
        .a(ready_PA),
        .b(_T_133)
    );
    wire _T_136;
    EQ_UNSIGNED #(.width(1)) u_eq_4941 (
        .y(_T_136),
        .a(cyc_B6_sqrt),
        .b(1'h0)
    );
    wire _T_137;
    BITWISEAND #(.width(1)) bitwiseand_4942 (
        .y(_T_137),
        .a(_T_134),
        .b(_T_136)
    );
    wire _T_139;
    EQ_UNSIGNED #(.width(1)) u_eq_4943 (
        .y(_T_139),
        .a(cyc_B5_sqrt),
        .b(1'h0)
    );
    wire _T_140;
    BITWISEAND #(.width(1)) bitwiseand_4944 (
        .y(_T_140),
        .a(_T_137),
        .b(_T_139)
    );
    wire _T_142;
    EQ_UNSIGNED #(.width(1)) u_eq_4945 (
        .y(_T_142),
        .a(cyc_B4_sqrt),
        .b(1'h0)
    );
    wire _T_143;
    BITWISEAND #(.width(1)) bitwiseand_4946 (
        .y(_T_143),
        .a(_T_140),
        .b(_T_142)
    );
    wire _T_145;
    EQ_UNSIGNED #(.width(1)) u_eq_4947 (
        .y(_T_145),
        .a(cyc_B3),
        .b(1'h0)
    );
    wire _T_146;
    BITWISEAND #(.width(1)) bitwiseand_4948 (
        .y(_T_146),
        .a(_T_143),
        .b(_T_145)
    );
    wire _T_148;
    EQ_UNSIGNED #(.width(1)) u_eq_4949 (
        .y(_T_148),
        .a(cyc_B2),
        .b(1'h0)
    );
    wire _T_149;
    BITWISEAND #(.width(1)) bitwiseand_4950 (
        .y(_T_149),
        .a(_T_146),
        .b(_T_148)
    );
    wire _T_151;
    EQ_UNSIGNED #(.width(1)) u_eq_4951 (
        .y(_T_151),
        .a(cyc_B1_sqrt),
        .b(1'h0)
    );
    wire _T_152;
    BITWISEAND #(.width(1)) bitwiseand_4952 (
        .y(_T_152),
        .a(_T_149),
        .b(_T_151)
    );
    wire _T_154;
    EQ_UNSIGNED #(.width(1)) u_eq_4953 (
        .y(_T_154),
        .a(cyc_C5),
        .b(1'h0)
    );
    wire _T_155;
    BITWISEAND #(.width(1)) bitwiseand_4954 (
        .y(_T_155),
        .a(_T_152),
        .b(_T_154)
    );
    wire _T_157;
    EQ_UNSIGNED #(.width(1)) u_eq_4955 (
        .y(_T_157),
        .a(cyc_C4),
        .b(1'h0)
    );
    wire _T_158;
    BITWISEAND #(.width(1)) bitwiseand_4956 (
        .y(_T_158),
        .a(_T_155),
        .b(_T_157)
    );
    wire _T_160;
    EQ_UNSIGNED #(.width(1)) u_eq_4957 (
        .y(_T_160),
        .a(cyc_B6_sqrt),
        .b(1'h0)
    );
    wire _T_161;
    BITWISEAND #(.width(1)) bitwiseand_4958 (
        .y(_T_161),
        .a(ready_PA),
        .b(_T_160)
    );
    wire _T_163;
    EQ_UNSIGNED #(.width(1)) u_eq_4959 (
        .y(_T_163),
        .a(cyc_B5_sqrt),
        .b(1'h0)
    );
    wire _T_164;
    BITWISEAND #(.width(1)) bitwiseand_4960 (
        .y(_T_164),
        .a(_T_161),
        .b(_T_163)
    );
    wire _T_166;
    EQ_UNSIGNED #(.width(1)) u_eq_4961 (
        .y(_T_166),
        .a(cyc_B4_sqrt),
        .b(1'h0)
    );
    wire _T_167;
    BITWISEAND #(.width(1)) bitwiseand_4962 (
        .y(_T_167),
        .a(_T_164),
        .b(_T_166)
    );
    wire _T_169;
    EQ_UNSIGNED #(.width(1)) u_eq_4963 (
        .y(_T_169),
        .a(cyc_B2_div),
        .b(1'h0)
    );
    wire _T_170;
    BITWISEAND #(.width(1)) bitwiseand_4964 (
        .y(_T_170),
        .a(_T_167),
        .b(_T_169)
    );
    wire _T_172;
    EQ_UNSIGNED #(.width(1)) u_eq_4965 (
        .y(_T_172),
        .a(cyc_B1_sqrt),
        .b(1'h0)
    );
    wire _T_173;
    BITWISEAND #(.width(1)) bitwiseand_4966 (
        .y(_T_173),
        .a(_T_170),
        .b(_T_172)
    );
    wire _T_174;
    BITWISEAND #(.width(1)) bitwiseand_4967 (
        .y(_T_174),
        .a(io_inReady_div),
        .b(io_inValid)
    );
    wire _T_176;
    EQ_UNSIGNED #(.width(1)) u_eq_4968 (
        .y(_T_176),
        .a(io_sqrtOp),
        .b(1'h0)
    );
    wire cyc_S_div;
    BITWISEAND #(.width(1)) bitwiseand_4969 (
        .y(cyc_S_div),
        .a(_T_174),
        .b(_T_176)
    );
    wire _T_177;
    BITWISEAND #(.width(1)) bitwiseand_4970 (
        .y(_T_177),
        .a(io_inReady_sqrt),
        .b(io_inValid)
    );
    wire cyc_S_sqrt;
    BITWISEAND #(.width(1)) bitwiseand_4971 (
        .y(cyc_S_sqrt),
        .a(_T_177),
        .b(io_sqrtOp)
    );
    wire cyc_S;
    BITWISEOR #(.width(1)) bitwiseor_4972 (
        .y(cyc_S),
        .a(cyc_S_div),
        .b(cyc_S_sqrt)
    );
    wire signA_S;
    BITS #(.width(65), .high(64), .low(64)) bits_4973 (
        .y(signA_S),
        .in(io_a)
    );
    wire [11:0] expA_S;
    BITS #(.width(65), .high(63), .low(52)) bits_4974 (
        .y(expA_S),
        .in(io_a)
    );
    wire [51:0] fractA_S;
    BITS #(.width(65), .high(51), .low(0)) bits_4975 (
        .y(fractA_S),
        .in(io_a)
    );
    wire [2:0] specialCodeA_S;
    BITS #(.width(12), .high(11), .low(9)) bits_4976 (
        .y(specialCodeA_S),
        .in(expA_S)
    );
    wire isZeroA_S;
    EQ_UNSIGNED #(.width(3)) u_eq_4977 (
        .y(isZeroA_S),
        .a(specialCodeA_S),
        .b(3'h0)
    );
    wire [1:0] _T_179;
    BITS #(.width(3), .high(2), .low(1)) bits_4978 (
        .y(_T_179),
        .in(specialCodeA_S)
    );
    wire isSpecialA_S;
    EQ_UNSIGNED #(.width(2)) u_eq_4979 (
        .y(isSpecialA_S),
        .a(_T_179),
        .b(2'h3)
    );
    wire signB_S;
    BITS #(.width(65), .high(64), .low(64)) bits_4980 (
        .y(signB_S),
        .in(io_b)
    );
    wire [11:0] expB_S;
    BITS #(.width(65), .high(63), .low(52)) bits_4981 (
        .y(expB_S),
        .in(io_b)
    );
    wire [51:0] fractB_S;
    BITS #(.width(65), .high(51), .low(0)) bits_4982 (
        .y(fractB_S),
        .in(io_b)
    );
    wire [2:0] specialCodeB_S;
    BITS #(.width(12), .high(11), .low(9)) bits_4983 (
        .y(specialCodeB_S),
        .in(expB_S)
    );
    wire isZeroB_S;
    EQ_UNSIGNED #(.width(3)) u_eq_4984 (
        .y(isZeroB_S),
        .a(specialCodeB_S),
        .b(3'h0)
    );
    wire [1:0] _T_182;
    BITS #(.width(3), .high(2), .low(1)) bits_4985 (
        .y(_T_182),
        .in(specialCodeB_S)
    );
    wire isSpecialB_S;
    EQ_UNSIGNED #(.width(2)) u_eq_4986 (
        .y(isSpecialB_S),
        .a(_T_182),
        .b(2'h3)
    );
    wire _T_184;
    BITWISEXOR #(.width(1)) bitwisexor_4987 (
        .y(_T_184),
        .a(signA_S),
        .b(signB_S)
    );
    wire sign_S;
    MUX_UNSIGNED #(.width(1)) u_mux_4988 (
        .y(sign_S),
        .sel(io_sqrtOp),
        .a(signB_S),
        .b(_T_184)
    );
    wire _T_186;
    EQ_UNSIGNED #(.width(1)) u_eq_4989 (
        .y(_T_186),
        .a(isSpecialA_S),
        .b(1'h0)
    );
    wire _T_188;
    EQ_UNSIGNED #(.width(1)) u_eq_4990 (
        .y(_T_188),
        .a(isSpecialB_S),
        .b(1'h0)
    );
    wire _T_189;
    BITWISEAND #(.width(1)) bitwiseand_4991 (
        .y(_T_189),
        .a(_T_186),
        .b(_T_188)
    );
    wire _T_191;
    EQ_UNSIGNED #(.width(1)) u_eq_4992 (
        .y(_T_191),
        .a(isZeroA_S),
        .b(1'h0)
    );
    wire _T_192;
    BITWISEAND #(.width(1)) bitwiseand_4993 (
        .y(_T_192),
        .a(_T_189),
        .b(_T_191)
    );
    wire _T_194;
    EQ_UNSIGNED #(.width(1)) u_eq_4994 (
        .y(_T_194),
        .a(isZeroB_S),
        .b(1'h0)
    );
    wire normalCase_S_div;
    BITWISEAND #(.width(1)) bitwiseand_4995 (
        .y(normalCase_S_div),
        .a(_T_192),
        .b(_T_194)
    );
    wire _T_196;
    EQ_UNSIGNED #(.width(1)) u_eq_4996 (
        .y(_T_196),
        .a(isSpecialB_S),
        .b(1'h0)
    );
    wire _T_198;
    EQ_UNSIGNED #(.width(1)) u_eq_4997 (
        .y(_T_198),
        .a(isZeroB_S),
        .b(1'h0)
    );
    wire _T_199;
    BITWISEAND #(.width(1)) bitwiseand_4998 (
        .y(_T_199),
        .a(_T_196),
        .b(_T_198)
    );
    wire _T_201;
    EQ_UNSIGNED #(.width(1)) u_eq_4999 (
        .y(_T_201),
        .a(signB_S),
        .b(1'h0)
    );
    wire normalCase_S_sqrt;
    BITWISEAND #(.width(1)) bitwiseand_5000 (
        .y(normalCase_S_sqrt),
        .a(_T_199),
        .b(_T_201)
    );
    wire normalCase_S;
    MUX_UNSIGNED #(.width(1)) u_mux_5001 (
        .y(normalCase_S),
        .sel(io_sqrtOp),
        .a(normalCase_S_sqrt),
        .b(normalCase_S_div)
    );
    wire cyc_A4_div;
    BITWISEAND #(.width(1)) bitwiseand_5002 (
        .y(cyc_A4_div),
        .a(cyc_S_div),
        .b(normalCase_S_div)
    );
    wire cyc_A7_sqrt;
    BITWISEAND #(.width(1)) bitwiseand_5003 (
        .y(cyc_A7_sqrt),
        .a(cyc_S_sqrt),
        .b(normalCase_S_sqrt)
    );
    wire entering_PA_normalCase;
    BITWISEOR #(.width(1)) bitwiseor_5004 (
        .y(entering_PA_normalCase),
        .a(cyc_A4_div),
        .b(cyc_A7_sqrt)
    );
    wire _T_203;
    EQ_UNSIGNED #(.width(1)) u_eq_5005 (
        .y(_T_203),
        .a(ready_PB),
        .b(1'h0)
    );
    wire _T_204;
    BITWISEOR #(.width(1)) bitwiseor_5006 (
        .y(_T_204),
        .a(_valid_PA__q),
        .b(_T_203)
    );
    wire _T_205;
    BITWISEAND #(.width(1)) bitwiseand_5007 (
        .y(_T_205),
        .a(cyc_S),
        .b(_T_204)
    );
    wire entering_PA;
    BITWISEOR #(.width(1)) bitwiseor_5008 (
        .y(entering_PA),
        .a(entering_PA_normalCase),
        .b(_T_205)
    );
    wire _T_207;
    EQ_UNSIGNED #(.width(1)) u_eq_5009 (
        .y(_T_207),
        .a(normalCase_S),
        .b(1'h0)
    );
    wire _T_208;
    BITWISEAND #(.width(1)) bitwiseand_5010 (
        .y(_T_208),
        .a(cyc_S),
        .b(_T_207)
    );
    wire _T_210;
    EQ_UNSIGNED #(.width(1)) u_eq_5011 (
        .y(_T_210),
        .a(_valid_PA__q),
        .b(1'h0)
    );
    wire _T_211;
    BITWISEAND #(.width(1)) bitwiseand_5012 (
        .y(_T_211),
        .a(_T_208),
        .b(_T_210)
    );
    wire _T_213;
    EQ_UNSIGNED #(.width(1)) u_eq_5013 (
        .y(_T_213),
        .a(_valid_PB__q),
        .b(1'h0)
    );
    wire _T_215;
    EQ_UNSIGNED #(.width(1)) u_eq_5014 (
        .y(_T_215),
        .a(ready_PC),
        .b(1'h0)
    );
    wire _T_216;
    BITWISEAND #(.width(1)) bitwiseand_5015 (
        .y(_T_216),
        .a(_T_213),
        .b(_T_215)
    );
    wire _T_217;
    BITWISEOR #(.width(1)) bitwiseor_5016 (
        .y(_T_217),
        .a(leaving_PB),
        .b(_T_216)
    );
    wire entering_PB_S;
    BITWISEAND #(.width(1)) bitwiseand_5017 (
        .y(entering_PB_S),
        .a(_T_211),
        .b(_T_217)
    );
    wire _T_219;
    EQ_UNSIGNED #(.width(1)) u_eq_5018 (
        .y(_T_219),
        .a(normalCase_S),
        .b(1'h0)
    );
    wire _T_220;
    BITWISEAND #(.width(1)) bitwiseand_5019 (
        .y(_T_220),
        .a(cyc_S),
        .b(_T_219)
    );
    wire _T_222;
    EQ_UNSIGNED #(.width(1)) u_eq_5020 (
        .y(_T_222),
        .a(_valid_PA__q),
        .b(1'h0)
    );
    wire _T_223;
    BITWISEAND #(.width(1)) bitwiseand_5021 (
        .y(_T_223),
        .a(_T_220),
        .b(_T_222)
    );
    wire _T_225;
    EQ_UNSIGNED #(.width(1)) u_eq_5022 (
        .y(_T_225),
        .a(_valid_PB__q),
        .b(1'h0)
    );
    wire _T_226;
    BITWISEAND #(.width(1)) bitwiseand_5023 (
        .y(_T_226),
        .a(_T_223),
        .b(_T_225)
    );
    wire entering_PC_S;
    BITWISEAND #(.width(1)) bitwiseand_5024 (
        .y(entering_PC_S),
        .a(_T_226),
        .b(ready_PC)
    );
    wire _T_227;
    BITWISEOR #(.width(1)) bitwiseor_5025 (
        .y(_T_227),
        .a(entering_PA),
        .b(leaving_PA)
    );
    wire _T_228;
    BITS #(.width(52), .high(51), .low(51)) bits_5026 (
        .y(_T_228),
        .in(fractB_S)
    );
    wire _T_230;
    EQ_UNSIGNED #(.width(1)) u_eq_5027 (
        .y(_T_230),
        .a(io_sqrtOp),
        .b(1'h0)
    );
    wire _T_231;
    BITWISEAND #(.width(1)) bitwiseand_5028 (
        .y(_T_231),
        .a(entering_PA),
        .b(_T_230)
    );
    wire _T_232;
    BITS #(.width(52), .high(51), .low(51)) bits_5029 (
        .y(_T_232),
        .in(fractA_S)
    );
    wire _T_233;
    BITS #(.width(12), .high(11), .low(11)) bits_5030 (
        .y(_T_233),
        .in(expB_S)
    );
    wire _T_234;
    BITS #(.width(1), .high(0), .low(0)) bits_5031 (
        .y(_T_234),
        .in(_T_233)
    );
    wire [2:0] _T_237;
    MUX_UNSIGNED #(.width(3)) u_mux_5032 (
        .y(_T_237),
        .sel(_T_234),
        .a(3'h7),
        .b(3'h0)
    );
    wire [10:0] _T_238;
    BITS #(.width(12), .high(10), .low(0)) bits_5033 (
        .y(_T_238),
        .in(expB_S)
    );
    wire [10:0] _T_239;
    BITWISENOT #(.width(11)) bitwisenot_5034 (
        .y(_T_239),
        .in(_T_238)
    );
    wire [13:0] _T_240;
    CAT #(.width_a(3), .width_b(11)) cat_5035 (
        .y(_T_240),
        .a(_T_237),
        .b(_T_239)
    );
    wire [14:0] _T_241;
    wire [13:0] _WTEMP_698;
    PAD_UNSIGNED #(.width(12), .n(14)) u_pad_5036 (
        .y(_WTEMP_698),
        .in(expA_S)
    );
    ADD_UNSIGNED #(.width(14)) u_add_5037 (
        .y(_T_241),
        .a(_WTEMP_698),
        .b(_T_240)
    );
    wire [13:0] _T_242;
    TAIL #(.width(15), .n(1)) tail_5038 (
        .y(_T_242),
        .in(_T_241)
    );
    wire [13:0] _T_243;
    wire [13:0] _WTEMP_699;
    PAD_UNSIGNED #(.width(12), .n(14)) u_pad_5039 (
        .y(_WTEMP_699),
        .in(expB_S)
    );
    MUX_UNSIGNED #(.width(14)) u_mux_5040 (
        .y(_T_243),
        .sel(io_sqrtOp),
        .a(_WTEMP_699),
        .b(_T_242)
    );
    wire [50:0] _T_244;
    BITS #(.width(52), .high(50), .low(0)) bits_5041 (
        .y(_T_244),
        .in(fractB_S)
    );
    wire [50:0] _T_245;
    BITS #(.width(52), .high(50), .low(0)) bits_5042 (
        .y(_T_245),
        .in(fractA_S)
    );
    wire isZeroA_PA;
    EQ_UNSIGNED #(.width(3)) u_eq_5043 (
        .y(isZeroA_PA),
        .a(_specialCodeA_PA__q),
        .b(3'h0)
    );
    wire [1:0] _T_247;
    BITS #(.width(3), .high(2), .low(1)) bits_5044 (
        .y(_T_247),
        .in(_specialCodeA_PA__q)
    );
    wire isSpecialA_PA;
    EQ_UNSIGNED #(.width(2)) u_eq_5045 (
        .y(isSpecialA_PA),
        .a(_T_247),
        .b(2'h3)
    );
    wire [1:0] _T_250;
    CAT #(.width_a(1), .width_b(1)) cat_5046 (
        .y(_T_250),
        .a(1'h1),
        .b(_fractA_51_PA__q)
    );
    wire [52:0] sigA_PA;
    CAT #(.width_a(2), .width_b(51)) cat_5047 (
        .y(sigA_PA),
        .a(_T_250),
        .b(_fractA_other_PA__q)
    );
    wire isZeroB_PA;
    EQ_UNSIGNED #(.width(3)) u_eq_5048 (
        .y(isZeroB_PA),
        .a(_specialCodeB_PA__q),
        .b(3'h0)
    );
    wire [1:0] _T_252;
    BITS #(.width(3), .high(2), .low(1)) bits_5049 (
        .y(_T_252),
        .in(_specialCodeB_PA__q)
    );
    wire isSpecialB_PA;
    EQ_UNSIGNED #(.width(2)) u_eq_5050 (
        .y(isSpecialB_PA),
        .a(_T_252),
        .b(2'h3)
    );
    wire [1:0] _T_255;
    CAT #(.width_a(1), .width_b(1)) cat_5051 (
        .y(_T_255),
        .a(1'h1),
        .b(_fractB_51_PA__q)
    );
    wire [52:0] sigB_PA;
    CAT #(.width_a(2), .width_b(51)) cat_5052 (
        .y(sigB_PA),
        .a(_T_255),
        .b(_fractB_other_PA__q)
    );
    wire _T_257;
    EQ_UNSIGNED #(.width(1)) u_eq_5053 (
        .y(_T_257),
        .a(isSpecialB_PA),
        .b(1'h0)
    );
    wire _T_259;
    EQ_UNSIGNED #(.width(1)) u_eq_5054 (
        .y(_T_259),
        .a(isZeroB_PA),
        .b(1'h0)
    );
    wire _T_260;
    BITWISEAND #(.width(1)) bitwiseand_5055 (
        .y(_T_260),
        .a(_T_257),
        .b(_T_259)
    );
    wire _T_262;
    EQ_UNSIGNED #(.width(1)) u_eq_5056 (
        .y(_T_262),
        .a(_sign_PA__q),
        .b(1'h0)
    );
    wire _T_263;
    BITWISEAND #(.width(1)) bitwiseand_5057 (
        .y(_T_263),
        .a(_T_260),
        .b(_T_262)
    );
    wire _T_265;
    EQ_UNSIGNED #(.width(1)) u_eq_5058 (
        .y(_T_265),
        .a(isSpecialA_PA),
        .b(1'h0)
    );
    wire _T_267;
    EQ_UNSIGNED #(.width(1)) u_eq_5059 (
        .y(_T_267),
        .a(isSpecialB_PA),
        .b(1'h0)
    );
    wire _T_268;
    BITWISEAND #(.width(1)) bitwiseand_5060 (
        .y(_T_268),
        .a(_T_265),
        .b(_T_267)
    );
    wire _T_270;
    EQ_UNSIGNED #(.width(1)) u_eq_5061 (
        .y(_T_270),
        .a(isZeroA_PA),
        .b(1'h0)
    );
    wire _T_271;
    BITWISEAND #(.width(1)) bitwiseand_5062 (
        .y(_T_271),
        .a(_T_268),
        .b(_T_270)
    );
    wire _T_273;
    EQ_UNSIGNED #(.width(1)) u_eq_5063 (
        .y(_T_273),
        .a(isZeroB_PA),
        .b(1'h0)
    );
    wire _T_274;
    BITWISEAND #(.width(1)) bitwiseand_5064 (
        .y(_T_274),
        .a(_T_271),
        .b(_T_273)
    );
    wire normalCase_PA;
    MUX_UNSIGNED #(.width(1)) u_mux_5065 (
        .y(normalCase_PA),
        .sel(_sqrtOp_PA__q),
        .a(_T_263),
        .b(_T_274)
    );
    wire valid_normalCase_leaving_PA;
    BITWISEOR #(.width(1)) bitwiseor_5066 (
        .y(valid_normalCase_leaving_PA),
        .a(cyc_B4_div),
        .b(cyc_B7_sqrt)
    );
    wire valid_leaving_PA;
    MUX_UNSIGNED #(.width(1)) u_mux_5067 (
        .y(valid_leaving_PA),
        .sel(normalCase_PA),
        .a(valid_normalCase_leaving_PA),
        .b(ready_PB)
    );
    wire _T_275;
    BITWISEAND #(.width(1)) bitwiseand_5068 (
        .y(_T_275),
        .a(_valid_PA__q),
        .b(valid_leaving_PA)
    );
    wire _T_277;
    EQ_UNSIGNED #(.width(1)) u_eq_5069 (
        .y(_T_277),
        .a(_valid_PA__q),
        .b(1'h0)
    );
    wire _T_278;
    BITWISEOR #(.width(1)) bitwiseor_5070 (
        .y(_T_278),
        .a(_T_277),
        .b(valid_leaving_PA)
    );
    wire _T_279;
    BITWISEAND #(.width(1)) bitwiseand_5071 (
        .y(_T_279),
        .a(_valid_PA__q),
        .b(normalCase_PA)
    );
    wire entering_PB_normalCase;
    BITWISEAND #(.width(1)) bitwiseand_5072 (
        .y(entering_PB_normalCase),
        .a(_T_279),
        .b(valid_normalCase_leaving_PA)
    );
    wire entering_PB;
    BITWISEOR #(.width(1)) bitwiseor_5073 (
        .y(entering_PB),
        .a(entering_PB_S),
        .b(leaving_PA)
    );
    wire _T_280;
    BITWISEOR #(.width(1)) bitwiseor_5074 (
        .y(_T_280),
        .a(entering_PB),
        .b(leaving_PB)
    );
    wire _T_281;
    MUX_UNSIGNED #(.width(1)) u_mux_5075 (
        .y(_T_281),
        .sel(_valid_PA__q),
        .a(_sqrtOp_PA__q),
        .b(io_sqrtOp)
    );
    wire _T_282;
    MUX_UNSIGNED #(.width(1)) u_mux_5076 (
        .y(_T_282),
        .sel(_valid_PA__q),
        .a(_sign_PA__q),
        .b(sign_S)
    );
    wire [2:0] _T_283;
    MUX_UNSIGNED #(.width(3)) u_mux_5077 (
        .y(_T_283),
        .sel(_valid_PA__q),
        .a(_specialCodeA_PA__q),
        .b(specialCodeA_S)
    );
    wire _T_284;
    BITS #(.width(52), .high(51), .low(51)) bits_5078 (
        .y(_T_284),
        .in(fractA_S)
    );
    wire _T_285;
    MUX_UNSIGNED #(.width(1)) u_mux_5079 (
        .y(_T_285),
        .sel(_valid_PA__q),
        .a(_fractA_51_PA__q),
        .b(_T_284)
    );
    wire [2:0] _T_286;
    MUX_UNSIGNED #(.width(3)) u_mux_5080 (
        .y(_T_286),
        .sel(_valid_PA__q),
        .a(_specialCodeB_PA__q),
        .b(specialCodeB_S)
    );
    wire _T_287;
    BITS #(.width(52), .high(51), .low(51)) bits_5081 (
        .y(_T_287),
        .in(fractB_S)
    );
    wire _T_288;
    MUX_UNSIGNED #(.width(1)) u_mux_5082 (
        .y(_T_288),
        .sel(_valid_PA__q),
        .a(_fractB_51_PA__q),
        .b(_T_287)
    );
    wire [1:0] _T_289;
    MUX_UNSIGNED #(.width(2)) u_mux_5083 (
        .y(_T_289),
        .sel(_valid_PA__q),
        .a(_roundingMode_PA__q),
        .b(io_roundingMode)
    );
    wire _T_290;
    BITS #(.width(51), .high(0), .low(0)) bits_5084 (
        .y(_T_290),
        .in(_fractA_other_PA__q)
    );
    wire isZeroA_PB;
    EQ_UNSIGNED #(.width(3)) u_eq_5085 (
        .y(isZeroA_PB),
        .a(_specialCodeA_PB__q),
        .b(3'h0)
    );
    wire [1:0] _T_292;
    BITS #(.width(3), .high(2), .low(1)) bits_5086 (
        .y(_T_292),
        .in(_specialCodeA_PB__q)
    );
    wire isSpecialA_PB;
    EQ_UNSIGNED #(.width(2)) u_eq_5087 (
        .y(isSpecialA_PB),
        .a(_T_292),
        .b(2'h3)
    );
    wire isZeroB_PB;
    EQ_UNSIGNED #(.width(3)) u_eq_5088 (
        .y(isZeroB_PB),
        .a(_specialCodeB_PB__q),
        .b(3'h0)
    );
    wire [1:0] _T_295;
    BITS #(.width(3), .high(2), .low(1)) bits_5089 (
        .y(_T_295),
        .in(_specialCodeB_PB__q)
    );
    wire isSpecialB_PB;
    EQ_UNSIGNED #(.width(2)) u_eq_5090 (
        .y(isSpecialB_PB),
        .a(_T_295),
        .b(2'h3)
    );
    wire _T_298;
    EQ_UNSIGNED #(.width(1)) u_eq_5091 (
        .y(_T_298),
        .a(isSpecialB_PB),
        .b(1'h0)
    );
    wire _T_300;
    EQ_UNSIGNED #(.width(1)) u_eq_5092 (
        .y(_T_300),
        .a(isZeroB_PB),
        .b(1'h0)
    );
    wire _T_301;
    BITWISEAND #(.width(1)) bitwiseand_5093 (
        .y(_T_301),
        .a(_T_298),
        .b(_T_300)
    );
    wire _T_303;
    EQ_UNSIGNED #(.width(1)) u_eq_5094 (
        .y(_T_303),
        .a(_sign_PB__q),
        .b(1'h0)
    );
    wire _T_304;
    BITWISEAND #(.width(1)) bitwiseand_5095 (
        .y(_T_304),
        .a(_T_301),
        .b(_T_303)
    );
    wire _T_306;
    EQ_UNSIGNED #(.width(1)) u_eq_5096 (
        .y(_T_306),
        .a(isSpecialA_PB),
        .b(1'h0)
    );
    wire _T_308;
    EQ_UNSIGNED #(.width(1)) u_eq_5097 (
        .y(_T_308),
        .a(isSpecialB_PB),
        .b(1'h0)
    );
    wire _T_309;
    BITWISEAND #(.width(1)) bitwiseand_5098 (
        .y(_T_309),
        .a(_T_306),
        .b(_T_308)
    );
    wire _T_311;
    EQ_UNSIGNED #(.width(1)) u_eq_5099 (
        .y(_T_311),
        .a(isZeroA_PB),
        .b(1'h0)
    );
    wire _T_312;
    BITWISEAND #(.width(1)) bitwiseand_5100 (
        .y(_T_312),
        .a(_T_309),
        .b(_T_311)
    );
    wire _T_314;
    EQ_UNSIGNED #(.width(1)) u_eq_5101 (
        .y(_T_314),
        .a(isZeroB_PB),
        .b(1'h0)
    );
    wire _T_315;
    BITWISEAND #(.width(1)) bitwiseand_5102 (
        .y(_T_315),
        .a(_T_312),
        .b(_T_314)
    );
    wire normalCase_PB;
    MUX_UNSIGNED #(.width(1)) u_mux_5103 (
        .y(normalCase_PB),
        .sel(_sqrtOp_PB__q),
        .a(_T_304),
        .b(_T_315)
    );
    wire valid_leaving_PB;
    MUX_UNSIGNED #(.width(1)) u_mux_5104 (
        .y(valid_leaving_PB),
        .sel(normalCase_PB),
        .a(cyc_C3),
        .b(ready_PC)
    );
    wire _T_316;
    BITWISEAND #(.width(1)) bitwiseand_5105 (
        .y(_T_316),
        .a(_valid_PB__q),
        .b(valid_leaving_PB)
    );
    wire _T_318;
    EQ_UNSIGNED #(.width(1)) u_eq_5106 (
        .y(_T_318),
        .a(_valid_PB__q),
        .b(1'h0)
    );
    wire _T_319;
    BITWISEOR #(.width(1)) bitwiseor_5107 (
        .y(_T_319),
        .a(_T_318),
        .b(valid_leaving_PB)
    );
    wire _T_320;
    BITWISEAND #(.width(1)) bitwiseand_5108 (
        .y(_T_320),
        .a(_valid_PB__q),
        .b(normalCase_PB)
    );
    wire entering_PC_normalCase;
    BITWISEAND #(.width(1)) bitwiseand_5109 (
        .y(entering_PC_normalCase),
        .a(_T_320),
        .b(cyc_C3)
    );
    wire entering_PC;
    BITWISEOR #(.width(1)) bitwiseor_5110 (
        .y(entering_PC),
        .a(entering_PC_S),
        .b(leaving_PB)
    );
    wire _T_321;
    BITWISEOR #(.width(1)) bitwiseor_5111 (
        .y(_T_321),
        .a(entering_PC),
        .b(leaving_PC)
    );
    wire _T_322;
    MUX_UNSIGNED #(.width(1)) u_mux_5112 (
        .y(_T_322),
        .sel(_valid_PB__q),
        .a(_sqrtOp_PB__q),
        .b(io_sqrtOp)
    );
    wire _T_323;
    MUX_UNSIGNED #(.width(1)) u_mux_5113 (
        .y(_T_323),
        .sel(_valid_PB__q),
        .a(_sign_PB__q),
        .b(sign_S)
    );
    wire [2:0] _T_324;
    MUX_UNSIGNED #(.width(3)) u_mux_5114 (
        .y(_T_324),
        .sel(_valid_PB__q),
        .a(_specialCodeA_PB__q),
        .b(specialCodeA_S)
    );
    wire _T_325;
    BITS #(.width(52), .high(51), .low(51)) bits_5115 (
        .y(_T_325),
        .in(fractA_S)
    );
    wire _T_326;
    MUX_UNSIGNED #(.width(1)) u_mux_5116 (
        .y(_T_326),
        .sel(_valid_PB__q),
        .a(_fractA_51_PB__q),
        .b(_T_325)
    );
    wire [2:0] _T_327;
    MUX_UNSIGNED #(.width(3)) u_mux_5117 (
        .y(_T_327),
        .sel(_valid_PB__q),
        .a(_specialCodeB_PB__q),
        .b(specialCodeB_S)
    );
    wire _T_328;
    BITS #(.width(52), .high(51), .low(51)) bits_5118 (
        .y(_T_328),
        .in(fractB_S)
    );
    wire _T_329;
    MUX_UNSIGNED #(.width(1)) u_mux_5119 (
        .y(_T_329),
        .sel(_valid_PB__q),
        .a(_fractB_51_PB__q),
        .b(_T_328)
    );
    wire [1:0] _T_330;
    MUX_UNSIGNED #(.width(2)) u_mux_5120 (
        .y(_T_330),
        .sel(_valid_PB__q),
        .a(_roundingMode_PB__q),
        .b(io_roundingMode)
    );
    wire isZeroA_PC;
    EQ_UNSIGNED #(.width(3)) u_eq_5121 (
        .y(isZeroA_PC),
        .a(_specialCodeA_PC__q),
        .b(3'h0)
    );
    wire [1:0] _T_332;
    BITS #(.width(3), .high(2), .low(1)) bits_5122 (
        .y(_T_332),
        .in(_specialCodeA_PC__q)
    );
    wire isSpecialA_PC;
    EQ_UNSIGNED #(.width(2)) u_eq_5123 (
        .y(isSpecialA_PC),
        .a(_T_332),
        .b(2'h3)
    );
    wire _T_334;
    BITS #(.width(3), .high(0), .low(0)) bits_5124 (
        .y(_T_334),
        .in(_specialCodeA_PC__q)
    );
    wire _T_336;
    EQ_UNSIGNED #(.width(1)) u_eq_5125 (
        .y(_T_336),
        .a(_T_334),
        .b(1'h0)
    );
    wire isInfA_PC;
    BITWISEAND #(.width(1)) bitwiseand_5126 (
        .y(isInfA_PC),
        .a(isSpecialA_PC),
        .b(_T_336)
    );
    wire _T_337;
    BITS #(.width(3), .high(0), .low(0)) bits_5127 (
        .y(_T_337),
        .in(_specialCodeA_PC__q)
    );
    wire isNaNA_PC;
    BITWISEAND #(.width(1)) bitwiseand_5128 (
        .y(isNaNA_PC),
        .a(isSpecialA_PC),
        .b(_T_337)
    );
    wire _T_339;
    EQ_UNSIGNED #(.width(1)) u_eq_5129 (
        .y(_T_339),
        .a(_fractA_51_PC__q),
        .b(1'h0)
    );
    wire isSigNaNA_PC;
    BITWISEAND #(.width(1)) bitwiseand_5130 (
        .y(isSigNaNA_PC),
        .a(isNaNA_PC),
        .b(_T_339)
    );
    wire isZeroB_PC;
    EQ_UNSIGNED #(.width(3)) u_eq_5131 (
        .y(isZeroB_PC),
        .a(_specialCodeB_PC__q),
        .b(3'h0)
    );
    wire [1:0] _T_341;
    BITS #(.width(3), .high(2), .low(1)) bits_5132 (
        .y(_T_341),
        .in(_specialCodeB_PC__q)
    );
    wire isSpecialB_PC;
    EQ_UNSIGNED #(.width(2)) u_eq_5133 (
        .y(isSpecialB_PC),
        .a(_T_341),
        .b(2'h3)
    );
    wire _T_343;
    BITS #(.width(3), .high(0), .low(0)) bits_5134 (
        .y(_T_343),
        .in(_specialCodeB_PC__q)
    );
    wire _T_345;
    EQ_UNSIGNED #(.width(1)) u_eq_5135 (
        .y(_T_345),
        .a(_T_343),
        .b(1'h0)
    );
    wire isInfB_PC;
    BITWISEAND #(.width(1)) bitwiseand_5136 (
        .y(isInfB_PC),
        .a(isSpecialB_PC),
        .b(_T_345)
    );
    wire _T_346;
    BITS #(.width(3), .high(0), .low(0)) bits_5137 (
        .y(_T_346),
        .in(_specialCodeB_PC__q)
    );
    wire isNaNB_PC;
    BITWISEAND #(.width(1)) bitwiseand_5138 (
        .y(isNaNB_PC),
        .a(isSpecialB_PC),
        .b(_T_346)
    );
    wire _T_348;
    EQ_UNSIGNED #(.width(1)) u_eq_5139 (
        .y(_T_348),
        .a(_fractB_51_PC__q),
        .b(1'h0)
    );
    wire isSigNaNB_PC;
    BITWISEAND #(.width(1)) bitwiseand_5140 (
        .y(isSigNaNB_PC),
        .a(isNaNB_PC),
        .b(_T_348)
    );
    wire [1:0] _T_350;
    CAT #(.width_a(1), .width_b(1)) cat_5141 (
        .y(_T_350),
        .a(1'h1),
        .b(_fractB_51_PC__q)
    );
    wire [52:0] sigB_PC;
    CAT #(.width_a(2), .width_b(51)) cat_5142 (
        .y(sigB_PC),
        .a(_T_350),
        .b(_fractB_other_PC__q)
    );
    wire _T_352;
    EQ_UNSIGNED #(.width(1)) u_eq_5143 (
        .y(_T_352),
        .a(isSpecialB_PC),
        .b(1'h0)
    );
    wire _T_354;
    EQ_UNSIGNED #(.width(1)) u_eq_5144 (
        .y(_T_354),
        .a(isZeroB_PC),
        .b(1'h0)
    );
    wire _T_355;
    BITWISEAND #(.width(1)) bitwiseand_5145 (
        .y(_T_355),
        .a(_T_352),
        .b(_T_354)
    );
    wire _T_357;
    EQ_UNSIGNED #(.width(1)) u_eq_5146 (
        .y(_T_357),
        .a(_sign_PC__q),
        .b(1'h0)
    );
    wire _T_358;
    BITWISEAND #(.width(1)) bitwiseand_5147 (
        .y(_T_358),
        .a(_T_355),
        .b(_T_357)
    );
    wire _T_360;
    EQ_UNSIGNED #(.width(1)) u_eq_5148 (
        .y(_T_360),
        .a(isSpecialA_PC),
        .b(1'h0)
    );
    wire _T_362;
    EQ_UNSIGNED #(.width(1)) u_eq_5149 (
        .y(_T_362),
        .a(isSpecialB_PC),
        .b(1'h0)
    );
    wire _T_363;
    BITWISEAND #(.width(1)) bitwiseand_5150 (
        .y(_T_363),
        .a(_T_360),
        .b(_T_362)
    );
    wire _T_365;
    EQ_UNSIGNED #(.width(1)) u_eq_5151 (
        .y(_T_365),
        .a(isZeroA_PC),
        .b(1'h0)
    );
    wire _T_366;
    BITWISEAND #(.width(1)) bitwiseand_5152 (
        .y(_T_366),
        .a(_T_363),
        .b(_T_365)
    );
    wire _T_368;
    EQ_UNSIGNED #(.width(1)) u_eq_5153 (
        .y(_T_368),
        .a(isZeroB_PC),
        .b(1'h0)
    );
    wire _T_369;
    BITWISEAND #(.width(1)) bitwiseand_5154 (
        .y(_T_369),
        .a(_T_366),
        .b(_T_368)
    );
    wire normalCase_PC;
    MUX_UNSIGNED #(.width(1)) u_mux_5155 (
        .y(normalCase_PC),
        .sel(_sqrtOp_PC__q),
        .a(_T_358),
        .b(_T_369)
    );
    wire [14:0] _T_371;
    wire [13:0] _WTEMP_700;
    PAD_UNSIGNED #(.width(2), .n(14)) u_pad_5156 (
        .y(_WTEMP_700),
        .in(2'h2)
    );
    ADD_UNSIGNED #(.width(14)) u_add_5157 (
        .y(_T_371),
        .a(_exp_PC__q),
        .b(_WTEMP_700)
    );
    wire [13:0] expP2_PC;
    TAIL #(.width(15), .n(1)) tail_5158 (
        .y(expP2_PC),
        .in(_T_371)
    );
    wire _T_372;
    BITS #(.width(14), .high(0), .low(0)) bits_5159 (
        .y(_T_372),
        .in(_exp_PC__q)
    );
    wire [12:0] _T_373;
    BITS #(.width(14), .high(13), .low(1)) bits_5160 (
        .y(_T_373),
        .in(expP2_PC)
    );
    wire [13:0] _T_375;
    CAT #(.width_a(13), .width_b(1)) cat_5161 (
        .y(_T_375),
        .a(_T_373),
        .b(1'h0)
    );
    wire [12:0] _T_376;
    BITS #(.width(14), .high(13), .low(1)) bits_5162 (
        .y(_T_376),
        .in(_exp_PC__q)
    );
    wire [13:0] _T_378;
    CAT #(.width_a(13), .width_b(1)) cat_5163 (
        .y(_T_378),
        .a(_T_376),
        .b(1'h1)
    );
    wire [13:0] expP1_PC;
    MUX_UNSIGNED #(.width(14)) u_mux_5164 (
        .y(expP1_PC),
        .sel(_T_372),
        .a(_T_375),
        .b(_T_378)
    );
    wire roundingMode_near_even_PC;
    EQ_UNSIGNED #(.width(2)) u_eq_5165 (
        .y(roundingMode_near_even_PC),
        .a(_roundingMode_PC__q),
        .b(2'h0)
    );
    wire roundingMode_minMag_PC;
    EQ_UNSIGNED #(.width(2)) u_eq_5166 (
        .y(roundingMode_minMag_PC),
        .a(_roundingMode_PC__q),
        .b(2'h1)
    );
    wire roundingMode_min_PC;
    EQ_UNSIGNED #(.width(2)) u_eq_5167 (
        .y(roundingMode_min_PC),
        .a(_roundingMode_PC__q),
        .b(2'h2)
    );
    wire roundingMode_max_PC;
    EQ_UNSIGNED #(.width(2)) u_eq_5168 (
        .y(roundingMode_max_PC),
        .a(_roundingMode_PC__q),
        .b(2'h3)
    );
    wire roundMagUp_PC;
    MUX_UNSIGNED #(.width(1)) u_mux_5169 (
        .y(roundMagUp_PC),
        .sel(_sign_PC__q),
        .a(roundingMode_min_PC),
        .b(roundingMode_max_PC)
    );
    wire overflowY_roundMagUp_PC;
    BITWISEOR #(.width(1)) bitwiseor_5170 (
        .y(overflowY_roundMagUp_PC),
        .a(roundingMode_near_even_PC),
        .b(roundMagUp_PC)
    );
    wire _T_380;
    EQ_UNSIGNED #(.width(1)) u_eq_5171 (
        .y(_T_380),
        .a(roundMagUp_PC),
        .b(1'h0)
    );
    wire _T_382;
    EQ_UNSIGNED #(.width(1)) u_eq_5172 (
        .y(_T_382),
        .a(roundingMode_near_even_PC),
        .b(1'h0)
    );
    wire roundMagDown_PC;
    BITWISEAND #(.width(1)) bitwiseand_5173 (
        .y(roundMagDown_PC),
        .a(_T_380),
        .b(_T_382)
    );
    wire _T_384;
    EQ_UNSIGNED #(.width(1)) u_eq_5174 (
        .y(_T_384),
        .a(normalCase_PC),
        .b(1'h0)
    );
    wire valid_leaving_PC;
    BITWISEOR #(.width(1)) bitwiseor_5175 (
        .y(valid_leaving_PC),
        .a(_T_384),
        .b(cyc_E1)
    );
    wire _T_385;
    BITWISEAND #(.width(1)) bitwiseand_5176 (
        .y(_T_385),
        .a(_valid_PC__q),
        .b(valid_leaving_PC)
    );
    wire _T_387;
    EQ_UNSIGNED #(.width(1)) u_eq_5177 (
        .y(_T_387),
        .a(_valid_PC__q),
        .b(1'h0)
    );
    wire _T_388;
    BITWISEOR #(.width(1)) bitwiseor_5178 (
        .y(_T_388),
        .a(_T_387),
        .b(valid_leaving_PC)
    );
    wire _T_390;
    EQ_UNSIGNED #(.width(1)) u_eq_5179 (
        .y(_T_390),
        .a(_sqrtOp_PC__q),
        .b(1'h0)
    );
    wire _T_391;
    BITWISEAND #(.width(1)) bitwiseand_5180 (
        .y(_T_391),
        .a(leaving_PC),
        .b(_T_390)
    );
    wire _T_392;
    BITWISEAND #(.width(1)) bitwiseand_5181 (
        .y(_T_392),
        .a(leaving_PC),
        .b(_sqrtOp_PC__q)
    );
    wire _T_394;
    wire [2:0] _WTEMP_701;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_5182 (
        .y(_WTEMP_701),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(3)) u_neq_5183 (
        .y(_T_394),
        .a(_cycleNum_A__q),
        .b(_WTEMP_701)
    );
    wire _T_395;
    BITWISEOR #(.width(1)) bitwiseor_5184 (
        .y(_T_395),
        .a(entering_PA_normalCase),
        .b(_T_394)
    );
    wire [1:0] _T_398;
    wire [1:0] _WTEMP_702;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_5185 (
        .y(_WTEMP_702),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_5186 (
        .y(_T_398),
        .sel(cyc_A4_div),
        .a(2'h3),
        .b(_WTEMP_702)
    );
    wire [2:0] _T_401;
    wire [2:0] _WTEMP_703;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_5187 (
        .y(_WTEMP_703),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(3)) u_mux_5188 (
        .y(_T_401),
        .sel(cyc_A7_sqrt),
        .a(3'h6),
        .b(_WTEMP_703)
    );
    wire [2:0] _T_402;
    wire [2:0] _WTEMP_704;
    PAD_UNSIGNED #(.width(2), .n(3)) u_pad_5189 (
        .y(_WTEMP_704),
        .in(_T_398)
    );
    BITWISEOR #(.width(3)) bitwiseor_5190 (
        .y(_T_402),
        .a(_WTEMP_704),
        .b(_T_401)
    );
    wire _T_404;
    EQ_UNSIGNED #(.width(1)) u_eq_5191 (
        .y(_T_404),
        .a(entering_PA_normalCase),
        .b(1'h0)
    );
    wire [3:0] _T_406;
    wire [2:0] _WTEMP_705;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_5192 (
        .y(_WTEMP_705),
        .in(1'h1)
    );
    SUB_UNSIGNED #(.width(3)) u_sub_5193 (
        .y(_T_406),
        .a(_cycleNum_A__q),
        .b(_WTEMP_705)
    );
    wire [3:0] _T_407;
    ASUINT #(.width(4)) asuint_5194 (
        .y(_T_407),
        .in(_T_406)
    );
    wire [2:0] _T_408;
    TAIL #(.width(4), .n(1)) tail_5195 (
        .y(_T_408),
        .in(_T_407)
    );
    wire [2:0] _T_410;
    wire [2:0] _WTEMP_706;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_5196 (
        .y(_WTEMP_706),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(3)) u_mux_5197 (
        .y(_T_410),
        .sel(_T_404),
        .a(_T_408),
        .b(_WTEMP_706)
    );
    wire [2:0] _T_411;
    BITWISEOR #(.width(3)) bitwiseor_5198 (
        .y(_T_411),
        .a(_T_402),
        .b(_T_410)
    );
    wire cyc_A6_sqrt;
    EQ_UNSIGNED #(.width(3)) u_eq_5199 (
        .y(cyc_A6_sqrt),
        .a(_cycleNum_A__q),
        .b(3'h6)
    );
    wire cyc_A5_sqrt;
    EQ_UNSIGNED #(.width(3)) u_eq_5200 (
        .y(cyc_A5_sqrt),
        .a(_cycleNum_A__q),
        .b(3'h5)
    );
    wire cyc_A4_sqrt;
    EQ_UNSIGNED #(.width(3)) u_eq_5201 (
        .y(cyc_A4_sqrt),
        .a(_cycleNum_A__q),
        .b(3'h4)
    );
    wire cyc_A4;
    BITWISEOR #(.width(1)) bitwiseor_5202 (
        .y(cyc_A4),
        .a(cyc_A4_sqrt),
        .b(cyc_A4_div)
    );
    wire cyc_A3;
    wire [2:0] _WTEMP_707;
    PAD_UNSIGNED #(.width(2), .n(3)) u_pad_5203 (
        .y(_WTEMP_707),
        .in(2'h3)
    );
    EQ_UNSIGNED #(.width(3)) u_eq_5204 (
        .y(cyc_A3),
        .a(_cycleNum_A__q),
        .b(_WTEMP_707)
    );
    wire cyc_A2;
    wire [2:0] _WTEMP_708;
    PAD_UNSIGNED #(.width(2), .n(3)) u_pad_5205 (
        .y(_WTEMP_708),
        .in(2'h2)
    );
    EQ_UNSIGNED #(.width(3)) u_eq_5206 (
        .y(cyc_A2),
        .a(_cycleNum_A__q),
        .b(_WTEMP_708)
    );
    wire cyc_A1;
    wire [2:0] _WTEMP_709;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_5207 (
        .y(_WTEMP_709),
        .in(1'h1)
    );
    EQ_UNSIGNED #(.width(3)) u_eq_5208 (
        .y(cyc_A1),
        .a(_cycleNum_A__q),
        .b(_WTEMP_709)
    );
    wire _T_419;
    EQ_UNSIGNED #(.width(1)) u_eq_5209 (
        .y(_T_419),
        .a(_sqrtOp_PA__q),
        .b(1'h0)
    );
    wire cyc_A3_div;
    BITWISEAND #(.width(1)) bitwiseand_5210 (
        .y(cyc_A3_div),
        .a(cyc_A3),
        .b(_T_419)
    );
    wire _T_421;
    EQ_UNSIGNED #(.width(1)) u_eq_5211 (
        .y(_T_421),
        .a(_sqrtOp_PA__q),
        .b(1'h0)
    );
    wire cyc_A2_div;
    BITWISEAND #(.width(1)) bitwiseand_5212 (
        .y(cyc_A2_div),
        .a(cyc_A2),
        .b(_T_421)
    );
    wire _T_423;
    EQ_UNSIGNED #(.width(1)) u_eq_5213 (
        .y(_T_423),
        .a(_sqrtOp_PA__q),
        .b(1'h0)
    );
    wire cyc_A1_div;
    BITWISEAND #(.width(1)) bitwiseand_5214 (
        .y(cyc_A1_div),
        .a(cyc_A1),
        .b(_T_423)
    );
    wire cyc_A3_sqrt;
    BITWISEAND #(.width(1)) bitwiseand_5215 (
        .y(cyc_A3_sqrt),
        .a(cyc_A3),
        .b(_sqrtOp_PA__q)
    );
    wire cyc_A2_sqrt;
    BITWISEAND #(.width(1)) bitwiseand_5216 (
        .y(cyc_A2_sqrt),
        .a(cyc_A2),
        .b(_sqrtOp_PA__q)
    );
    wire cyc_A1_sqrt;
    BITWISEAND #(.width(1)) bitwiseand_5217 (
        .y(cyc_A1_sqrt),
        .a(cyc_A1),
        .b(_sqrtOp_PA__q)
    );
    wire _T_425;
    wire [3:0] _WTEMP_710;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_5218 (
        .y(_WTEMP_710),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_5219 (
        .y(_T_425),
        .a(_cycleNum_B__q),
        .b(_WTEMP_710)
    );
    wire _T_426;
    BITWISEOR #(.width(1)) bitwiseor_5220 (
        .y(_T_426),
        .a(cyc_A1),
        .b(_T_425)
    );
    wire [3:0] _T_429;
    wire [3:0] _WTEMP_711;
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_5221 (
        .y(_WTEMP_711),
        .in(3'h6)
    );
    MUX_UNSIGNED #(.width(4)) u_mux_5222 (
        .y(_T_429),
        .sel(_sqrtOp_PA__q),
        .a(4'hA),
        .b(_WTEMP_711)
    );
    wire [4:0] _T_431;
    wire [3:0] _WTEMP_712;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_5223 (
        .y(_WTEMP_712),
        .in(1'h1)
    );
    SUB_UNSIGNED #(.width(4)) u_sub_5224 (
        .y(_T_431),
        .a(_cycleNum_B__q),
        .b(_WTEMP_712)
    );
    wire [4:0] _T_432;
    ASUINT #(.width(5)) asuint_5225 (
        .y(_T_432),
        .in(_T_431)
    );
    wire [3:0] _T_433;
    TAIL #(.width(5), .n(1)) tail_5226 (
        .y(_T_433),
        .in(_T_432)
    );
    wire [3:0] _T_434;
    MUX_UNSIGNED #(.width(4)) u_mux_5227 (
        .y(_T_434),
        .sel(cyc_A1),
        .a(_T_429),
        .b(_T_433)
    );
    wire _T_436;
    EQ_UNSIGNED #(.width(4)) u_eq_5228 (
        .y(_T_436),
        .a(_cycleNum_B__q),
        .b(4'hA)
    );
    wire _T_438;
    EQ_UNSIGNED #(.width(4)) u_eq_5229 (
        .y(_T_438),
        .a(_cycleNum_B__q),
        .b(4'h9)
    );
    wire _T_440;
    EQ_UNSIGNED #(.width(4)) u_eq_5230 (
        .y(_T_440),
        .a(_cycleNum_B__q),
        .b(4'h8)
    );
    wire _T_442;
    wire [3:0] _WTEMP_713;
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_5231 (
        .y(_WTEMP_713),
        .in(3'h7)
    );
    EQ_UNSIGNED #(.width(4)) u_eq_5232 (
        .y(_T_442),
        .a(_cycleNum_B__q),
        .b(_WTEMP_713)
    );
    wire _T_444;
    wire [3:0] _WTEMP_714;
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_5233 (
        .y(_WTEMP_714),
        .in(3'h6)
    );
    EQ_UNSIGNED #(.width(4)) u_eq_5234 (
        .y(_T_444),
        .a(_cycleNum_B__q),
        .b(_WTEMP_714)
    );
    wire _T_446;
    wire [3:0] _WTEMP_715;
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_5235 (
        .y(_WTEMP_715),
        .in(3'h5)
    );
    EQ_UNSIGNED #(.width(4)) u_eq_5236 (
        .y(_T_446),
        .a(_cycleNum_B__q),
        .b(_WTEMP_715)
    );
    wire _T_448;
    wire [3:0] _WTEMP_716;
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_5237 (
        .y(_WTEMP_716),
        .in(3'h4)
    );
    EQ_UNSIGNED #(.width(4)) u_eq_5238 (
        .y(_T_448),
        .a(_cycleNum_B__q),
        .b(_WTEMP_716)
    );
    wire _T_450;
    wire [3:0] _WTEMP_717;
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_5239 (
        .y(_WTEMP_717),
        .in(2'h3)
    );
    EQ_UNSIGNED #(.width(4)) u_eq_5240 (
        .y(_T_450),
        .a(_cycleNum_B__q),
        .b(_WTEMP_717)
    );
    wire _T_452;
    wire [3:0] _WTEMP_718;
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_5241 (
        .y(_WTEMP_718),
        .in(2'h2)
    );
    EQ_UNSIGNED #(.width(4)) u_eq_5242 (
        .y(_T_452),
        .a(_cycleNum_B__q),
        .b(_WTEMP_718)
    );
    wire _T_454;
    wire [3:0] _WTEMP_719;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_5243 (
        .y(_WTEMP_719),
        .in(1'h1)
    );
    EQ_UNSIGNED #(.width(4)) u_eq_5244 (
        .y(_T_454),
        .a(_cycleNum_B__q),
        .b(_WTEMP_719)
    );
    wire _T_455;
    BITWISEAND #(.width(1)) bitwiseand_5245 (
        .y(_T_455),
        .a(cyc_B6),
        .b(_valid_PA__q)
    );
    wire _T_457;
    EQ_UNSIGNED #(.width(1)) u_eq_5246 (
        .y(_T_457),
        .a(_sqrtOp_PA__q),
        .b(1'h0)
    );
    wire _T_458;
    BITWISEAND #(.width(1)) bitwiseand_5247 (
        .y(_T_458),
        .a(_T_455),
        .b(_T_457)
    );
    wire _T_459;
    BITWISEAND #(.width(1)) bitwiseand_5248 (
        .y(_T_459),
        .a(cyc_B5),
        .b(_valid_PA__q)
    );
    wire _T_461;
    EQ_UNSIGNED #(.width(1)) u_eq_5249 (
        .y(_T_461),
        .a(_sqrtOp_PA__q),
        .b(1'h0)
    );
    wire _T_462;
    BITWISEAND #(.width(1)) bitwiseand_5250 (
        .y(_T_462),
        .a(_T_459),
        .b(_T_461)
    );
    wire _T_463;
    BITWISEAND #(.width(1)) bitwiseand_5251 (
        .y(_T_463),
        .a(cyc_B4),
        .b(_valid_PA__q)
    );
    wire _T_465;
    EQ_UNSIGNED #(.width(1)) u_eq_5252 (
        .y(_T_465),
        .a(_sqrtOp_PA__q),
        .b(1'h0)
    );
    wire _T_466;
    BITWISEAND #(.width(1)) bitwiseand_5253 (
        .y(_T_466),
        .a(_T_463),
        .b(_T_465)
    );
    wire _T_468;
    EQ_UNSIGNED #(.width(1)) u_eq_5254 (
        .y(_T_468),
        .a(_sqrtOp_PB__q),
        .b(1'h0)
    );
    wire _T_469;
    BITWISEAND #(.width(1)) bitwiseand_5255 (
        .y(_T_469),
        .a(cyc_B3),
        .b(_T_468)
    );
    wire _T_471;
    EQ_UNSIGNED #(.width(1)) u_eq_5256 (
        .y(_T_471),
        .a(_sqrtOp_PB__q),
        .b(1'h0)
    );
    wire _T_472;
    BITWISEAND #(.width(1)) bitwiseand_5257 (
        .y(_T_472),
        .a(cyc_B2),
        .b(_T_471)
    );
    wire _T_474;
    EQ_UNSIGNED #(.width(1)) u_eq_5258 (
        .y(_T_474),
        .a(_sqrtOp_PB__q),
        .b(1'h0)
    );
    wire _T_475;
    BITWISEAND #(.width(1)) bitwiseand_5259 (
        .y(_T_475),
        .a(cyc_B1),
        .b(_T_474)
    );
    wire _T_476;
    BITWISEAND #(.width(1)) bitwiseand_5260 (
        .y(_T_476),
        .a(cyc_B6),
        .b(_valid_PB__q)
    );
    wire _T_477;
    BITWISEAND #(.width(1)) bitwiseand_5261 (
        .y(_T_477),
        .a(_T_476),
        .b(_sqrtOp_PB__q)
    );
    wire _T_478;
    BITWISEAND #(.width(1)) bitwiseand_5262 (
        .y(_T_478),
        .a(cyc_B5),
        .b(_valid_PB__q)
    );
    wire _T_479;
    BITWISEAND #(.width(1)) bitwiseand_5263 (
        .y(_T_479),
        .a(_T_478),
        .b(_sqrtOp_PB__q)
    );
    wire _T_480;
    BITWISEAND #(.width(1)) bitwiseand_5264 (
        .y(_T_480),
        .a(cyc_B4),
        .b(_valid_PB__q)
    );
    wire _T_481;
    BITWISEAND #(.width(1)) bitwiseand_5265 (
        .y(_T_481),
        .a(_T_480),
        .b(_sqrtOp_PB__q)
    );
    wire _T_482;
    BITWISEAND #(.width(1)) bitwiseand_5266 (
        .y(_T_482),
        .a(cyc_B3),
        .b(_sqrtOp_PB__q)
    );
    wire _T_483;
    BITWISEAND #(.width(1)) bitwiseand_5267 (
        .y(_T_483),
        .a(cyc_B2),
        .b(_sqrtOp_PB__q)
    );
    wire _T_484;
    BITWISEAND #(.width(1)) bitwiseand_5268 (
        .y(_T_484),
        .a(cyc_B1),
        .b(_sqrtOp_PB__q)
    );
    wire _T_486;
    wire [2:0] _WTEMP_720;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_5269 (
        .y(_WTEMP_720),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(3)) u_neq_5270 (
        .y(_T_486),
        .a(_cycleNum_C__q),
        .b(_WTEMP_720)
    );
    wire _T_487;
    BITWISEOR #(.width(1)) bitwiseor_5271 (
        .y(_T_487),
        .a(cyc_B1),
        .b(_T_486)
    );
    wire [2:0] _T_490;
    MUX_UNSIGNED #(.width(3)) u_mux_5272 (
        .y(_T_490),
        .sel(_sqrtOp_PB__q),
        .a(3'h6),
        .b(3'h5)
    );
    wire [3:0] _T_492;
    wire [2:0] _WTEMP_721;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_5273 (
        .y(_WTEMP_721),
        .in(1'h1)
    );
    SUB_UNSIGNED #(.width(3)) u_sub_5274 (
        .y(_T_492),
        .a(_cycleNum_C__q),
        .b(_WTEMP_721)
    );
    wire [3:0] _T_493;
    ASUINT #(.width(4)) asuint_5275 (
        .y(_T_493),
        .in(_T_492)
    );
    wire [2:0] _T_494;
    TAIL #(.width(4), .n(1)) tail_5276 (
        .y(_T_494),
        .in(_T_493)
    );
    wire [2:0] _T_495;
    MUX_UNSIGNED #(.width(3)) u_mux_5277 (
        .y(_T_495),
        .sel(cyc_B1),
        .a(_T_490),
        .b(_T_494)
    );
    wire cyc_C6_sqrt;
    EQ_UNSIGNED #(.width(3)) u_eq_5278 (
        .y(cyc_C6_sqrt),
        .a(_cycleNum_C__q),
        .b(3'h6)
    );
    wire _T_498;
    EQ_UNSIGNED #(.width(3)) u_eq_5279 (
        .y(_T_498),
        .a(_cycleNum_C__q),
        .b(3'h5)
    );
    wire _T_500;
    EQ_UNSIGNED #(.width(3)) u_eq_5280 (
        .y(_T_500),
        .a(_cycleNum_C__q),
        .b(3'h4)
    );
    wire _T_502;
    wire [2:0] _WTEMP_722;
    PAD_UNSIGNED #(.width(2), .n(3)) u_pad_5281 (
        .y(_WTEMP_722),
        .in(2'h3)
    );
    EQ_UNSIGNED #(.width(3)) u_eq_5282 (
        .y(_T_502),
        .a(_cycleNum_C__q),
        .b(_WTEMP_722)
    );
    wire _T_504;
    wire [2:0] _WTEMP_723;
    PAD_UNSIGNED #(.width(2), .n(3)) u_pad_5283 (
        .y(_WTEMP_723),
        .in(2'h2)
    );
    EQ_UNSIGNED #(.width(3)) u_eq_5284 (
        .y(_T_504),
        .a(_cycleNum_C__q),
        .b(_WTEMP_723)
    );
    wire _T_506;
    wire [2:0] _WTEMP_724;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_5285 (
        .y(_WTEMP_724),
        .in(1'h1)
    );
    EQ_UNSIGNED #(.width(3)) u_eq_5286 (
        .y(_T_506),
        .a(_cycleNum_C__q),
        .b(_WTEMP_724)
    );
    wire _T_508;
    EQ_UNSIGNED #(.width(1)) u_eq_5287 (
        .y(_T_508),
        .a(_sqrtOp_PB__q),
        .b(1'h0)
    );
    wire cyc_C5_div;
    BITWISEAND #(.width(1)) bitwiseand_5288 (
        .y(cyc_C5_div),
        .a(cyc_C5),
        .b(_T_508)
    );
    wire _T_510;
    EQ_UNSIGNED #(.width(1)) u_eq_5289 (
        .y(_T_510),
        .a(_sqrtOp_PB__q),
        .b(1'h0)
    );
    wire cyc_C4_div;
    BITWISEAND #(.width(1)) bitwiseand_5290 (
        .y(cyc_C4_div),
        .a(cyc_C4),
        .b(_T_510)
    );
    wire _T_512;
    EQ_UNSIGNED #(.width(1)) u_eq_5291 (
        .y(_T_512),
        .a(_sqrtOp_PB__q),
        .b(1'h0)
    );
    wire cyc_C3_div;
    BITWISEAND #(.width(1)) bitwiseand_5292 (
        .y(cyc_C3_div),
        .a(cyc_C3),
        .b(_T_512)
    );
    wire _T_514;
    EQ_UNSIGNED #(.width(1)) u_eq_5293 (
        .y(_T_514),
        .a(_sqrtOp_PC__q),
        .b(1'h0)
    );
    wire cyc_C2_div;
    BITWISEAND #(.width(1)) bitwiseand_5294 (
        .y(cyc_C2_div),
        .a(cyc_C2),
        .b(_T_514)
    );
    wire _T_516;
    EQ_UNSIGNED #(.width(1)) u_eq_5295 (
        .y(_T_516),
        .a(_sqrtOp_PC__q),
        .b(1'h0)
    );
    wire cyc_C1_div;
    BITWISEAND #(.width(1)) bitwiseand_5296 (
        .y(cyc_C1_div),
        .a(cyc_C1),
        .b(_T_516)
    );
    wire cyc_C5_sqrt;
    BITWISEAND #(.width(1)) bitwiseand_5297 (
        .y(cyc_C5_sqrt),
        .a(cyc_C5),
        .b(_sqrtOp_PB__q)
    );
    wire cyc_C4_sqrt;
    BITWISEAND #(.width(1)) bitwiseand_5298 (
        .y(cyc_C4_sqrt),
        .a(cyc_C4),
        .b(_sqrtOp_PB__q)
    );
    wire cyc_C3_sqrt;
    BITWISEAND #(.width(1)) bitwiseand_5299 (
        .y(cyc_C3_sqrt),
        .a(cyc_C3),
        .b(_sqrtOp_PB__q)
    );
    wire cyc_C2_sqrt;
    BITWISEAND #(.width(1)) bitwiseand_5300 (
        .y(cyc_C2_sqrt),
        .a(cyc_C2),
        .b(_sqrtOp_PC__q)
    );
    wire cyc_C1_sqrt;
    BITWISEAND #(.width(1)) bitwiseand_5301 (
        .y(cyc_C1_sqrt),
        .a(cyc_C1),
        .b(_sqrtOp_PC__q)
    );
    wire _T_518;
    wire [2:0] _WTEMP_725;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_5302 (
        .y(_WTEMP_725),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(3)) u_neq_5303 (
        .y(_T_518),
        .a(_cycleNum_E__q),
        .b(_WTEMP_725)
    );
    wire _T_519;
    BITWISEOR #(.width(1)) bitwiseor_5304 (
        .y(_T_519),
        .a(cyc_C1),
        .b(_T_518)
    );
    wire [3:0] _T_522;
    wire [2:0] _WTEMP_726;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_5305 (
        .y(_WTEMP_726),
        .in(1'h1)
    );
    SUB_UNSIGNED #(.width(3)) u_sub_5306 (
        .y(_T_522),
        .a(_cycleNum_E__q),
        .b(_WTEMP_726)
    );
    wire [3:0] _T_523;
    ASUINT #(.width(4)) asuint_5307 (
        .y(_T_523),
        .in(_T_522)
    );
    wire [2:0] _T_524;
    TAIL #(.width(4), .n(1)) tail_5308 (
        .y(_T_524),
        .in(_T_523)
    );
    wire [2:0] _T_525;
    MUX_UNSIGNED #(.width(3)) u_mux_5309 (
        .y(_T_525),
        .sel(cyc_C1),
        .a(3'h4),
        .b(_T_524)
    );
    wire _T_527;
    EQ_UNSIGNED #(.width(3)) u_eq_5310 (
        .y(_T_527),
        .a(_cycleNum_E__q),
        .b(3'h4)
    );
    wire _T_529;
    wire [2:0] _WTEMP_727;
    PAD_UNSIGNED #(.width(2), .n(3)) u_pad_5311 (
        .y(_WTEMP_727),
        .in(2'h3)
    );
    EQ_UNSIGNED #(.width(3)) u_eq_5312 (
        .y(_T_529),
        .a(_cycleNum_E__q),
        .b(_WTEMP_727)
    );
    wire _T_531;
    wire [2:0] _WTEMP_728;
    PAD_UNSIGNED #(.width(2), .n(3)) u_pad_5313 (
        .y(_WTEMP_728),
        .in(2'h2)
    );
    EQ_UNSIGNED #(.width(3)) u_eq_5314 (
        .y(_T_531),
        .a(_cycleNum_E__q),
        .b(_WTEMP_728)
    );
    wire _T_533;
    wire [2:0] _WTEMP_729;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_5315 (
        .y(_WTEMP_729),
        .in(1'h1)
    );
    EQ_UNSIGNED #(.width(3)) u_eq_5316 (
        .y(_T_533),
        .a(_cycleNum_E__q),
        .b(_WTEMP_729)
    );
    wire _T_535;
    EQ_UNSIGNED #(.width(1)) u_eq_5317 (
        .y(_T_535),
        .a(_sqrtOp_PC__q),
        .b(1'h0)
    );
    wire cyc_E4_div;
    BITWISEAND #(.width(1)) bitwiseand_5318 (
        .y(cyc_E4_div),
        .a(cyc_E4),
        .b(_T_535)
    );
    wire _T_537;
    EQ_UNSIGNED #(.width(1)) u_eq_5319 (
        .y(_T_537),
        .a(_sqrtOp_PC__q),
        .b(1'h0)
    );
    wire cyc_E3_div;
    BITWISEAND #(.width(1)) bitwiseand_5320 (
        .y(cyc_E3_div),
        .a(cyc_E3),
        .b(_T_537)
    );
    wire _T_539;
    EQ_UNSIGNED #(.width(1)) u_eq_5321 (
        .y(_T_539),
        .a(_sqrtOp_PC__q),
        .b(1'h0)
    );
    wire cyc_E2_div;
    BITWISEAND #(.width(1)) bitwiseand_5322 (
        .y(cyc_E2_div),
        .a(cyc_E2),
        .b(_T_539)
    );
    wire _T_541;
    EQ_UNSIGNED #(.width(1)) u_eq_5323 (
        .y(_T_541),
        .a(_sqrtOp_PC__q),
        .b(1'h0)
    );
    wire cyc_E1_div;
    BITWISEAND #(.width(1)) bitwiseand_5324 (
        .y(cyc_E1_div),
        .a(cyc_E1),
        .b(_T_541)
    );
    wire cyc_E4_sqrt;
    BITWISEAND #(.width(1)) bitwiseand_5325 (
        .y(cyc_E4_sqrt),
        .a(cyc_E4),
        .b(_sqrtOp_PC__q)
    );
    wire cyc_E3_sqrt;
    BITWISEAND #(.width(1)) bitwiseand_5326 (
        .y(cyc_E3_sqrt),
        .a(cyc_E3),
        .b(_sqrtOp_PC__q)
    );
    wire cyc_E2_sqrt;
    BITWISEAND #(.width(1)) bitwiseand_5327 (
        .y(cyc_E2_sqrt),
        .a(cyc_E2),
        .b(_sqrtOp_PC__q)
    );
    wire cyc_E1_sqrt;
    BITWISEAND #(.width(1)) bitwiseand_5328 (
        .y(cyc_E1_sqrt),
        .a(cyc_E1),
        .b(_sqrtOp_PC__q)
    );
    wire [51:0] zFractB_A4_div;
    wire [51:0] _WTEMP_730;
    PAD_UNSIGNED #(.width(1), .n(52)) u_pad_5329 (
        .y(_WTEMP_730),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(52)) u_mux_5330 (
        .y(zFractB_A4_div),
        .sel(cyc_A4_div),
        .a(fractB_S),
        .b(_WTEMP_730)
    );
    wire [2:0] _T_543;
    BITS #(.width(52), .high(51), .low(49)) bits_5331 (
        .y(_T_543),
        .in(fractB_S)
    );
    wire _T_545;
    wire [2:0] _WTEMP_731;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_5332 (
        .y(_WTEMP_731),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(3)) u_eq_5333 (
        .y(_T_545),
        .a(_T_543),
        .b(_WTEMP_731)
    );
    wire zLinPiece_0_A4_div;
    BITWISEAND #(.width(1)) bitwiseand_5334 (
        .y(zLinPiece_0_A4_div),
        .a(cyc_A4_div),
        .b(_T_545)
    );
    wire [2:0] _T_546;
    BITS #(.width(52), .high(51), .low(49)) bits_5335 (
        .y(_T_546),
        .in(fractB_S)
    );
    wire _T_548;
    wire [2:0] _WTEMP_732;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_5336 (
        .y(_WTEMP_732),
        .in(1'h1)
    );
    EQ_UNSIGNED #(.width(3)) u_eq_5337 (
        .y(_T_548),
        .a(_T_546),
        .b(_WTEMP_732)
    );
    wire zLinPiece_1_A4_div;
    BITWISEAND #(.width(1)) bitwiseand_5338 (
        .y(zLinPiece_1_A4_div),
        .a(cyc_A4_div),
        .b(_T_548)
    );
    wire [2:0] _T_549;
    BITS #(.width(52), .high(51), .low(49)) bits_5339 (
        .y(_T_549),
        .in(fractB_S)
    );
    wire _T_551;
    wire [2:0] _WTEMP_733;
    PAD_UNSIGNED #(.width(2), .n(3)) u_pad_5340 (
        .y(_WTEMP_733),
        .in(2'h2)
    );
    EQ_UNSIGNED #(.width(3)) u_eq_5341 (
        .y(_T_551),
        .a(_T_549),
        .b(_WTEMP_733)
    );
    wire zLinPiece_2_A4_div;
    BITWISEAND #(.width(1)) bitwiseand_5342 (
        .y(zLinPiece_2_A4_div),
        .a(cyc_A4_div),
        .b(_T_551)
    );
    wire [2:0] _T_552;
    BITS #(.width(52), .high(51), .low(49)) bits_5343 (
        .y(_T_552),
        .in(fractB_S)
    );
    wire _T_554;
    wire [2:0] _WTEMP_734;
    PAD_UNSIGNED #(.width(2), .n(3)) u_pad_5344 (
        .y(_WTEMP_734),
        .in(2'h3)
    );
    EQ_UNSIGNED #(.width(3)) u_eq_5345 (
        .y(_T_554),
        .a(_T_552),
        .b(_WTEMP_734)
    );
    wire zLinPiece_3_A4_div;
    BITWISEAND #(.width(1)) bitwiseand_5346 (
        .y(zLinPiece_3_A4_div),
        .a(cyc_A4_div),
        .b(_T_554)
    );
    wire [2:0] _T_555;
    BITS #(.width(52), .high(51), .low(49)) bits_5347 (
        .y(_T_555),
        .in(fractB_S)
    );
    wire _T_557;
    EQ_UNSIGNED #(.width(3)) u_eq_5348 (
        .y(_T_557),
        .a(_T_555),
        .b(3'h4)
    );
    wire zLinPiece_4_A4_div;
    BITWISEAND #(.width(1)) bitwiseand_5349 (
        .y(zLinPiece_4_A4_div),
        .a(cyc_A4_div),
        .b(_T_557)
    );
    wire [2:0] _T_558;
    BITS #(.width(52), .high(51), .low(49)) bits_5350 (
        .y(_T_558),
        .in(fractB_S)
    );
    wire _T_560;
    EQ_UNSIGNED #(.width(3)) u_eq_5351 (
        .y(_T_560),
        .a(_T_558),
        .b(3'h5)
    );
    wire zLinPiece_5_A4_div;
    BITWISEAND #(.width(1)) bitwiseand_5352 (
        .y(zLinPiece_5_A4_div),
        .a(cyc_A4_div),
        .b(_T_560)
    );
    wire [2:0] _T_561;
    BITS #(.width(52), .high(51), .low(49)) bits_5353 (
        .y(_T_561),
        .in(fractB_S)
    );
    wire _T_563;
    EQ_UNSIGNED #(.width(3)) u_eq_5354 (
        .y(_T_563),
        .a(_T_561),
        .b(3'h6)
    );
    wire zLinPiece_6_A4_div;
    BITWISEAND #(.width(1)) bitwiseand_5355 (
        .y(zLinPiece_6_A4_div),
        .a(cyc_A4_div),
        .b(_T_563)
    );
    wire [2:0] _T_564;
    BITS #(.width(52), .high(51), .low(49)) bits_5356 (
        .y(_T_564),
        .in(fractB_S)
    );
    wire _T_566;
    EQ_UNSIGNED #(.width(3)) u_eq_5357 (
        .y(_T_566),
        .a(_T_564),
        .b(3'h7)
    );
    wire zLinPiece_7_A4_div;
    BITWISEAND #(.width(1)) bitwiseand_5358 (
        .y(zLinPiece_7_A4_div),
        .a(cyc_A4_div),
        .b(_T_566)
    );
    wire [8:0] _T_569;
    wire [8:0] _WTEMP_735;
    PAD_UNSIGNED #(.width(1), .n(9)) u_pad_5359 (
        .y(_WTEMP_735),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(9)) u_mux_5360 (
        .y(_T_569),
        .sel(zLinPiece_0_A4_div),
        .a(9'h1C7),
        .b(_WTEMP_735)
    );
    wire [8:0] _T_572;
    wire [8:0] _WTEMP_736;
    PAD_UNSIGNED #(.width(1), .n(9)) u_pad_5361 (
        .y(_WTEMP_736),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(9)) u_mux_5362 (
        .y(_T_572),
        .sel(zLinPiece_1_A4_div),
        .a(9'h16C),
        .b(_WTEMP_736)
    );
    wire [8:0] _T_573;
    BITWISEOR #(.width(9)) bitwiseor_5363 (
        .y(_T_573),
        .a(_T_569),
        .b(_T_572)
    );
    wire [8:0] _T_576;
    wire [8:0] _WTEMP_737;
    PAD_UNSIGNED #(.width(1), .n(9)) u_pad_5364 (
        .y(_WTEMP_737),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(9)) u_mux_5365 (
        .y(_T_576),
        .sel(zLinPiece_2_A4_div),
        .a(9'h12A),
        .b(_WTEMP_737)
    );
    wire [8:0] _T_577;
    BITWISEOR #(.width(9)) bitwiseor_5366 (
        .y(_T_577),
        .a(_T_573),
        .b(_T_576)
    );
    wire [8:0] _T_580;
    wire [8:0] _WTEMP_738;
    PAD_UNSIGNED #(.width(1), .n(9)) u_pad_5367 (
        .y(_WTEMP_738),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(9)) u_mux_5368 (
        .y(_T_580),
        .sel(zLinPiece_3_A4_div),
        .a(9'hF8),
        .b(_WTEMP_738)
    );
    wire [8:0] _T_581;
    BITWISEOR #(.width(9)) bitwiseor_5369 (
        .y(_T_581),
        .a(_T_577),
        .b(_T_580)
    );
    wire [8:0] _T_584;
    wire [8:0] _WTEMP_739;
    PAD_UNSIGNED #(.width(1), .n(9)) u_pad_5370 (
        .y(_WTEMP_739),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(9)) u_mux_5371 (
        .y(_T_584),
        .sel(zLinPiece_4_A4_div),
        .a(9'hD2),
        .b(_WTEMP_739)
    );
    wire [8:0] _T_585;
    BITWISEOR #(.width(9)) bitwiseor_5372 (
        .y(_T_585),
        .a(_T_581),
        .b(_T_584)
    );
    wire [8:0] _T_588;
    wire [8:0] _WTEMP_740;
    PAD_UNSIGNED #(.width(1), .n(9)) u_pad_5373 (
        .y(_WTEMP_740),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(9)) u_mux_5374 (
        .y(_T_588),
        .sel(zLinPiece_5_A4_div),
        .a(9'hB4),
        .b(_WTEMP_740)
    );
    wire [8:0] _T_589;
    BITWISEOR #(.width(9)) bitwiseor_5375 (
        .y(_T_589),
        .a(_T_585),
        .b(_T_588)
    );
    wire [8:0] _T_592;
    wire [8:0] _WTEMP_741;
    PAD_UNSIGNED #(.width(1), .n(9)) u_pad_5376 (
        .y(_WTEMP_741),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(9)) u_mux_5377 (
        .y(_T_592),
        .sel(zLinPiece_6_A4_div),
        .a(9'h9C),
        .b(_WTEMP_741)
    );
    wire [8:0] _T_593;
    BITWISEOR #(.width(9)) bitwiseor_5378 (
        .y(_T_593),
        .a(_T_589),
        .b(_T_592)
    );
    wire [8:0] _T_596;
    wire [8:0] _WTEMP_742;
    PAD_UNSIGNED #(.width(1), .n(9)) u_pad_5379 (
        .y(_WTEMP_742),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(9)) u_mux_5380 (
        .y(_T_596),
        .sel(zLinPiece_7_A4_div),
        .a(9'h89),
        .b(_WTEMP_742)
    );
    wire [8:0] zK1_A4_div;
    BITWISEOR #(.width(9)) bitwiseor_5381 (
        .y(zK1_A4_div),
        .a(_T_593),
        .b(_T_596)
    );
    wire [11:0] _T_598;
    assign _T_598 = 12'h1C;
    wire [11:0] _T_600;
    wire [11:0] _WTEMP_743;
    PAD_UNSIGNED #(.width(1), .n(12)) u_pad_5382 (
        .y(_WTEMP_743),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(12)) u_mux_5383 (
        .y(_T_600),
        .sel(zLinPiece_0_A4_div),
        .a(_T_598),
        .b(_WTEMP_743)
    );
    wire [11:0] _T_602;
    assign _T_602 = 12'h3A2;
    wire [11:0] _T_604;
    wire [11:0] _WTEMP_744;
    PAD_UNSIGNED #(.width(1), .n(12)) u_pad_5384 (
        .y(_WTEMP_744),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(12)) u_mux_5385 (
        .y(_T_604),
        .sel(zLinPiece_1_A4_div),
        .a(_T_602),
        .b(_WTEMP_744)
    );
    wire [11:0] _T_605;
    BITWISEOR #(.width(12)) bitwiseor_5386 (
        .y(_T_605),
        .a(_T_600),
        .b(_T_604)
    );
    wire [11:0] _T_607;
    assign _T_607 = 12'h675;
    wire [11:0] _T_609;
    wire [11:0] _WTEMP_745;
    PAD_UNSIGNED #(.width(1), .n(12)) u_pad_5387 (
        .y(_WTEMP_745),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(12)) u_mux_5388 (
        .y(_T_609),
        .sel(zLinPiece_2_A4_div),
        .a(_T_607),
        .b(_WTEMP_745)
    );
    wire [11:0] _T_610;
    BITWISEOR #(.width(12)) bitwiseor_5389 (
        .y(_T_610),
        .a(_T_605),
        .b(_T_609)
    );
    wire [11:0] _T_612;
    assign _T_612 = 12'h8C6;
    wire [11:0] _T_614;
    wire [11:0] _WTEMP_746;
    PAD_UNSIGNED #(.width(1), .n(12)) u_pad_5390 (
        .y(_WTEMP_746),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(12)) u_mux_5391 (
        .y(_T_614),
        .sel(zLinPiece_3_A4_div),
        .a(_T_612),
        .b(_WTEMP_746)
    );
    wire [11:0] _T_615;
    BITWISEOR #(.width(12)) bitwiseor_5392 (
        .y(_T_615),
        .a(_T_610),
        .b(_T_614)
    );
    wire [11:0] _T_617;
    assign _T_617 = 12'hAB4;
    wire [11:0] _T_619;
    wire [11:0] _WTEMP_747;
    PAD_UNSIGNED #(.width(1), .n(12)) u_pad_5393 (
        .y(_WTEMP_747),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(12)) u_mux_5394 (
        .y(_T_619),
        .sel(zLinPiece_4_A4_div),
        .a(_T_617),
        .b(_WTEMP_747)
    );
    wire [11:0] _T_620;
    BITWISEOR #(.width(12)) bitwiseor_5395 (
        .y(_T_620),
        .a(_T_615),
        .b(_T_619)
    );
    wire [11:0] _T_622;
    assign _T_622 = 12'hC56;
    wire [11:0] _T_624;
    wire [11:0] _WTEMP_748;
    PAD_UNSIGNED #(.width(1), .n(12)) u_pad_5396 (
        .y(_WTEMP_748),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(12)) u_mux_5397 (
        .y(_T_624),
        .sel(zLinPiece_5_A4_div),
        .a(_T_622),
        .b(_WTEMP_748)
    );
    wire [11:0] _T_625;
    BITWISEOR #(.width(12)) bitwiseor_5398 (
        .y(_T_625),
        .a(_T_620),
        .b(_T_624)
    );
    wire [11:0] _T_627;
    assign _T_627 = 12'hDBD;
    wire [11:0] _T_629;
    wire [11:0] _WTEMP_749;
    PAD_UNSIGNED #(.width(1), .n(12)) u_pad_5399 (
        .y(_WTEMP_749),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(12)) u_mux_5400 (
        .y(_T_629),
        .sel(zLinPiece_6_A4_div),
        .a(_T_627),
        .b(_WTEMP_749)
    );
    wire [11:0] _T_630;
    BITWISEOR #(.width(12)) bitwiseor_5401 (
        .y(_T_630),
        .a(_T_625),
        .b(_T_629)
    );
    wire [11:0] _T_632;
    assign _T_632 = 12'hEF4;
    wire [11:0] _T_634;
    wire [11:0] _WTEMP_750;
    PAD_UNSIGNED #(.width(1), .n(12)) u_pad_5402 (
        .y(_WTEMP_750),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(12)) u_mux_5403 (
        .y(_T_634),
        .sel(zLinPiece_7_A4_div),
        .a(_T_632),
        .b(_WTEMP_750)
    );
    wire [11:0] zComplFractK0_A4_div;
    BITWISEOR #(.width(12)) bitwiseor_5404 (
        .y(zComplFractK0_A4_div),
        .a(_T_630),
        .b(_T_634)
    );
    wire [51:0] zFractB_A7_sqrt;
    wire [51:0] _WTEMP_751;
    PAD_UNSIGNED #(.width(1), .n(52)) u_pad_5405 (
        .y(_WTEMP_751),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(52)) u_mux_5406 (
        .y(zFractB_A7_sqrt),
        .sel(cyc_A7_sqrt),
        .a(fractB_S),
        .b(_WTEMP_751)
    );
    wire _T_636;
    BITS #(.width(12), .high(0), .low(0)) bits_5407 (
        .y(_T_636),
        .in(expB_S)
    );
    wire _T_638;
    EQ_UNSIGNED #(.width(1)) u_eq_5408 (
        .y(_T_638),
        .a(_T_636),
        .b(1'h0)
    );
    wire _T_639;
    BITWISEAND #(.width(1)) bitwiseand_5409 (
        .y(_T_639),
        .a(cyc_A7_sqrt),
        .b(_T_638)
    );
    wire _T_640;
    BITS #(.width(52), .high(51), .low(51)) bits_5410 (
        .y(_T_640),
        .in(fractB_S)
    );
    wire _T_642;
    EQ_UNSIGNED #(.width(1)) u_eq_5411 (
        .y(_T_642),
        .a(_T_640),
        .b(1'h0)
    );
    wire zQuadPiece_0_A7_sqrt;
    BITWISEAND #(.width(1)) bitwiseand_5412 (
        .y(zQuadPiece_0_A7_sqrt),
        .a(_T_639),
        .b(_T_642)
    );
    wire _T_643;
    BITS #(.width(12), .high(0), .low(0)) bits_5413 (
        .y(_T_643),
        .in(expB_S)
    );
    wire _T_645;
    EQ_UNSIGNED #(.width(1)) u_eq_5414 (
        .y(_T_645),
        .a(_T_643),
        .b(1'h0)
    );
    wire _T_646;
    BITWISEAND #(.width(1)) bitwiseand_5415 (
        .y(_T_646),
        .a(cyc_A7_sqrt),
        .b(_T_645)
    );
    wire _T_647;
    BITS #(.width(52), .high(51), .low(51)) bits_5416 (
        .y(_T_647),
        .in(fractB_S)
    );
    wire zQuadPiece_1_A7_sqrt;
    BITWISEAND #(.width(1)) bitwiseand_5417 (
        .y(zQuadPiece_1_A7_sqrt),
        .a(_T_646),
        .b(_T_647)
    );
    wire _T_648;
    BITS #(.width(12), .high(0), .low(0)) bits_5418 (
        .y(_T_648),
        .in(expB_S)
    );
    wire _T_649;
    BITWISEAND #(.width(1)) bitwiseand_5419 (
        .y(_T_649),
        .a(cyc_A7_sqrt),
        .b(_T_648)
    );
    wire _T_650;
    BITS #(.width(52), .high(51), .low(51)) bits_5420 (
        .y(_T_650),
        .in(fractB_S)
    );
    wire _T_652;
    EQ_UNSIGNED #(.width(1)) u_eq_5421 (
        .y(_T_652),
        .a(_T_650),
        .b(1'h0)
    );
    wire zQuadPiece_2_A7_sqrt;
    BITWISEAND #(.width(1)) bitwiseand_5422 (
        .y(zQuadPiece_2_A7_sqrt),
        .a(_T_649),
        .b(_T_652)
    );
    wire _T_653;
    BITS #(.width(12), .high(0), .low(0)) bits_5423 (
        .y(_T_653),
        .in(expB_S)
    );
    wire _T_654;
    BITWISEAND #(.width(1)) bitwiseand_5424 (
        .y(_T_654),
        .a(cyc_A7_sqrt),
        .b(_T_653)
    );
    wire _T_655;
    BITS #(.width(52), .high(51), .low(51)) bits_5425 (
        .y(_T_655),
        .in(fractB_S)
    );
    wire zQuadPiece_3_A7_sqrt;
    BITWISEAND #(.width(1)) bitwiseand_5426 (
        .y(zQuadPiece_3_A7_sqrt),
        .a(_T_654),
        .b(_T_655)
    );
    wire [8:0] _T_658;
    wire [8:0] _WTEMP_752;
    PAD_UNSIGNED #(.width(1), .n(9)) u_pad_5427 (
        .y(_WTEMP_752),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(9)) u_mux_5428 (
        .y(_T_658),
        .sel(zQuadPiece_0_A7_sqrt),
        .a(9'h1C8),
        .b(_WTEMP_752)
    );
    wire [8:0] _T_661;
    wire [8:0] _WTEMP_753;
    PAD_UNSIGNED #(.width(1), .n(9)) u_pad_5429 (
        .y(_WTEMP_753),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(9)) u_mux_5430 (
        .y(_T_661),
        .sel(zQuadPiece_1_A7_sqrt),
        .a(9'hC1),
        .b(_WTEMP_753)
    );
    wire [8:0] _T_662;
    BITWISEOR #(.width(9)) bitwiseor_5431 (
        .y(_T_662),
        .a(_T_658),
        .b(_T_661)
    );
    wire [8:0] _T_665;
    wire [8:0] _WTEMP_754;
    PAD_UNSIGNED #(.width(1), .n(9)) u_pad_5432 (
        .y(_WTEMP_754),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(9)) u_mux_5433 (
        .y(_T_665),
        .sel(zQuadPiece_2_A7_sqrt),
        .a(9'h143),
        .b(_WTEMP_754)
    );
    wire [8:0] _T_666;
    BITWISEOR #(.width(9)) bitwiseor_5434 (
        .y(_T_666),
        .a(_T_662),
        .b(_T_665)
    );
    wire [8:0] _T_669;
    wire [8:0] _WTEMP_755;
    PAD_UNSIGNED #(.width(1), .n(9)) u_pad_5435 (
        .y(_WTEMP_755),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(9)) u_mux_5436 (
        .y(_T_669),
        .sel(zQuadPiece_3_A7_sqrt),
        .a(9'h89),
        .b(_WTEMP_755)
    );
    wire [8:0] zK2_A7_sqrt;
    BITWISEOR #(.width(9)) bitwiseor_5437 (
        .y(zK2_A7_sqrt),
        .a(_T_666),
        .b(_T_669)
    );
    wire [9:0] _T_671;
    assign _T_671 = 10'h2F;
    wire [9:0] _T_673;
    wire [9:0] _WTEMP_756;
    PAD_UNSIGNED #(.width(1), .n(10)) u_pad_5438 (
        .y(_WTEMP_756),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(10)) u_mux_5439 (
        .y(_T_673),
        .sel(zQuadPiece_0_A7_sqrt),
        .a(_T_671),
        .b(_WTEMP_756)
    );
    wire [9:0] _T_675;
    assign _T_675 = 10'h1DF;
    wire [9:0] _T_677;
    wire [9:0] _WTEMP_757;
    PAD_UNSIGNED #(.width(1), .n(10)) u_pad_5440 (
        .y(_WTEMP_757),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(10)) u_mux_5441 (
        .y(_T_677),
        .sel(zQuadPiece_1_A7_sqrt),
        .a(_T_675),
        .b(_WTEMP_757)
    );
    wire [9:0] _T_678;
    BITWISEOR #(.width(10)) bitwiseor_5442 (
        .y(_T_678),
        .a(_T_673),
        .b(_T_677)
    );
    wire [9:0] _T_680;
    assign _T_680 = 10'h14D;
    wire [9:0] _T_682;
    wire [9:0] _WTEMP_758;
    PAD_UNSIGNED #(.width(1), .n(10)) u_pad_5443 (
        .y(_WTEMP_758),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(10)) u_mux_5444 (
        .y(_T_682),
        .sel(zQuadPiece_2_A7_sqrt),
        .a(_T_680),
        .b(_WTEMP_758)
    );
    wire [9:0] _T_683;
    BITWISEOR #(.width(10)) bitwiseor_5445 (
        .y(_T_683),
        .a(_T_678),
        .b(_T_682)
    );
    wire [9:0] _T_685;
    assign _T_685 = 10'h27E;
    wire [9:0] _T_687;
    wire [9:0] _WTEMP_759;
    PAD_UNSIGNED #(.width(1), .n(10)) u_pad_5446 (
        .y(_WTEMP_759),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(10)) u_mux_5447 (
        .y(_T_687),
        .sel(zQuadPiece_3_A7_sqrt),
        .a(_T_685),
        .b(_WTEMP_759)
    );
    wire [9:0] zComplK1_A7_sqrt;
    BITWISEOR #(.width(10)) bitwiseor_5448 (
        .y(zComplK1_A7_sqrt),
        .a(_T_683),
        .b(_T_687)
    );
    wire _T_688;
    BITS #(.width(14), .high(0), .low(0)) bits_5449 (
        .y(_T_688),
        .in(_exp_PA__q)
    );
    wire _T_690;
    EQ_UNSIGNED #(.width(1)) u_eq_5450 (
        .y(_T_690),
        .a(_T_688),
        .b(1'h0)
    );
    wire _T_691;
    BITWISEAND #(.width(1)) bitwiseand_5451 (
        .y(_T_691),
        .a(cyc_A6_sqrt),
        .b(_T_690)
    );
    wire _T_692;
    BITS #(.width(53), .high(51), .low(51)) bits_5452 (
        .y(_T_692),
        .in(sigB_PA)
    );
    wire _T_694;
    EQ_UNSIGNED #(.width(1)) u_eq_5453 (
        .y(_T_694),
        .a(_T_692),
        .b(1'h0)
    );
    wire zQuadPiece_0_A6_sqrt;
    BITWISEAND #(.width(1)) bitwiseand_5454 (
        .y(zQuadPiece_0_A6_sqrt),
        .a(_T_691),
        .b(_T_694)
    );
    wire _T_695;
    BITS #(.width(14), .high(0), .low(0)) bits_5455 (
        .y(_T_695),
        .in(_exp_PA__q)
    );
    wire _T_697;
    EQ_UNSIGNED #(.width(1)) u_eq_5456 (
        .y(_T_697),
        .a(_T_695),
        .b(1'h0)
    );
    wire _T_698;
    BITWISEAND #(.width(1)) bitwiseand_5457 (
        .y(_T_698),
        .a(cyc_A6_sqrt),
        .b(_T_697)
    );
    wire _T_699;
    BITS #(.width(53), .high(51), .low(51)) bits_5458 (
        .y(_T_699),
        .in(sigB_PA)
    );
    wire zQuadPiece_1_A6_sqrt;
    BITWISEAND #(.width(1)) bitwiseand_5459 (
        .y(zQuadPiece_1_A6_sqrt),
        .a(_T_698),
        .b(_T_699)
    );
    wire _T_700;
    BITS #(.width(14), .high(0), .low(0)) bits_5460 (
        .y(_T_700),
        .in(_exp_PA__q)
    );
    wire _T_701;
    BITWISEAND #(.width(1)) bitwiseand_5461 (
        .y(_T_701),
        .a(cyc_A6_sqrt),
        .b(_T_700)
    );
    wire _T_702;
    BITS #(.width(53), .high(51), .low(51)) bits_5462 (
        .y(_T_702),
        .in(sigB_PA)
    );
    wire _T_704;
    EQ_UNSIGNED #(.width(1)) u_eq_5463 (
        .y(_T_704),
        .a(_T_702),
        .b(1'h0)
    );
    wire zQuadPiece_2_A6_sqrt;
    BITWISEAND #(.width(1)) bitwiseand_5464 (
        .y(zQuadPiece_2_A6_sqrt),
        .a(_T_701),
        .b(_T_704)
    );
    wire _T_705;
    BITS #(.width(14), .high(0), .low(0)) bits_5465 (
        .y(_T_705),
        .in(_exp_PA__q)
    );
    wire _T_706;
    BITWISEAND #(.width(1)) bitwiseand_5466 (
        .y(_T_706),
        .a(cyc_A6_sqrt),
        .b(_T_705)
    );
    wire _T_707;
    BITS #(.width(53), .high(51), .low(51)) bits_5467 (
        .y(_T_707),
        .in(sigB_PA)
    );
    wire zQuadPiece_3_A6_sqrt;
    BITWISEAND #(.width(1)) bitwiseand_5468 (
        .y(zQuadPiece_3_A6_sqrt),
        .a(_T_706),
        .b(_T_707)
    );
    wire [12:0] _T_709;
    assign _T_709 = 13'h1A;
    wire [12:0] _T_711;
    wire [12:0] _WTEMP_760;
    PAD_UNSIGNED #(.width(1), .n(13)) u_pad_5469 (
        .y(_WTEMP_760),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(13)) u_mux_5470 (
        .y(_T_711),
        .sel(zQuadPiece_0_A6_sqrt),
        .a(_T_709),
        .b(_WTEMP_760)
    );
    wire [12:0] _T_713;
    assign _T_713 = 13'hBCA;
    wire [12:0] _T_715;
    wire [12:0] _WTEMP_761;
    PAD_UNSIGNED #(.width(1), .n(13)) u_pad_5471 (
        .y(_WTEMP_761),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(13)) u_mux_5472 (
        .y(_T_715),
        .sel(zQuadPiece_1_A6_sqrt),
        .a(_T_713),
        .b(_WTEMP_761)
    );
    wire [12:0] _T_716;
    BITWISEOR #(.width(13)) bitwiseor_5473 (
        .y(_T_716),
        .a(_T_711),
        .b(_T_715)
    );
    wire [12:0] _T_718;
    assign _T_718 = 13'h12D3;
    wire [12:0] _T_720;
    wire [12:0] _WTEMP_762;
    PAD_UNSIGNED #(.width(1), .n(13)) u_pad_5474 (
        .y(_WTEMP_762),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(13)) u_mux_5475 (
        .y(_T_720),
        .sel(zQuadPiece_2_A6_sqrt),
        .a(_T_718),
        .b(_WTEMP_762)
    );
    wire [12:0] _T_721;
    BITWISEOR #(.width(13)) bitwiseor_5476 (
        .y(_T_721),
        .a(_T_716),
        .b(_T_720)
    );
    wire [12:0] _T_723;
    assign _T_723 = 13'h1B17;
    wire [12:0] _T_725;
    wire [12:0] _WTEMP_763;
    PAD_UNSIGNED #(.width(1), .n(13)) u_pad_5477 (
        .y(_WTEMP_763),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(13)) u_mux_5478 (
        .y(_T_725),
        .sel(zQuadPiece_3_A6_sqrt),
        .a(_T_723),
        .b(_WTEMP_763)
    );
    wire [12:0] zComplFractK0_A6_sqrt;
    BITWISEOR #(.width(13)) bitwiseor_5479 (
        .y(zComplFractK0_A6_sqrt),
        .a(_T_721),
        .b(_T_725)
    );
    wire [8:0] _T_726;
    BITS #(.width(52), .high(48), .low(40)) bits_5480 (
        .y(_T_726),
        .in(zFractB_A4_div)
    );
    wire [8:0] _T_727;
    BITWISEOR #(.width(9)) bitwiseor_5481 (
        .y(_T_727),
        .a(_T_726),
        .b(zK2_A7_sqrt)
    );
    wire _T_729;
    EQ_UNSIGNED #(.width(1)) u_eq_5482 (
        .y(_T_729),
        .a(cyc_S),
        .b(1'h0)
    );
    wire [8:0] _T_731;
    wire [8:0] _WTEMP_764;
    PAD_UNSIGNED #(.width(1), .n(9)) u_pad_5483 (
        .y(_WTEMP_764),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(9)) u_mux_5484 (
        .y(_T_731),
        .sel(_T_729),
        .a(_nextMulAdd9A_A__q),
        .b(_WTEMP_764)
    );
    wire [8:0] mulAdd9A_A;
    BITWISEOR #(.width(9)) bitwiseor_5485 (
        .y(mulAdd9A_A),
        .a(_T_727),
        .b(_T_731)
    );
    wire [8:0] _T_732;
    BITS #(.width(52), .high(50), .low(42)) bits_5486 (
        .y(_T_732),
        .in(zFractB_A7_sqrt)
    );
    wire [8:0] _T_733;
    BITWISEOR #(.width(9)) bitwiseor_5487 (
        .y(_T_733),
        .a(zK1_A4_div),
        .b(_T_732)
    );
    wire _T_735;
    EQ_UNSIGNED #(.width(1)) u_eq_5488 (
        .y(_T_735),
        .a(cyc_S),
        .b(1'h0)
    );
    wire [8:0] _T_737;
    wire [8:0] _WTEMP_765;
    PAD_UNSIGNED #(.width(1), .n(9)) u_pad_5489 (
        .y(_WTEMP_765),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(9)) u_mux_5490 (
        .y(_T_737),
        .sel(_T_735),
        .a(_nextMulAdd9B_A__q),
        .b(_WTEMP_765)
    );
    wire [8:0] mulAdd9B_A;
    BITWISEOR #(.width(9)) bitwiseor_5491 (
        .y(mulAdd9B_A),
        .a(_T_733),
        .b(_T_737)
    );
    wire _T_738;
    BITS #(.width(1), .high(0), .low(0)) bits_5492 (
        .y(_T_738),
        .in(cyc_A7_sqrt)
    );
    wire [9:0] _T_741;
    MUX_UNSIGNED #(.width(10)) u_mux_5493 (
        .y(_T_741),
        .sel(_T_738),
        .a(10'h3FF),
        .b(10'h0)
    );
    wire [19:0] _T_742;
    CAT #(.width_a(10), .width_b(10)) cat_5494 (
        .y(_T_742),
        .a(zComplK1_A7_sqrt),
        .b(_T_741)
    );
    wire _T_743;
    BITS #(.width(1), .high(0), .low(0)) bits_5495 (
        .y(_T_743),
        .in(cyc_A6_sqrt)
    );
    wire [5:0] _T_746;
    MUX_UNSIGNED #(.width(6)) u_mux_5496 (
        .y(_T_746),
        .sel(_T_743),
        .a(6'h3F),
        .b(6'h0)
    );
    wire [13:0] _T_747;
    CAT #(.width_a(1), .width_b(13)) cat_5497 (
        .y(_T_747),
        .a(cyc_A6_sqrt),
        .b(zComplFractK0_A6_sqrt)
    );
    wire [19:0] _T_748;
    CAT #(.width_a(14), .width_b(6)) cat_5498 (
        .y(_T_748),
        .a(_T_747),
        .b(_T_746)
    );
    wire [19:0] _T_749;
    BITWISEOR #(.width(20)) bitwiseor_5499 (
        .y(_T_749),
        .a(_T_742),
        .b(_T_748)
    );
    wire _T_750;
    BITS #(.width(1), .high(0), .low(0)) bits_5500 (
        .y(_T_750),
        .in(cyc_A4_div)
    );
    wire [7:0] _T_753;
    MUX_UNSIGNED #(.width(8)) u_mux_5501 (
        .y(_T_753),
        .sel(_T_750),
        .a(8'hFF),
        .b(8'h0)
    );
    wire [12:0] _T_754;
    CAT #(.width_a(1), .width_b(12)) cat_5502 (
        .y(_T_754),
        .a(cyc_A4_div),
        .b(zComplFractK0_A4_div)
    );
    wire [20:0] _T_755;
    CAT #(.width_a(13), .width_b(8)) cat_5503 (
        .y(_T_755),
        .a(_T_754),
        .b(_T_753)
    );
    wire [20:0] _T_756;
    wire [20:0] _WTEMP_766;
    PAD_UNSIGNED #(.width(20), .n(21)) u_pad_5504 (
        .y(_WTEMP_766),
        .in(_T_749)
    );
    BITWISEOR #(.width(21)) bitwiseor_5505 (
        .y(_T_756),
        .a(_WTEMP_766),
        .b(_T_755)
    );
    wire [18:0] _T_758;
    SHL_UNSIGNED #(.width(9), .n(10)) u_shl_5506 (
        .y(_T_758),
        .in(_fractR0_A__q)
    );
    wire [20:0] _T_759;
    wire [19:0] _WTEMP_767;
    PAD_UNSIGNED #(.width(19), .n(20)) u_pad_5507 (
        .y(_WTEMP_767),
        .in(_T_758)
    );
    ADD_UNSIGNED #(.width(20)) u_add_5508 (
        .y(_T_759),
        .a(20'h40000),
        .b(_WTEMP_767)
    );
    wire [19:0] _T_760;
    TAIL #(.width(21), .n(1)) tail_5509 (
        .y(_T_760),
        .in(_T_759)
    );
    wire [19:0] _T_762;
    wire [19:0] _WTEMP_768;
    PAD_UNSIGNED #(.width(1), .n(20)) u_pad_5510 (
        .y(_WTEMP_768),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(20)) u_mux_5511 (
        .y(_T_762),
        .sel(cyc_A5_sqrt),
        .a(_T_760),
        .b(_WTEMP_768)
    );
    wire [20:0] _T_763;
    wire [20:0] _WTEMP_769;
    PAD_UNSIGNED #(.width(20), .n(21)) u_pad_5512 (
        .y(_WTEMP_769),
        .in(_T_762)
    );
    BITWISEOR #(.width(21)) bitwiseor_5513 (
        .y(_T_763),
        .a(_T_756),
        .b(_WTEMP_769)
    );
    wire _T_764;
    BITS #(.width(10), .high(9), .low(9)) bits_5514 (
        .y(_T_764),
        .in(_hiSqrR0_A_sqrt__q)
    );
    wire _T_766;
    EQ_UNSIGNED #(.width(1)) u_eq_5515 (
        .y(_T_766),
        .a(_T_764),
        .b(1'h0)
    );
    wire _T_767;
    BITWISEAND #(.width(1)) bitwiseand_5516 (
        .y(_T_767),
        .a(cyc_A4_sqrt),
        .b(_T_766)
    );
    wire [10:0] _T_770;
    wire [10:0] _WTEMP_770;
    PAD_UNSIGNED #(.width(1), .n(11)) u_pad_5517 (
        .y(_WTEMP_770),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(11)) u_mux_5518 (
        .y(_T_770),
        .sel(_T_767),
        .a(11'h400),
        .b(_WTEMP_770)
    );
    wire [20:0] _T_771;
    wire [20:0] _WTEMP_771;
    PAD_UNSIGNED #(.width(11), .n(21)) u_pad_5519 (
        .y(_WTEMP_771),
        .in(_T_770)
    );
    BITWISEOR #(.width(21)) bitwiseor_5520 (
        .y(_T_771),
        .a(_T_763),
        .b(_WTEMP_771)
    );
    wire _T_772;
    BITS #(.width(10), .high(9), .low(9)) bits_5521 (
        .y(_T_772),
        .in(_hiSqrR0_A_sqrt__q)
    );
    wire _T_773;
    BITWISEAND #(.width(1)) bitwiseand_5522 (
        .y(_T_773),
        .a(cyc_A4_sqrt),
        .b(_T_772)
    );
    wire _T_774;
    BITWISEOR #(.width(1)) bitwiseor_5523 (
        .y(_T_774),
        .a(_T_773),
        .b(cyc_A3_div)
    );
    wire [20:0] _T_775;
    BITS #(.width(53), .high(46), .low(26)) bits_5524 (
        .y(_T_775),
        .in(sigB_PA)
    );
    wire [21:0] _T_777;
    wire [20:0] _WTEMP_772;
    PAD_UNSIGNED #(.width(11), .n(21)) u_pad_5525 (
        .y(_WTEMP_772),
        .in(11'h400)
    );
    ADD_UNSIGNED #(.width(21)) u_add_5526 (
        .y(_T_777),
        .a(_T_775),
        .b(_WTEMP_772)
    );
    wire [20:0] _T_778;
    TAIL #(.width(22), .n(1)) tail_5527 (
        .y(_T_778),
        .in(_T_777)
    );
    wire [20:0] _T_780;
    wire [20:0] _WTEMP_773;
    PAD_UNSIGNED #(.width(1), .n(21)) u_pad_5528 (
        .y(_WTEMP_773),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(21)) u_mux_5529 (
        .y(_T_780),
        .sel(_T_774),
        .a(_T_778),
        .b(_WTEMP_773)
    );
    wire [20:0] _T_781;
    BITWISEOR #(.width(21)) bitwiseor_5530 (
        .y(_T_781),
        .a(_T_771),
        .b(_T_780)
    );
    wire _T_782;
    BITWISEOR #(.width(1)) bitwiseor_5531 (
        .y(_T_782),
        .a(cyc_A3_sqrt),
        .b(cyc_A2)
    );
    wire [20:0] _T_784;
    wire [20:0] _WTEMP_774;
    PAD_UNSIGNED #(.width(1), .n(21)) u_pad_5532 (
        .y(_WTEMP_774),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(21)) u_mux_5533 (
        .y(_T_784),
        .sel(_T_782),
        .a(_partNegSigma0_A__q),
        .b(_WTEMP_774)
    );
    wire [20:0] _T_785;
    BITWISEOR #(.width(21)) bitwiseor_5534 (
        .y(_T_785),
        .a(_T_781),
        .b(_T_784)
    );
    wire [24:0] _T_786;
    SHL_UNSIGNED #(.width(9), .n(16)) u_shl_5535 (
        .y(_T_786),
        .in(_fractR0_A__q)
    );
    wire [24:0] _T_788;
    wire [24:0] _WTEMP_775;
    PAD_UNSIGNED #(.width(1), .n(25)) u_pad_5536 (
        .y(_WTEMP_775),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(25)) u_mux_5537 (
        .y(_T_788),
        .sel(cyc_A1_sqrt),
        .a(_T_786),
        .b(_WTEMP_775)
    );
    wire [24:0] _T_789;
    wire [24:0] _WTEMP_776;
    PAD_UNSIGNED #(.width(21), .n(25)) u_pad_5538 (
        .y(_WTEMP_776),
        .in(_T_785)
    );
    BITWISEOR #(.width(25)) bitwiseor_5539 (
        .y(_T_789),
        .a(_WTEMP_776),
        .b(_T_788)
    );
    wire [23:0] _T_790;
    SHL_UNSIGNED #(.width(9), .n(15)) u_shl_5540 (
        .y(_T_790),
        .in(_fractR0_A__q)
    );
    wire [23:0] _T_792;
    wire [23:0] _WTEMP_777;
    PAD_UNSIGNED #(.width(1), .n(24)) u_pad_5541 (
        .y(_WTEMP_777),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(24)) u_mux_5542 (
        .y(_T_792),
        .sel(cyc_A1_div),
        .a(_T_790),
        .b(_WTEMP_777)
    );
    wire [24:0] mulAdd9C_A;
    wire [24:0] _WTEMP_778;
    PAD_UNSIGNED #(.width(24), .n(25)) u_pad_5543 (
        .y(_WTEMP_778),
        .in(_T_792)
    );
    BITWISEOR #(.width(25)) bitwiseor_5544 (
        .y(mulAdd9C_A),
        .a(_T_789),
        .b(_WTEMP_778)
    );
    wire [17:0] _T_793;
    MUL2_UNSIGNED #(.width_a(9), .width_b(9)) u_mul2_5545 (
        .y(_T_793),
        .a(mulAdd9A_A),
        .b(mulAdd9B_A)
    );
    wire [17:0] _T_795;
    BITS #(.width(25), .high(17), .low(0)) bits_5546 (
        .y(_T_795),
        .in(mulAdd9C_A)
    );
    wire [18:0] _T_796;
    CAT #(.width_a(1), .width_b(18)) cat_5547 (
        .y(_T_796),
        .a(1'h0),
        .b(_T_795)
    );
    wire [19:0] _T_797;
    wire [18:0] _WTEMP_779;
    PAD_UNSIGNED #(.width(18), .n(19)) u_pad_5548 (
        .y(_WTEMP_779),
        .in(_T_793)
    );
    ADD_UNSIGNED #(.width(19)) u_add_5549 (
        .y(_T_797),
        .a(_WTEMP_779),
        .b(_T_796)
    );
    wire [18:0] loMulAdd9Out_A;
    TAIL #(.width(20), .n(1)) tail_5550 (
        .y(loMulAdd9Out_A),
        .in(_T_797)
    );
    wire _T_798;
    BITS #(.width(19), .high(18), .low(18)) bits_5551 (
        .y(_T_798),
        .in(loMulAdd9Out_A)
    );
    wire [6:0] _T_799;
    BITS #(.width(25), .high(24), .low(18)) bits_5552 (
        .y(_T_799),
        .in(mulAdd9C_A)
    );
    wire [7:0] _T_801;
    wire [6:0] _WTEMP_780;
    PAD_UNSIGNED #(.width(1), .n(7)) u_pad_5553 (
        .y(_WTEMP_780),
        .in(1'h1)
    );
    ADD_UNSIGNED #(.width(7)) u_add_5554 (
        .y(_T_801),
        .a(_T_799),
        .b(_WTEMP_780)
    );
    wire [6:0] _T_802;
    TAIL #(.width(8), .n(1)) tail_5555 (
        .y(_T_802),
        .in(_T_801)
    );
    wire [6:0] _T_803;
    BITS #(.width(25), .high(24), .low(18)) bits_5556 (
        .y(_T_803),
        .in(mulAdd9C_A)
    );
    wire [6:0] _T_804;
    MUX_UNSIGNED #(.width(7)) u_mux_5557 (
        .y(_T_804),
        .sel(_T_798),
        .a(_T_802),
        .b(_T_803)
    );
    wire [17:0] _T_805;
    BITS #(.width(19), .high(17), .low(0)) bits_5558 (
        .y(_T_805),
        .in(loMulAdd9Out_A)
    );
    wire [24:0] mulAdd9Out_A;
    CAT #(.width_a(7), .width_b(18)) cat_5559 (
        .y(mulAdd9Out_A),
        .a(_T_804),
        .b(_T_805)
    );
    wire _T_806;
    BITS #(.width(25), .high(19), .low(19)) bits_5560 (
        .y(_T_806),
        .in(mulAdd9Out_A)
    );
    wire _T_807;
    BITWISEAND #(.width(1)) bitwiseand_5561 (
        .y(_T_807),
        .a(cyc_A6_sqrt),
        .b(_T_806)
    );
    wire [24:0] _T_808;
    BITWISENOT #(.width(25)) bitwisenot_5562 (
        .y(_T_808),
        .in(mulAdd9Out_A)
    );
    wire [14:0] _T_809;
    SHR_UNSIGNED #(.width(25), .n(10)) u_shr_5563 (
        .y(_T_809),
        .in(_T_808)
    );
    wire [14:0] _T_811;
    wire [14:0] _WTEMP_781;
    PAD_UNSIGNED #(.width(1), .n(15)) u_pad_5564 (
        .y(_WTEMP_781),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(15)) u_mux_5565 (
        .y(_T_811),
        .sel(_T_807),
        .a(_T_809),
        .b(_WTEMP_781)
    );
    wire [8:0] zFractR0_A6_sqrt;
    BITS #(.width(15), .high(8), .low(0)) bits_5566 (
        .y(zFractR0_A6_sqrt),
        .in(_T_811)
    );
    wire _T_812;
    BITS #(.width(14), .high(0), .low(0)) bits_5567 (
        .y(_T_812),
        .in(_exp_PA__q)
    );
    wire [25:0] _T_813;
    SHL_UNSIGNED #(.width(25), .n(1)) u_shl_5568 (
        .y(_T_813),
        .in(mulAdd9Out_A)
    );
    wire [25:0] sqrR0_A5_sqrt;
    wire [25:0] _WTEMP_782;
    PAD_UNSIGNED #(.width(25), .n(26)) u_pad_5569 (
        .y(_WTEMP_782),
        .in(mulAdd9Out_A)
    );
    MUX_UNSIGNED #(.width(26)) u_mux_5570 (
        .y(sqrR0_A5_sqrt),
        .sel(_T_812),
        .a(_T_813),
        .b(_WTEMP_782)
    );
    wire _T_814;
    BITS #(.width(25), .high(20), .low(20)) bits_5571 (
        .y(_T_814),
        .in(mulAdd9Out_A)
    );
    wire _T_815;
    BITWISEAND #(.width(1)) bitwiseand_5572 (
        .y(_T_815),
        .a(cyc_A4_div),
        .b(_T_814)
    );
    wire [24:0] _T_816;
    BITWISENOT #(.width(25)) bitwisenot_5573 (
        .y(_T_816),
        .in(mulAdd9Out_A)
    );
    wire [13:0] _T_817;
    SHR_UNSIGNED #(.width(25), .n(11)) u_shr_5574 (
        .y(_T_817),
        .in(_T_816)
    );
    wire [13:0] _T_819;
    wire [13:0] _WTEMP_783;
    PAD_UNSIGNED #(.width(1), .n(14)) u_pad_5575 (
        .y(_WTEMP_783),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(14)) u_mux_5576 (
        .y(_T_819),
        .sel(_T_815),
        .a(_T_817),
        .b(_WTEMP_783)
    );
    wire [8:0] zFractR0_A4_div;
    BITS #(.width(14), .high(8), .low(0)) bits_5577 (
        .y(zFractR0_A4_div),
        .in(_T_819)
    );
    wire _T_820;
    BITS #(.width(25), .high(11), .low(11)) bits_5578 (
        .y(_T_820),
        .in(mulAdd9Out_A)
    );
    wire _T_821;
    BITWISEAND #(.width(1)) bitwiseand_5579 (
        .y(_T_821),
        .a(cyc_A2),
        .b(_T_820)
    );
    wire [24:0] _T_822;
    BITWISENOT #(.width(25)) bitwisenot_5580 (
        .y(_T_822),
        .in(mulAdd9Out_A)
    );
    wire [22:0] _T_823;
    SHR_UNSIGNED #(.width(25), .n(2)) u_shr_5581 (
        .y(_T_823),
        .in(_T_822)
    );
    wire [22:0] _T_825;
    wire [22:0] _WTEMP_784;
    PAD_UNSIGNED #(.width(1), .n(23)) u_pad_5582 (
        .y(_WTEMP_784),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(23)) u_mux_5583 (
        .y(_T_825),
        .sel(_T_821),
        .a(_T_823),
        .b(_WTEMP_784)
    );
    wire [8:0] zSigma0_A2;
    BITS #(.width(23), .high(8), .low(0)) bits_5584 (
        .y(zSigma0_A2),
        .in(_T_825)
    );
    wire [14:0] _T_826;
    SHR_UNSIGNED #(.width(25), .n(10)) u_shr_5585 (
        .y(_T_826),
        .in(mulAdd9Out_A)
    );
    wire [15:0] _T_827;
    SHR_UNSIGNED #(.width(25), .n(9)) u_shr_5586 (
        .y(_T_827),
        .in(mulAdd9Out_A)
    );
    wire [15:0] _T_828;
    wire [15:0] _WTEMP_785;
    PAD_UNSIGNED #(.width(15), .n(16)) u_pad_5587 (
        .y(_WTEMP_785),
        .in(_T_826)
    );
    MUX_UNSIGNED #(.width(16)) u_mux_5588 (
        .y(_T_828),
        .sel(_sqrtOp_PA__q),
        .a(_WTEMP_785),
        .b(_T_827)
    );
    wire [14:0] fractR1_A1;
    BITS #(.width(16), .high(14), .low(0)) bits_5589 (
        .y(fractR1_A1),
        .in(_T_828)
    );
    wire [15:0] r1_A1;
    CAT #(.width_a(1), .width_b(15)) cat_5590 (
        .y(r1_A1),
        .a(1'h1),
        .b(fractR1_A1)
    );
    wire _T_830;
    BITS #(.width(14), .high(0), .low(0)) bits_5591 (
        .y(_T_830),
        .in(_exp_PA__q)
    );
    wire [16:0] _T_831;
    SHL_UNSIGNED #(.width(16), .n(1)) u_shl_5592 (
        .y(_T_831),
        .in(r1_A1)
    );
    wire [16:0] ER1_A1_sqrt;
    wire [16:0] _WTEMP_786;
    PAD_UNSIGNED #(.width(16), .n(17)) u_pad_5593 (
        .y(_WTEMP_786),
        .in(r1_A1)
    );
    MUX_UNSIGNED #(.width(17)) u_mux_5594 (
        .y(ER1_A1_sqrt),
        .sel(_T_830),
        .a(_T_831),
        .b(_WTEMP_786)
    );
    wire _T_832;
    BITWISEOR #(.width(1)) bitwiseor_5595 (
        .y(_T_832),
        .a(cyc_A6_sqrt),
        .b(cyc_A4_div)
    );
    wire [8:0] _T_833;
    BITWISEOR #(.width(9)) bitwiseor_5596 (
        .y(_T_833),
        .a(zFractR0_A6_sqrt),
        .b(zFractR0_A4_div)
    );
    wire [15:0] _T_834;
    SHR_UNSIGNED #(.width(26), .n(10)) u_shr_5597 (
        .y(_T_834),
        .in(sqrR0_A5_sqrt)
    );
    wire _T_835;
    BITWISEOR #(.width(1)) bitwiseor_5598 (
        .y(_T_835),
        .a(cyc_A4_sqrt),
        .b(cyc_A3)
    );
    wire [15:0] _T_836;
    SHR_UNSIGNED #(.width(25), .n(9)) u_shr_5599 (
        .y(_T_836),
        .in(mulAdd9Out_A)
    );
    wire [24:0] _T_837;
    wire [24:0] _WTEMP_787;
    PAD_UNSIGNED #(.width(16), .n(25)) u_pad_5600 (
        .y(_WTEMP_787),
        .in(_T_836)
    );
    MUX_UNSIGNED #(.width(25)) u_mux_5601 (
        .y(_T_837),
        .sel(cyc_A4_sqrt),
        .a(mulAdd9Out_A),
        .b(_WTEMP_787)
    );
    wire [20:0] _T_838;
    BITS #(.width(25), .high(20), .low(0)) bits_5602 (
        .y(_T_838),
        .in(_T_837)
    );
    wire _T_839;
    BITWISEOR #(.width(1)) bitwiseor_5603 (
        .y(_T_839),
        .a(cyc_A7_sqrt),
        .b(cyc_A6_sqrt)
    );
    wire _T_840;
    BITWISEOR #(.width(1)) bitwiseor_5604 (
        .y(_T_840),
        .a(_T_839),
        .b(cyc_A5_sqrt)
    );
    wire _T_841;
    BITWISEOR #(.width(1)) bitwiseor_5605 (
        .y(_T_841),
        .a(_T_840),
        .b(cyc_A4)
    );
    wire _T_842;
    BITWISEOR #(.width(1)) bitwiseor_5606 (
        .y(_T_842),
        .a(_T_841),
        .b(cyc_A3)
    );
    wire _T_843;
    BITWISEOR #(.width(1)) bitwiseor_5607 (
        .y(_T_843),
        .a(_T_842),
        .b(cyc_A2)
    );
    wire [24:0] _T_844;
    BITWISENOT #(.width(25)) bitwisenot_5608 (
        .y(_T_844),
        .in(mulAdd9Out_A)
    );
    wire [13:0] _T_845;
    SHR_UNSIGNED #(.width(25), .n(11)) u_shr_5609 (
        .y(_T_845),
        .in(_T_844)
    );
    wire [13:0] _T_847;
    wire [13:0] _WTEMP_788;
    PAD_UNSIGNED #(.width(1), .n(14)) u_pad_5610 (
        .y(_WTEMP_788),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(14)) u_mux_5611 (
        .y(_T_847),
        .sel(cyc_A7_sqrt),
        .a(_T_845),
        .b(_WTEMP_788)
    );
    wire [13:0] _T_848;
    wire [13:0] _WTEMP_789;
    PAD_UNSIGNED #(.width(9), .n(14)) u_pad_5612 (
        .y(_WTEMP_789),
        .in(zFractR0_A6_sqrt)
    );
    BITWISEOR #(.width(14)) bitwiseor_5613 (
        .y(_T_848),
        .a(_T_847),
        .b(_WTEMP_789)
    );
    wire [8:0] _T_849;
    BITS #(.width(53), .high(43), .low(35)) bits_5614 (
        .y(_T_849),
        .in(sigB_PA)
    );
    wire [8:0] _T_851;
    wire [8:0] _WTEMP_790;
    PAD_UNSIGNED #(.width(1), .n(9)) u_pad_5615 (
        .y(_WTEMP_790),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(9)) u_mux_5616 (
        .y(_T_851),
        .sel(cyc_A4_sqrt),
        .a(_T_849),
        .b(_WTEMP_790)
    );
    wire [13:0] _T_852;
    wire [13:0] _WTEMP_791;
    PAD_UNSIGNED #(.width(9), .n(14)) u_pad_5617 (
        .y(_WTEMP_791),
        .in(_T_851)
    );
    BITWISEOR #(.width(14)) bitwiseor_5618 (
        .y(_T_852),
        .a(_T_848),
        .b(_WTEMP_791)
    );
    wire [8:0] _T_853;
    BITS #(.width(52), .high(43), .low(35)) bits_5619 (
        .y(_T_853),
        .in(zFractB_A4_div)
    );
    wire [13:0] _T_854;
    wire [13:0] _WTEMP_792;
    PAD_UNSIGNED #(.width(9), .n(14)) u_pad_5620 (
        .y(_WTEMP_792),
        .in(_T_853)
    );
    BITWISEOR #(.width(14)) bitwiseor_5621 (
        .y(_T_854),
        .a(_T_852),
        .b(_WTEMP_792)
    );
    wire _T_855;
    BITWISEOR #(.width(1)) bitwiseor_5622 (
        .y(_T_855),
        .a(cyc_A5_sqrt),
        .b(cyc_A3)
    );
    wire [8:0] _T_856;
    BITS #(.width(53), .high(52), .low(44)) bits_5623 (
        .y(_T_856),
        .in(sigB_PA)
    );
    wire [8:0] _T_858;
    wire [8:0] _WTEMP_793;
    PAD_UNSIGNED #(.width(1), .n(9)) u_pad_5624 (
        .y(_WTEMP_793),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(9)) u_mux_5625 (
        .y(_T_858),
        .sel(_T_855),
        .a(_T_856),
        .b(_WTEMP_793)
    );
    wire [13:0] _T_859;
    wire [13:0] _WTEMP_794;
    PAD_UNSIGNED #(.width(9), .n(14)) u_pad_5626 (
        .y(_WTEMP_794),
        .in(_T_858)
    );
    BITWISEOR #(.width(14)) bitwiseor_5627 (
        .y(_T_859),
        .a(_T_854),
        .b(_WTEMP_794)
    );
    wire [13:0] _T_860;
    wire [13:0] _WTEMP_795;
    PAD_UNSIGNED #(.width(9), .n(14)) u_pad_5628 (
        .y(_WTEMP_795),
        .in(zSigma0_A2)
    );
    BITWISEOR #(.width(14)) bitwiseor_5629 (
        .y(_T_860),
        .a(_T_859),
        .b(_WTEMP_795)
    );
    wire _T_861;
    BITWISEOR #(.width(1)) bitwiseor_5630 (
        .y(_T_861),
        .a(cyc_A7_sqrt),
        .b(cyc_A6_sqrt)
    );
    wire _T_862;
    BITWISEOR #(.width(1)) bitwiseor_5631 (
        .y(_T_862),
        .a(_T_861),
        .b(cyc_A5_sqrt)
    );
    wire _T_863;
    BITWISEOR #(.width(1)) bitwiseor_5632 (
        .y(_T_863),
        .a(_T_862),
        .b(cyc_A4)
    );
    wire _T_864;
    BITWISEOR #(.width(1)) bitwiseor_5633 (
        .y(_T_864),
        .a(_T_863),
        .b(cyc_A2)
    );
    wire [8:0] _T_865;
    BITS #(.width(52), .high(50), .low(42)) bits_5634 (
        .y(_T_865),
        .in(zFractB_A7_sqrt)
    );
    wire [8:0] _T_866;
    BITWISEOR #(.width(9)) bitwiseor_5635 (
        .y(_T_866),
        .a(_T_865),
        .b(zFractR0_A6_sqrt)
    );
    wire [8:0] _T_867;
    BITS #(.width(26), .high(9), .low(1)) bits_5636 (
        .y(_T_867),
        .in(sqrR0_A5_sqrt)
    );
    wire [8:0] _T_869;
    wire [8:0] _WTEMP_796;
    PAD_UNSIGNED #(.width(1), .n(9)) u_pad_5637 (
        .y(_WTEMP_796),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(9)) u_mux_5638 (
        .y(_T_869),
        .sel(cyc_A5_sqrt),
        .a(_T_867),
        .b(_WTEMP_796)
    );
    wire [8:0] _T_870;
    BITWISEOR #(.width(9)) bitwiseor_5639 (
        .y(_T_870),
        .a(_T_866),
        .b(_T_869)
    );
    wire [8:0] _T_871;
    BITWISEOR #(.width(9)) bitwiseor_5640 (
        .y(_T_871),
        .a(_T_870),
        .b(zFractR0_A4_div)
    );
    wire [8:0] _T_872;
    BITS #(.width(10), .high(8), .low(0)) bits_5641 (
        .y(_T_872),
        .in(_hiSqrR0_A_sqrt__q)
    );
    wire [8:0] _T_874;
    wire [8:0] _WTEMP_797;
    PAD_UNSIGNED #(.width(1), .n(9)) u_pad_5642 (
        .y(_WTEMP_797),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(9)) u_mux_5643 (
        .y(_T_874),
        .sel(cyc_A4_sqrt),
        .a(_T_872),
        .b(_WTEMP_797)
    );
    wire [8:0] _T_875;
    BITWISEOR #(.width(9)) bitwiseor_5644 (
        .y(_T_875),
        .a(_T_871),
        .b(_T_874)
    );
    wire [7:0] _T_877;
    BITS #(.width(9), .high(8), .low(1)) bits_5645 (
        .y(_T_877),
        .in(_fractR0_A__q)
    );
    wire [8:0] _T_878;
    CAT #(.width_a(1), .width_b(8)) cat_5646 (
        .y(_T_878),
        .a(1'h1),
        .b(_T_877)
    );
    wire [8:0] _T_880;
    wire [8:0] _WTEMP_798;
    PAD_UNSIGNED #(.width(1), .n(9)) u_pad_5647 (
        .y(_WTEMP_798),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(9)) u_mux_5648 (
        .y(_T_880),
        .sel(cyc_A2),
        .a(_T_878),
        .b(_WTEMP_798)
    );
    wire [8:0] _T_881;
    BITWISEOR #(.width(9)) bitwiseor_5649 (
        .y(_T_881),
        .a(_T_875),
        .b(_T_880)
    );
    wire _T_882;
    BITWISEOR #(.width(1)) bitwiseor_5650 (
        .y(_T_882),
        .a(cyc_A1),
        .b(cyc_B7_sqrt)
    );
    wire _T_883;
    BITWISEOR #(.width(1)) bitwiseor_5651 (
        .y(_T_883),
        .a(_T_882),
        .b(cyc_B6_div)
    );
    wire _T_884;
    BITWISEOR #(.width(1)) bitwiseor_5652 (
        .y(_T_884),
        .a(_T_883),
        .b(cyc_B4)
    );
    wire _T_885;
    BITWISEOR #(.width(1)) bitwiseor_5653 (
        .y(_T_885),
        .a(_T_884),
        .b(cyc_B3)
    );
    wire _T_886;
    BITWISEOR #(.width(1)) bitwiseor_5654 (
        .y(_T_886),
        .a(_T_885),
        .b(cyc_C6_sqrt)
    );
    wire _T_887;
    BITWISEOR #(.width(1)) bitwiseor_5655 (
        .y(_T_887),
        .a(_T_886),
        .b(cyc_C4)
    );
    wire _T_888;
    BITWISEOR #(.width(1)) bitwiseor_5656 (
        .y(_T_888),
        .a(_T_887),
        .b(cyc_C1)
    );
    wire [52:0] _T_889;
    SHL_UNSIGNED #(.width(17), .n(36)) u_shl_5657 (
        .y(_T_889),
        .in(ER1_A1_sqrt)
    );
    wire [52:0] _T_891;
    wire [52:0] _WTEMP_799;
    PAD_UNSIGNED #(.width(1), .n(53)) u_pad_5658 (
        .y(_WTEMP_799),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(53)) u_mux_5659 (
        .y(_T_891),
        .sel(cyc_A1_sqrt),
        .a(_T_889),
        .b(_WTEMP_799)
    );
    wire _T_892;
    BITWISEOR #(.width(1)) bitwiseor_5660 (
        .y(_T_892),
        .a(cyc_B7_sqrt),
        .b(cyc_A1_div)
    );
    wire [52:0] _T_894;
    wire [52:0] _WTEMP_800;
    PAD_UNSIGNED #(.width(1), .n(53)) u_pad_5661 (
        .y(_WTEMP_800),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(53)) u_mux_5662 (
        .y(_T_894),
        .sel(_T_892),
        .a(sigB_PA),
        .b(_WTEMP_800)
    );
    wire [52:0] _T_895;
    BITWISEOR #(.width(53)) bitwiseor_5663 (
        .y(_T_895),
        .a(_T_891),
        .b(_T_894)
    );
    wire [52:0] _T_897;
    wire [52:0] _WTEMP_801;
    PAD_UNSIGNED #(.width(1), .n(53)) u_pad_5664 (
        .y(_WTEMP_801),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(53)) u_mux_5665 (
        .y(_T_897),
        .sel(cyc_B6_div),
        .a(sigA_PA),
        .b(_WTEMP_801)
    );
    wire [52:0] _T_898;
    BITWISEOR #(.width(53)) bitwiseor_5666 (
        .y(_T_898),
        .a(_T_895),
        .b(_T_897)
    );
    wire [33:0] _T_899;
    BITS #(.width(46), .high(45), .low(12)) bits_5667 (
        .y(_T_899),
        .in(zSigma1_B4)
    );
    wire [52:0] _T_900;
    wire [52:0] _WTEMP_802;
    PAD_UNSIGNED #(.width(34), .n(53)) u_pad_5668 (
        .y(_WTEMP_802),
        .in(_T_899)
    );
    BITWISEOR #(.width(53)) bitwiseor_5669 (
        .y(_T_900),
        .a(_T_898),
        .b(_WTEMP_802)
    );
    wire _T_901;
    BITWISEOR #(.width(1)) bitwiseor_5670 (
        .y(_T_901),
        .a(cyc_B3),
        .b(cyc_C6_sqrt)
    );
    wire [45:0] _T_902;
    BITS #(.width(58), .high(57), .low(12)) bits_5671 (
        .y(_T_902),
        .in(sigXNU_B3_CX)
    );
    wire [45:0] _T_904;
    wire [45:0] _WTEMP_803;
    PAD_UNSIGNED #(.width(1), .n(46)) u_pad_5672 (
        .y(_WTEMP_803),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(46)) u_mux_5673 (
        .y(_T_904),
        .sel(_T_901),
        .a(_T_902),
        .b(_WTEMP_803)
    );
    wire [52:0] _T_905;
    wire [52:0] _WTEMP_804;
    PAD_UNSIGNED #(.width(46), .n(53)) u_pad_5674 (
        .y(_WTEMP_804),
        .in(_T_904)
    );
    BITWISEOR #(.width(53)) bitwiseor_5675 (
        .y(_T_905),
        .a(_T_900),
        .b(_WTEMP_804)
    );
    wire [32:0] _T_906;
    BITS #(.width(58), .high(57), .low(25)) bits_5676 (
        .y(_T_906),
        .in(_sigXN_C__q)
    );
    wire [45:0] _T_907;
    SHL_UNSIGNED #(.width(33), .n(13)) u_shl_5677 (
        .y(_T_907),
        .in(_T_906)
    );
    wire [45:0] _T_909;
    wire [45:0] _WTEMP_805;
    PAD_UNSIGNED #(.width(1), .n(46)) u_pad_5678 (
        .y(_WTEMP_805),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(46)) u_mux_5679 (
        .y(_T_909),
        .sel(cyc_C4_div),
        .a(_T_907),
        .b(_WTEMP_805)
    );
    wire [52:0] _T_910;
    wire [52:0] _WTEMP_806;
    PAD_UNSIGNED #(.width(46), .n(53)) u_pad_5680 (
        .y(_WTEMP_806),
        .in(_T_909)
    );
    BITWISEOR #(.width(53)) bitwiseor_5681 (
        .y(_T_910),
        .a(_T_905),
        .b(_WTEMP_806)
    );
    wire [45:0] _T_911;
    SHL_UNSIGNED #(.width(31), .n(15)) u_shl_5682 (
        .y(_T_911),
        .in(_u_C_sqrt__q)
    );
    wire [45:0] _T_913;
    wire [45:0] _WTEMP_807;
    PAD_UNSIGNED #(.width(1), .n(46)) u_pad_5683 (
        .y(_WTEMP_807),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(46)) u_mux_5684 (
        .y(_T_913),
        .sel(cyc_C4_sqrt),
        .a(_T_911),
        .b(_WTEMP_807)
    );
    wire [52:0] _T_914;
    wire [52:0] _WTEMP_808;
    PAD_UNSIGNED #(.width(46), .n(53)) u_pad_5685 (
        .y(_WTEMP_808),
        .in(_T_913)
    );
    BITWISEOR #(.width(53)) bitwiseor_5686 (
        .y(_T_914),
        .a(_T_910),
        .b(_WTEMP_808)
    );
    wire [52:0] _T_916;
    wire [52:0] _WTEMP_809;
    PAD_UNSIGNED #(.width(1), .n(53)) u_pad_5687 (
        .y(_WTEMP_809),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(53)) u_mux_5688 (
        .y(_T_916),
        .sel(cyc_C1_div),
        .a(sigB_PC),
        .b(_WTEMP_809)
    );
    wire [52:0] _T_917;
    BITWISEOR #(.width(53)) bitwiseor_5689 (
        .y(_T_917),
        .a(_T_914),
        .b(_T_916)
    );
    wire [53:0] _T_918;
    wire [53:0] _WTEMP_810;
    PAD_UNSIGNED #(.width(53), .n(54)) u_pad_5690 (
        .y(_WTEMP_810),
        .in(_T_917)
    );
    BITWISEOR #(.width(54)) bitwiseor_5691 (
        .y(_T_918),
        .a(_WTEMP_810),
        .b(zComplSigT_C1_sqrt)
    );
    wire _T_919;
    BITWISEOR #(.width(1)) bitwiseor_5692 (
        .y(_T_919),
        .a(cyc_A1),
        .b(cyc_B7_sqrt)
    );
    wire _T_920;
    BITWISEOR #(.width(1)) bitwiseor_5693 (
        .y(_T_920),
        .a(_T_919),
        .b(cyc_B6_sqrt)
    );
    wire _T_921;
    BITWISEOR #(.width(1)) bitwiseor_5694 (
        .y(_T_921),
        .a(_T_920),
        .b(cyc_B4)
    );
    wire _T_922;
    BITWISEOR #(.width(1)) bitwiseor_5695 (
        .y(_T_922),
        .a(_T_921),
        .b(cyc_C6_sqrt)
    );
    wire _T_923;
    BITWISEOR #(.width(1)) bitwiseor_5696 (
        .y(_T_923),
        .a(_T_922),
        .b(cyc_C4)
    );
    wire _T_924;
    BITWISEOR #(.width(1)) bitwiseor_5697 (
        .y(_T_924),
        .a(_T_923),
        .b(cyc_C1)
    );
    wire [51:0] _T_925;
    SHL_UNSIGNED #(.width(16), .n(36)) u_shl_5698 (
        .y(_T_925),
        .in(r1_A1)
    );
    wire [51:0] _T_927;
    wire [51:0] _WTEMP_811;
    PAD_UNSIGNED #(.width(1), .n(52)) u_pad_5699 (
        .y(_WTEMP_811),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(52)) u_mux_5700 (
        .y(_T_927),
        .sel(cyc_A1),
        .a(_T_925),
        .b(_WTEMP_811)
    );
    wire [50:0] _T_928;
    SHL_UNSIGNED #(.width(32), .n(19)) u_shl_5701 (
        .y(_T_928),
        .in(_ESqrR1_B_sqrt__q)
    );
    wire [50:0] _T_930;
    wire [50:0] _WTEMP_812;
    PAD_UNSIGNED #(.width(1), .n(51)) u_pad_5702 (
        .y(_WTEMP_812),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(51)) u_mux_5703 (
        .y(_T_930),
        .sel(cyc_B7_sqrt),
        .a(_T_928),
        .b(_WTEMP_812)
    );
    wire [51:0] _T_931;
    wire [51:0] _WTEMP_813;
    PAD_UNSIGNED #(.width(51), .n(52)) u_pad_5704 (
        .y(_WTEMP_813),
        .in(_T_930)
    );
    BITWISEOR #(.width(52)) bitwiseor_5705 (
        .y(_T_931),
        .a(_T_927),
        .b(_WTEMP_813)
    );
    wire [52:0] _T_932;
    SHL_UNSIGNED #(.width(17), .n(36)) u_shl_5706 (
        .y(_T_932),
        .in(_ER1_B_sqrt__q)
    );
    wire [52:0] _T_934;
    wire [52:0] _WTEMP_814;
    PAD_UNSIGNED #(.width(1), .n(53)) u_pad_5707 (
        .y(_WTEMP_814),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(53)) u_mux_5708 (
        .y(_T_934),
        .sel(cyc_B6_sqrt),
        .a(_T_932),
        .b(_WTEMP_814)
    );
    wire [52:0] _T_935;
    wire [52:0] _WTEMP_815;
    PAD_UNSIGNED #(.width(52), .n(53)) u_pad_5709 (
        .y(_WTEMP_815),
        .in(_T_931)
    );
    BITWISEOR #(.width(53)) bitwiseor_5710 (
        .y(_T_935),
        .a(_WTEMP_815),
        .b(_T_934)
    );
    wire [52:0] _T_936;
    wire [52:0] _WTEMP_816;
    PAD_UNSIGNED #(.width(46), .n(53)) u_pad_5711 (
        .y(_WTEMP_816),
        .in(zSigma1_B4)
    );
    BITWISEOR #(.width(53)) bitwiseor_5712 (
        .y(_T_936),
        .a(_T_935),
        .b(_WTEMP_816)
    );
    wire [29:0] _T_937;
    BITS #(.width(33), .high(30), .low(1)) bits_5713 (
        .y(_T_937),
        .in(_sqrSigma1_C__q)
    );
    wire [29:0] _T_939;
    wire [29:0] _WTEMP_817;
    PAD_UNSIGNED #(.width(1), .n(30)) u_pad_5714 (
        .y(_WTEMP_817),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(30)) u_mux_5715 (
        .y(_T_939),
        .sel(cyc_C6_sqrt),
        .a(_T_937),
        .b(_WTEMP_817)
    );
    wire [52:0] _T_940;
    wire [52:0] _WTEMP_818;
    PAD_UNSIGNED #(.width(30), .n(53)) u_pad_5716 (
        .y(_WTEMP_818),
        .in(_T_939)
    );
    BITWISEOR #(.width(53)) bitwiseor_5717 (
        .y(_T_940),
        .a(_T_936),
        .b(_WTEMP_818)
    );
    wire [32:0] _T_942;
    wire [32:0] _WTEMP_819;
    PAD_UNSIGNED #(.width(1), .n(33)) u_pad_5718 (
        .y(_WTEMP_819),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(33)) u_mux_5719 (
        .y(_T_942),
        .sel(cyc_C4),
        .a(_sqrSigma1_C__q),
        .b(_WTEMP_819)
    );
    wire [52:0] _T_943;
    wire [52:0] _WTEMP_820;
    PAD_UNSIGNED #(.width(33), .n(53)) u_pad_5720 (
        .y(_WTEMP_820),
        .in(_T_942)
    );
    BITWISEOR #(.width(53)) bitwiseor_5721 (
        .y(_T_943),
        .a(_T_940),
        .b(_WTEMP_820)
    );
    wire [53:0] _T_944;
    wire [53:0] _WTEMP_821;
    PAD_UNSIGNED #(.width(53), .n(54)) u_pad_5722 (
        .y(_WTEMP_821),
        .in(_T_943)
    );
    BITWISEOR #(.width(54)) bitwiseor_5723 (
        .y(_T_944),
        .a(_WTEMP_821),
        .b(zComplSigT_C1)
    );
    wire _T_945;
    BITWISEOR #(.width(1)) bitwiseor_5724 (
        .y(_T_945),
        .a(cyc_A4),
        .b(cyc_A3_div)
    );
    wire _T_946;
    BITWISEOR #(.width(1)) bitwiseor_5725 (
        .y(_T_946),
        .a(_T_945),
        .b(cyc_A1_div)
    );
    wire _T_947;
    BITWISEOR #(.width(1)) bitwiseor_5726 (
        .y(_T_947),
        .a(_T_946),
        .b(cyc_B10_sqrt)
    );
    wire _T_948;
    BITWISEOR #(.width(1)) bitwiseor_5727 (
        .y(_T_948),
        .a(_T_947),
        .b(cyc_B9_sqrt)
    );
    wire _T_949;
    BITWISEOR #(.width(1)) bitwiseor_5728 (
        .y(_T_949),
        .a(_T_948),
        .b(cyc_B7_sqrt)
    );
    wire _T_950;
    BITWISEOR #(.width(1)) bitwiseor_5729 (
        .y(_T_950),
        .a(_T_949),
        .b(cyc_B6)
    );
    wire _T_951;
    BITWISEOR #(.width(1)) bitwiseor_5730 (
        .y(_T_951),
        .a(_T_950),
        .b(cyc_B5_sqrt)
    );
    wire _T_952;
    BITWISEOR #(.width(1)) bitwiseor_5731 (
        .y(_T_952),
        .a(_T_951),
        .b(cyc_B3_sqrt)
    );
    wire _T_953;
    BITWISEOR #(.width(1)) bitwiseor_5732 (
        .y(_T_953),
        .a(_T_952),
        .b(cyc_B2_div)
    );
    wire _T_954;
    BITWISEOR #(.width(1)) bitwiseor_5733 (
        .y(_T_954),
        .a(_T_953),
        .b(cyc_B1_sqrt)
    );
    wire _T_955;
    BITWISEOR #(.width(1)) bitwiseor_5734 (
        .y(_T_955),
        .a(_T_954),
        .b(cyc_C4)
    );
    wire _T_956;
    BITWISEOR #(.width(1)) bitwiseor_5735 (
        .y(_T_956),
        .a(cyc_A3),
        .b(cyc_A2_div)
    );
    wire _T_957;
    BITWISEOR #(.width(1)) bitwiseor_5736 (
        .y(_T_957),
        .a(_T_956),
        .b(cyc_B9_sqrt)
    );
    wire _T_958;
    BITWISEOR #(.width(1)) bitwiseor_5737 (
        .y(_T_958),
        .a(_T_957),
        .b(cyc_B8_sqrt)
    );
    wire _T_959;
    BITWISEOR #(.width(1)) bitwiseor_5738 (
        .y(_T_959),
        .a(_T_958),
        .b(cyc_B6)
    );
    wire _T_960;
    BITWISEOR #(.width(1)) bitwiseor_5739 (
        .y(_T_960),
        .a(_T_959),
        .b(cyc_B5)
    );
    wire _T_961;
    BITWISEOR #(.width(1)) bitwiseor_5740 (
        .y(_T_961),
        .a(_T_960),
        .b(cyc_B4_sqrt)
    );
    wire _T_962;
    BITWISEOR #(.width(1)) bitwiseor_5741 (
        .y(_T_962),
        .a(_T_961),
        .b(cyc_B2_sqrt)
    );
    wire _T_963;
    BITWISEOR #(.width(1)) bitwiseor_5742 (
        .y(_T_963),
        .a(_T_962),
        .b(cyc_B1_div)
    );
    wire _T_964;
    BITWISEOR #(.width(1)) bitwiseor_5743 (
        .y(_T_964),
        .a(_T_963),
        .b(cyc_C6_sqrt)
    );
    wire _T_965;
    BITWISEOR #(.width(1)) bitwiseor_5744 (
        .y(_T_965),
        .a(_T_964),
        .b(cyc_C3)
    );
    wire _T_966;
    BITWISEOR #(.width(1)) bitwiseor_5745 (
        .y(_T_966),
        .a(cyc_A2),
        .b(cyc_A1_div)
    );
    wire _T_967;
    BITWISEOR #(.width(1)) bitwiseor_5746 (
        .y(_T_967),
        .a(_T_966),
        .b(cyc_B8_sqrt)
    );
    wire _T_968;
    BITWISEOR #(.width(1)) bitwiseor_5747 (
        .y(_T_968),
        .a(_T_967),
        .b(cyc_B7_sqrt)
    );
    wire _T_969;
    BITWISEOR #(.width(1)) bitwiseor_5748 (
        .y(_T_969),
        .a(_T_968),
        .b(cyc_B5)
    );
    wire _T_970;
    BITWISEOR #(.width(1)) bitwiseor_5749 (
        .y(_T_970),
        .a(_T_969),
        .b(cyc_B4)
    );
    wire _T_971;
    BITWISEOR #(.width(1)) bitwiseor_5750 (
        .y(_T_971),
        .a(_T_970),
        .b(cyc_B3_sqrt)
    );
    wire _T_972;
    BITWISEOR #(.width(1)) bitwiseor_5751 (
        .y(_T_972),
        .a(_T_971),
        .b(cyc_B1_sqrt)
    );
    wire _T_973;
    BITWISEOR #(.width(1)) bitwiseor_5752 (
        .y(_T_973),
        .a(_T_972),
        .b(cyc_C5)
    );
    wire _T_974;
    BITWISEOR #(.width(1)) bitwiseor_5753 (
        .y(_T_974),
        .a(_T_973),
        .b(cyc_C2)
    );
    wire _T_975;
    BITWISEOR #(.width(1)) bitwiseor_5754 (
        .y(_T_975),
        .a(io_latchMulAddA_0),
        .b(cyc_B6)
    );
    wire _T_976;
    BITWISEOR #(.width(1)) bitwiseor_5755 (
        .y(_T_976),
        .a(_T_975),
        .b(cyc_B2_sqrt)
    );
    wire [1:0] _T_977;
    CAT #(.width_a(1), .width_b(1)) cat_5756 (
        .y(_T_977),
        .a(_T_974),
        .b(_T_976)
    );
    wire [1:0] _T_978;
    CAT #(.width_a(1), .width_b(1)) cat_5757 (
        .y(_T_978),
        .a(_T_955),
        .b(_T_965)
    );
    wire [3:0] _T_979;
    CAT #(.width_a(2), .width_b(2)) cat_5758 (
        .y(_T_979),
        .a(_T_978),
        .b(_T_977)
    );
    wire [104:0] _T_980;
    SHL_UNSIGNED #(.width(58), .n(47)) u_shl_5759 (
        .y(_T_980),
        .in(_sigX1_B__q)
    );
    wire [104:0] _T_982;
    wire [104:0] _WTEMP_822;
    PAD_UNSIGNED #(.width(1), .n(105)) u_pad_5760 (
        .y(_WTEMP_822),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(105)) u_mux_5761 (
        .y(_T_982),
        .sel(cyc_B1),
        .a(_T_980),
        .b(_WTEMP_822)
    );
    wire [103:0] _T_983;
    SHL_UNSIGNED #(.width(58), .n(46)) u_shl_5762 (
        .y(_T_983),
        .in(_sigX1_B__q)
    );
    wire [103:0] _T_985;
    wire [103:0] _WTEMP_823;
    PAD_UNSIGNED #(.width(1), .n(104)) u_pad_5763 (
        .y(_WTEMP_823),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(104)) u_mux_5764 (
        .y(_T_985),
        .sel(cyc_C6_sqrt),
        .a(_T_983),
        .b(_WTEMP_823)
    );
    wire [104:0] _T_986;
    wire [104:0] _WTEMP_824;
    PAD_UNSIGNED #(.width(104), .n(105)) u_pad_5765 (
        .y(_WTEMP_824),
        .in(_T_985)
    );
    BITWISEOR #(.width(105)) bitwiseor_5766 (
        .y(_T_986),
        .a(_T_982),
        .b(_WTEMP_824)
    );
    wire _T_987;
    BITWISEOR #(.width(1)) bitwiseor_5767 (
        .y(_T_987),
        .a(cyc_C4_sqrt),
        .b(cyc_C2)
    );
    wire [104:0] _T_988;
    SHL_UNSIGNED #(.width(58), .n(47)) u_shl_5768 (
        .y(_T_988),
        .in(_sigXN_C__q)
    );
    wire [104:0] _T_990;
    wire [104:0] _WTEMP_825;
    PAD_UNSIGNED #(.width(1), .n(105)) u_pad_5769 (
        .y(_WTEMP_825),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(105)) u_mux_5770 (
        .y(_T_990),
        .sel(_T_987),
        .a(_T_988),
        .b(_WTEMP_825)
    );
    wire [104:0] _T_991;
    BITWISEOR #(.width(105)) bitwiseor_5771 (
        .y(_T_991),
        .a(_T_986),
        .b(_T_990)
    );
    wire _T_993;
    EQ_UNSIGNED #(.width(1)) u_eq_5772 (
        .y(_T_993),
        .a(_E_E_div__q),
        .b(1'h0)
    );
    wire _T_994;
    BITWISEAND #(.width(1)) bitwiseand_5773 (
        .y(_T_994),
        .a(cyc_E3_div),
        .b(_T_993)
    );
    wire [53:0] _T_995;
    SHL_UNSIGNED #(.width(1), .n(53)) u_shl_5774 (
        .y(_T_995),
        .in(_fractA_0_PC__q)
    );
    wire [53:0] _T_997;
    wire [53:0] _WTEMP_826;
    PAD_UNSIGNED #(.width(1), .n(54)) u_pad_5775 (
        .y(_WTEMP_826),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(54)) u_mux_5776 (
        .y(_T_997),
        .sel(_T_994),
        .a(_T_995),
        .b(_WTEMP_826)
    );
    wire [104:0] _T_998;
    wire [104:0] _WTEMP_827;
    PAD_UNSIGNED #(.width(54), .n(105)) u_pad_5777 (
        .y(_WTEMP_827),
        .in(_T_997)
    );
    BITWISEOR #(.width(105)) bitwiseor_5778 (
        .y(_T_998),
        .a(_T_991),
        .b(_WTEMP_827)
    );
    wire _T_999;
    BITS #(.width(14), .high(0), .low(0)) bits_5779 (
        .y(_T_999),
        .in(_exp_PC__q)
    );
    wire _T_1000;
    BITS #(.width(53), .high(0), .low(0)) bits_5780 (
        .y(_T_1000),
        .in(sigB_PC)
    );
    wire [1:0] _T_1002;
    CAT #(.width_a(1), .width_b(1)) cat_5781 (
        .y(_T_1002),
        .a(_T_1000),
        .b(1'h0)
    );
    wire _T_1003;
    BITS #(.width(53), .high(1), .low(1)) bits_5782 (
        .y(_T_1003),
        .in(sigB_PC)
    );
    wire _T_1004;
    BITS #(.width(53), .high(0), .low(0)) bits_5783 (
        .y(_T_1004),
        .in(sigB_PC)
    );
    wire _T_1005;
    BITWISEXOR #(.width(1)) bitwisexor_5784 (
        .y(_T_1005),
        .a(_T_1003),
        .b(_T_1004)
    );
    wire _T_1006;
    BITS #(.width(53), .high(0), .low(0)) bits_5785 (
        .y(_T_1006),
        .in(sigB_PC)
    );
    wire [1:0] _T_1007;
    CAT #(.width_a(1), .width_b(1)) cat_5786 (
        .y(_T_1007),
        .a(_T_1005),
        .b(_T_1006)
    );
    wire [1:0] _T_1008;
    MUX_UNSIGNED #(.width(2)) u_mux_5787 (
        .y(_T_1008),
        .sel(_T_999),
        .a(_T_1002),
        .b(_T_1007)
    );
    wire _T_1010;
    EQ_UNSIGNED #(.width(1)) u_eq_5788 (
        .y(_T_1010),
        .a(_extraT_E__q),
        .b(1'h0)
    );
    wire [1:0] _T_1012;
    CAT #(.width_a(1), .width_b(1)) cat_5789 (
        .y(_T_1012),
        .a(_T_1010),
        .b(1'h0)
    );
    wire [1:0] _T_1013;
    BITWISEXOR #(.width(2)) bitwisexor_5790 (
        .y(_T_1013),
        .a(_T_1008),
        .b(_T_1012)
    );
    wire [55:0] _T_1014;
    SHL_UNSIGNED #(.width(2), .n(54)) u_shl_5791 (
        .y(_T_1014),
        .in(_T_1013)
    );
    wire [55:0] _T_1016;
    wire [55:0] _WTEMP_828;
    PAD_UNSIGNED #(.width(1), .n(56)) u_pad_5792 (
        .y(_WTEMP_828),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(56)) u_mux_5793 (
        .y(_T_1016),
        .sel(cyc_E3_sqrt),
        .a(_T_1014),
        .b(_WTEMP_828)
    );
    wire [104:0] _T_1017;
    wire [104:0] _WTEMP_829;
    PAD_UNSIGNED #(.width(56), .n(105)) u_pad_5794 (
        .y(_WTEMP_829),
        .in(_T_1016)
    );
    BITWISEOR #(.width(105)) bitwiseor_5795 (
        .y(_T_1017),
        .a(_T_998),
        .b(_WTEMP_829)
    );
    wire [31:0] ESqrR1_B8_sqrt;
    BITS #(.width(105), .high(103), .low(72)) bits_5796 (
        .y(ESqrR1_B8_sqrt),
        .in(io_mulAddResult_3)
    );
    wire [45:0] _T_1018;
    BITS #(.width(105), .high(90), .low(45)) bits_5797 (
        .y(_T_1018),
        .in(io_mulAddResult_3)
    );
    wire [45:0] _T_1019;
    BITWISENOT #(.width(46)) bitwisenot_5798 (
        .y(_T_1019),
        .in(_T_1018)
    );
    wire [45:0] _T_1021;
    wire [45:0] _WTEMP_830;
    PAD_UNSIGNED #(.width(1), .n(46)) u_pad_5799 (
        .y(_WTEMP_830),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(46)) u_mux_5800 (
        .y(_T_1021),
        .sel(cyc_B4),
        .a(_T_1019),
        .b(_WTEMP_830)
    );
    wire [32:0] sqrSigma1_B1;
    BITS #(.width(105), .high(79), .low(47)) bits_5801 (
        .y(sqrSigma1_B1),
        .in(io_mulAddResult_3)
    );
    wire [57:0] _T_1022;
    BITS #(.width(105), .high(104), .low(47)) bits_5802 (
        .y(_T_1022),
        .in(io_mulAddResult_3)
    );
    wire _T_1023;
    BITS #(.width(105), .high(104), .low(104)) bits_5803 (
        .y(_T_1023),
        .in(io_mulAddResult_3)
    );
    wire E_C1_div;
    EQ_UNSIGNED #(.width(1)) u_eq_5804 (
        .y(E_C1_div),
        .a(_T_1023),
        .b(1'h0)
    );
    wire _T_1026;
    EQ_UNSIGNED #(.width(1)) u_eq_5805 (
        .y(_T_1026),
        .a(E_C1_div),
        .b(1'h0)
    );
    wire _T_1027;
    BITWISEAND #(.width(1)) bitwiseand_5806 (
        .y(_T_1027),
        .a(cyc_C1_div),
        .b(_T_1026)
    );
    wire _T_1028;
    BITWISEOR #(.width(1)) bitwiseor_5807 (
        .y(_T_1028),
        .a(_T_1027),
        .b(cyc_C1_sqrt)
    );
    wire [53:0] _T_1029;
    BITS #(.width(105), .high(104), .low(51)) bits_5808 (
        .y(_T_1029),
        .in(io_mulAddResult_3)
    );
    wire [53:0] _T_1030;
    BITWISENOT #(.width(54)) bitwisenot_5809 (
        .y(_T_1030),
        .in(_T_1029)
    );
    wire [53:0] _T_1032;
    wire [53:0] _WTEMP_831;
    PAD_UNSIGNED #(.width(1), .n(54)) u_pad_5810 (
        .y(_WTEMP_831),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(54)) u_mux_5811 (
        .y(_T_1032),
        .sel(_T_1028),
        .a(_T_1030),
        .b(_WTEMP_831)
    );
    wire _T_1033;
    BITWISEAND #(.width(1)) bitwiseand_5812 (
        .y(_T_1033),
        .a(cyc_C1_div),
        .b(E_C1_div)
    );
    wire [52:0] _T_1035;
    BITS #(.width(105), .high(102), .low(50)) bits_5813 (
        .y(_T_1035),
        .in(io_mulAddResult_3)
    );
    wire [52:0] _T_1036;
    BITWISENOT #(.width(53)) bitwisenot_5814 (
        .y(_T_1036),
        .in(_T_1035)
    );
    wire [53:0] _T_1037;
    CAT #(.width_a(1), .width_b(53)) cat_5815 (
        .y(_T_1037),
        .a(1'h0),
        .b(_T_1036)
    );
    wire [53:0] _T_1039;
    wire [53:0] _WTEMP_832;
    PAD_UNSIGNED #(.width(1), .n(54)) u_pad_5816 (
        .y(_WTEMP_832),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(54)) u_mux_5817 (
        .y(_T_1039),
        .sel(_T_1033),
        .a(_T_1037),
        .b(_WTEMP_832)
    );
    wire [53:0] _T_1040;
    BITWISEOR #(.width(54)) bitwiseor_5818 (
        .y(_T_1040),
        .a(_T_1032),
        .b(_T_1039)
    );
    wire [53:0] _T_1041;
    BITS #(.width(105), .high(104), .low(51)) bits_5819 (
        .y(_T_1041),
        .in(io_mulAddResult_3)
    );
    wire [53:0] _T_1042;
    BITWISENOT #(.width(54)) bitwisenot_5820 (
        .y(_T_1042),
        .in(_T_1041)
    );
    wire [53:0] _T_1044;
    wire [53:0] _WTEMP_833;
    PAD_UNSIGNED #(.width(1), .n(54)) u_pad_5821 (
        .y(_WTEMP_833),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(54)) u_mux_5822 (
        .y(_T_1044),
        .sel(cyc_C1_sqrt),
        .a(_T_1042),
        .b(_WTEMP_833)
    );
    wire [53:0] sigT_C1;
    BITWISENOT #(.width(54)) bitwisenot_5823 (
        .y(sigT_C1),
        .in(zComplSigT_C1)
    );
    wire [55:0] remT_E2;
    BITS #(.width(105), .high(55), .low(0)) bits_5824 (
        .y(remT_E2),
        .in(io_mulAddResult_3)
    );
    wire _T_1045;
    BITWISEOR #(.width(1)) bitwiseor_5825 (
        .y(_T_1045),
        .a(cyc_C6_sqrt),
        .b(cyc_C5_div)
    );
    wire _T_1046;
    BITWISEOR #(.width(1)) bitwiseor_5826 (
        .y(_T_1046),
        .a(_T_1045),
        .b(cyc_C3_sqrt)
    );
    wire [30:0] _T_1047;
    BITS #(.width(58), .high(56), .low(26)) bits_5827 (
        .y(_T_1047),
        .in(sigXNU_B3_CX)
    );
    wire [52:0] _T_1048;
    BITS #(.width(54), .high(53), .low(1)) bits_5828 (
        .y(_T_1048),
        .in(sigT_C1)
    );
    wire _T_1049;
    BITS #(.width(54), .high(0), .low(0)) bits_5829 (
        .y(_T_1049),
        .in(sigT_C1)
    );
    wire _T_1050;
    BITS #(.width(56), .high(55), .low(55)) bits_5830 (
        .y(_T_1050),
        .in(remT_E2)
    );
    wire _T_1051;
    BITS #(.width(56), .high(53), .low(53)) bits_5831 (
        .y(_T_1051),
        .in(remT_E2)
    );
    wire _T_1052;
    MUX_UNSIGNED #(.width(1)) u_mux_5832 (
        .y(_T_1052),
        .sel(_sqrtOp_PC__q),
        .a(_T_1050),
        .b(_T_1051)
    );
    wire [53:0] _T_1053;
    BITS #(.width(56), .high(53), .low(0)) bits_5833 (
        .y(_T_1053),
        .in(remT_E2)
    );
    wire _T_1055;
    wire [53:0] _WTEMP_834;
    PAD_UNSIGNED #(.width(1), .n(54)) u_pad_5834 (
        .y(_WTEMP_834),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(54)) u_eq_5835 (
        .y(_T_1055),
        .a(_T_1053),
        .b(_WTEMP_834)
    );
    wire _T_1057;
    EQ_UNSIGNED #(.width(1)) u_eq_5836 (
        .y(_T_1057),
        .a(_sqrtOp_PC__q),
        .b(1'h0)
    );
    wire [1:0] _T_1058;
    BITS #(.width(56), .high(55), .low(54)) bits_5837 (
        .y(_T_1058),
        .in(remT_E2)
    );
    wire _T_1060;
    wire [1:0] _WTEMP_835;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_5838 (
        .y(_WTEMP_835),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(2)) u_eq_5839 (
        .y(_T_1060),
        .a(_T_1058),
        .b(_WTEMP_835)
    );
    wire _T_1061;
    BITWISEOR #(.width(1)) bitwiseor_5840 (
        .y(_T_1061),
        .a(_T_1057),
        .b(_T_1060)
    );
    wire _T_1062;
    BITWISEAND #(.width(1)) bitwiseand_5841 (
        .y(_T_1062),
        .a(_T_1055),
        .b(_T_1061)
    );
    wire _T_1064;
    EQ_UNSIGNED #(.width(1)) u_eq_5842 (
        .y(_T_1064),
        .a(_sqrtOp_PC__q),
        .b(1'h0)
    );
    wire _T_1065;
    BITWISEAND #(.width(1)) bitwiseand_5843 (
        .y(_T_1065),
        .a(_T_1064),
        .b(_E_E_div__q)
    );
    wire [13:0] _T_1067;
    wire [13:0] _WTEMP_836;
    PAD_UNSIGNED #(.width(1), .n(14)) u_pad_5844 (
        .y(_WTEMP_836),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(14)) u_mux_5845 (
        .y(_T_1067),
        .sel(_T_1065),
        .a(_exp_PC__q),
        .b(_WTEMP_836)
    );
    wire _T_1069;
    EQ_UNSIGNED #(.width(1)) u_eq_5846 (
        .y(_T_1069),
        .a(_sqrtOp_PC__q),
        .b(1'h0)
    );
    wire _T_1071;
    EQ_UNSIGNED #(.width(1)) u_eq_5847 (
        .y(_T_1071),
        .a(_E_E_div__q),
        .b(1'h0)
    );
    wire _T_1072;
    BITWISEAND #(.width(1)) bitwiseand_5848 (
        .y(_T_1072),
        .a(_T_1069),
        .b(_T_1071)
    );
    wire [13:0] _T_1074;
    wire [13:0] _WTEMP_837;
    PAD_UNSIGNED #(.width(1), .n(14)) u_pad_5849 (
        .y(_WTEMP_837),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(14)) u_mux_5850 (
        .y(_T_1074),
        .sel(_T_1072),
        .a(expP1_PC),
        .b(_WTEMP_837)
    );
    wire [13:0] _T_1075;
    BITWISEOR #(.width(14)) bitwiseor_5851 (
        .y(_T_1075),
        .a(_T_1067),
        .b(_T_1074)
    );
    wire [12:0] _T_1076;
    SHR_UNSIGNED #(.width(14), .n(1)) u_shr_5852 (
        .y(_T_1076),
        .in(_exp_PC__q)
    );
    wire [13:0] _T_1078;
    wire [12:0] _WTEMP_838;
    PAD_UNSIGNED #(.width(12), .n(13)) u_pad_5853 (
        .y(_WTEMP_838),
        .in(12'h400)
    );
    ADD_UNSIGNED #(.width(13)) u_add_5854 (
        .y(_T_1078),
        .a(_T_1076),
        .b(_WTEMP_838)
    );
    wire [12:0] _T_1079;
    TAIL #(.width(14), .n(1)) tail_5855 (
        .y(_T_1079),
        .in(_T_1078)
    );
    wire [12:0] _T_1081;
    wire [12:0] _WTEMP_839;
    PAD_UNSIGNED #(.width(1), .n(13)) u_pad_5856 (
        .y(_WTEMP_839),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(13)) u_mux_5857 (
        .y(_T_1081),
        .sel(_sqrtOp_PC__q),
        .a(_T_1079),
        .b(_WTEMP_839)
    );
    wire [13:0] sExpX_E;
    wire [13:0] _WTEMP_840;
    PAD_UNSIGNED #(.width(13), .n(14)) u_pad_5858 (
        .y(_WTEMP_840),
        .in(_T_1081)
    );
    BITWISEOR #(.width(14)) bitwiseor_5859 (
        .y(sExpX_E),
        .a(_T_1075),
        .b(_WTEMP_840)
    );
    wire [12:0] posExpX_E;
    BITS #(.width(14), .high(12), .low(0)) bits_5860 (
        .y(posExpX_E),
        .in(sExpX_E)
    );
    wire [12:0] _T_1082;
    BITWISENOT #(.width(13)) bitwisenot_5861 (
        .y(_T_1082),
        .in(posExpX_E)
    );
    wire _T_1083;
    BITS #(.width(13), .high(12), .low(12)) bits_5862 (
        .y(_T_1083),
        .in(_T_1082)
    );
    wire [11:0] _T_1084;
    BITS #(.width(13), .high(11), .low(0)) bits_5863 (
        .y(_T_1084),
        .in(_T_1082)
    );
    wire _T_1085;
    BITS #(.width(12), .high(11), .low(11)) bits_5864 (
        .y(_T_1085),
        .in(_T_1084)
    );
    wire [10:0] _T_1086;
    BITS #(.width(12), .high(10), .low(0)) bits_5865 (
        .y(_T_1086),
        .in(_T_1084)
    );
    wire _T_1087;
    BITS #(.width(11), .high(10), .low(10)) bits_5866 (
        .y(_T_1087),
        .in(_T_1086)
    );
    wire [9:0] _T_1088;
    BITS #(.width(11), .high(9), .low(0)) bits_5867 (
        .y(_T_1088),
        .in(_T_1086)
    );
    wire _T_1089;
    BITS #(.width(10), .high(9), .low(9)) bits_5868 (
        .y(_T_1089),
        .in(_T_1088)
    );
    wire [8:0] _T_1090;
    BITS #(.width(10), .high(8), .low(0)) bits_5869 (
        .y(_T_1090),
        .in(_T_1088)
    );
    wire _T_1092;
    BITS #(.width(9), .high(8), .low(8)) bits_5870 (
        .y(_T_1092),
        .in(_T_1090)
    );
    wire [7:0] _T_1093;
    BITS #(.width(9), .high(7), .low(0)) bits_5871 (
        .y(_T_1093),
        .in(_T_1090)
    );
    wire _T_1095;
    BITS #(.width(8), .high(7), .low(7)) bits_5872 (
        .y(_T_1095),
        .in(_T_1093)
    );
    wire [6:0] _T_1096;
    BITS #(.width(8), .high(6), .low(0)) bits_5873 (
        .y(_T_1096),
        .in(_T_1093)
    );
    wire _T_1098;
    BITS #(.width(7), .high(6), .low(6)) bits_5874 (
        .y(_T_1098),
        .in(_T_1096)
    );
    wire [5:0] _T_1099;
    BITS #(.width(7), .high(5), .low(0)) bits_5875 (
        .y(_T_1099),
        .in(_T_1096)
    );
    wire [64:0] _T_1102;
    DSHR_SIGNED #(.width_in(65), .width_n(6)) s_dshr_5876 (
        .y(_T_1102),
        .in(-65'sh10000000000000000),
        .n(_T_1099)
    );
    wire [49:0] _T_1103;
    BITS #(.width(65), .high(63), .low(14)) bits_5877 (
        .y(_T_1103),
        .in(_T_1102)
    );
    wire [31:0] _T_1104;
    BITS #(.width(50), .high(31), .low(0)) bits_5878 (
        .y(_T_1104),
        .in(_T_1103)
    );
    wire [31:0] _T_1107;
    assign _T_1107 = 32'hFFFF0000;
    wire [31:0] _T_1108;
    assign _T_1108 = 32'hFFFF;
    wire [15:0] _T_1109;
    SHR_UNSIGNED #(.width(32), .n(16)) u_shr_5879 (
        .y(_T_1109),
        .in(_T_1104)
    );
    wire [31:0] _T_1110;
    wire [31:0] _WTEMP_841;
    PAD_UNSIGNED #(.width(16), .n(32)) u_pad_5880 (
        .y(_WTEMP_841),
        .in(_T_1109)
    );
    BITWISEAND #(.width(32)) bitwiseand_5881 (
        .y(_T_1110),
        .a(_WTEMP_841),
        .b(_T_1108)
    );
    wire [15:0] _T_1111;
    BITS #(.width(32), .high(15), .low(0)) bits_5882 (
        .y(_T_1111),
        .in(_T_1104)
    );
    wire [31:0] _T_1112;
    SHL_UNSIGNED #(.width(16), .n(16)) u_shl_5883 (
        .y(_T_1112),
        .in(_T_1111)
    );
    wire [31:0] _T_1113;
    assign _T_1113 = 32'hFFFF0000;
    wire [31:0] _T_1114;
    BITWISEAND #(.width(32)) bitwiseand_5884 (
        .y(_T_1114),
        .a(_T_1112),
        .b(_T_1113)
    );
    wire [31:0] _T_1115;
    BITWISEOR #(.width(32)) bitwiseor_5885 (
        .y(_T_1115),
        .a(_T_1110),
        .b(_T_1114)
    );
    wire [23:0] _T_1116;
    assign _T_1116 = 24'hFFFF;
    wire [31:0] _T_1117;
    assign _T_1117 = 32'hFFFF00;
    wire [31:0] _T_1118;
    assign _T_1118 = 32'hFF00FF;
    wire [23:0] _T_1119;
    SHR_UNSIGNED #(.width(32), .n(8)) u_shr_5886 (
        .y(_T_1119),
        .in(_T_1115)
    );
    wire [31:0] _T_1120;
    wire [31:0] _WTEMP_842;
    PAD_UNSIGNED #(.width(24), .n(32)) u_pad_5887 (
        .y(_WTEMP_842),
        .in(_T_1119)
    );
    BITWISEAND #(.width(32)) bitwiseand_5888 (
        .y(_T_1120),
        .a(_WTEMP_842),
        .b(_T_1118)
    );
    wire [23:0] _T_1121;
    BITS #(.width(32), .high(23), .low(0)) bits_5889 (
        .y(_T_1121),
        .in(_T_1115)
    );
    wire [31:0] _T_1122;
    SHL_UNSIGNED #(.width(24), .n(8)) u_shl_5890 (
        .y(_T_1122),
        .in(_T_1121)
    );
    wire [31:0] _T_1123;
    assign _T_1123 = 32'hFF00FF00;
    wire [31:0] _T_1124;
    BITWISEAND #(.width(32)) bitwiseand_5891 (
        .y(_T_1124),
        .a(_T_1122),
        .b(_T_1123)
    );
    wire [31:0] _T_1125;
    BITWISEOR #(.width(32)) bitwiseor_5892 (
        .y(_T_1125),
        .a(_T_1120),
        .b(_T_1124)
    );
    wire [27:0] _T_1126;
    assign _T_1126 = 28'hFF00FF;
    wire [31:0] _T_1127;
    assign _T_1127 = 32'hFF00FF0;
    wire [31:0] _T_1128;
    assign _T_1128 = 32'hF0F0F0F;
    wire [27:0] _T_1129;
    SHR_UNSIGNED #(.width(32), .n(4)) u_shr_5893 (
        .y(_T_1129),
        .in(_T_1125)
    );
    wire [31:0] _T_1130;
    wire [31:0] _WTEMP_843;
    PAD_UNSIGNED #(.width(28), .n(32)) u_pad_5894 (
        .y(_WTEMP_843),
        .in(_T_1129)
    );
    BITWISEAND #(.width(32)) bitwiseand_5895 (
        .y(_T_1130),
        .a(_WTEMP_843),
        .b(_T_1128)
    );
    wire [27:0] _T_1131;
    BITS #(.width(32), .high(27), .low(0)) bits_5896 (
        .y(_T_1131),
        .in(_T_1125)
    );
    wire [31:0] _T_1132;
    SHL_UNSIGNED #(.width(28), .n(4)) u_shl_5897 (
        .y(_T_1132),
        .in(_T_1131)
    );
    wire [31:0] _T_1133;
    assign _T_1133 = 32'hF0F0F0F0;
    wire [31:0] _T_1134;
    BITWISEAND #(.width(32)) bitwiseand_5898 (
        .y(_T_1134),
        .a(_T_1132),
        .b(_T_1133)
    );
    wire [31:0] _T_1135;
    BITWISEOR #(.width(32)) bitwiseor_5899 (
        .y(_T_1135),
        .a(_T_1130),
        .b(_T_1134)
    );
    wire [29:0] _T_1136;
    assign _T_1136 = 30'hF0F0F0F;
    wire [31:0] _T_1137;
    assign _T_1137 = 32'h3C3C3C3C;
    wire [31:0] _T_1138;
    assign _T_1138 = 32'h33333333;
    wire [29:0] _T_1139;
    SHR_UNSIGNED #(.width(32), .n(2)) u_shr_5900 (
        .y(_T_1139),
        .in(_T_1135)
    );
    wire [31:0] _T_1140;
    wire [31:0] _WTEMP_844;
    PAD_UNSIGNED #(.width(30), .n(32)) u_pad_5901 (
        .y(_WTEMP_844),
        .in(_T_1139)
    );
    BITWISEAND #(.width(32)) bitwiseand_5902 (
        .y(_T_1140),
        .a(_WTEMP_844),
        .b(_T_1138)
    );
    wire [29:0] _T_1141;
    BITS #(.width(32), .high(29), .low(0)) bits_5903 (
        .y(_T_1141),
        .in(_T_1135)
    );
    wire [31:0] _T_1142;
    SHL_UNSIGNED #(.width(30), .n(2)) u_shl_5904 (
        .y(_T_1142),
        .in(_T_1141)
    );
    wire [31:0] _T_1143;
    assign _T_1143 = 32'hCCCCCCCC;
    wire [31:0] _T_1144;
    BITWISEAND #(.width(32)) bitwiseand_5905 (
        .y(_T_1144),
        .a(_T_1142),
        .b(_T_1143)
    );
    wire [31:0] _T_1145;
    BITWISEOR #(.width(32)) bitwiseor_5906 (
        .y(_T_1145),
        .a(_T_1140),
        .b(_T_1144)
    );
    wire [30:0] _T_1146;
    assign _T_1146 = 31'h33333333;
    wire [31:0] _T_1147;
    assign _T_1147 = 32'h66666666;
    wire [31:0] _T_1148;
    assign _T_1148 = 32'h55555555;
    wire [30:0] _T_1149;
    SHR_UNSIGNED #(.width(32), .n(1)) u_shr_5907 (
        .y(_T_1149),
        .in(_T_1145)
    );
    wire [31:0] _T_1150;
    wire [31:0] _WTEMP_845;
    PAD_UNSIGNED #(.width(31), .n(32)) u_pad_5908 (
        .y(_WTEMP_845),
        .in(_T_1149)
    );
    BITWISEAND #(.width(32)) bitwiseand_5909 (
        .y(_T_1150),
        .a(_WTEMP_845),
        .b(_T_1148)
    );
    wire [30:0] _T_1151;
    BITS #(.width(32), .high(30), .low(0)) bits_5910 (
        .y(_T_1151),
        .in(_T_1145)
    );
    wire [31:0] _T_1152;
    SHL_UNSIGNED #(.width(31), .n(1)) u_shl_5911 (
        .y(_T_1152),
        .in(_T_1151)
    );
    wire [31:0] _T_1153;
    assign _T_1153 = 32'hAAAAAAAA;
    wire [31:0] _T_1154;
    BITWISEAND #(.width(32)) bitwiseand_5912 (
        .y(_T_1154),
        .a(_T_1152),
        .b(_T_1153)
    );
    wire [31:0] _T_1155;
    BITWISEOR #(.width(32)) bitwiseor_5913 (
        .y(_T_1155),
        .a(_T_1150),
        .b(_T_1154)
    );
    wire [17:0] _T_1156;
    BITS #(.width(50), .high(49), .low(32)) bits_5914 (
        .y(_T_1156),
        .in(_T_1103)
    );
    wire [15:0] _T_1157;
    BITS #(.width(18), .high(15), .low(0)) bits_5915 (
        .y(_T_1157),
        .in(_T_1156)
    );
    wire [15:0] _T_1160;
    assign _T_1160 = 16'hFF00;
    wire [15:0] _T_1161;
    assign _T_1161 = 16'hFF;
    wire [7:0] _T_1162;
    SHR_UNSIGNED #(.width(16), .n(8)) u_shr_5916 (
        .y(_T_1162),
        .in(_T_1157)
    );
    wire [15:0] _T_1163;
    wire [15:0] _WTEMP_846;
    PAD_UNSIGNED #(.width(8), .n(16)) u_pad_5917 (
        .y(_WTEMP_846),
        .in(_T_1162)
    );
    BITWISEAND #(.width(16)) bitwiseand_5918 (
        .y(_T_1163),
        .a(_WTEMP_846),
        .b(_T_1161)
    );
    wire [7:0] _T_1164;
    BITS #(.width(16), .high(7), .low(0)) bits_5919 (
        .y(_T_1164),
        .in(_T_1157)
    );
    wire [15:0] _T_1165;
    SHL_UNSIGNED #(.width(8), .n(8)) u_shl_5920 (
        .y(_T_1165),
        .in(_T_1164)
    );
    wire [15:0] _T_1166;
    assign _T_1166 = 16'hFF00;
    wire [15:0] _T_1167;
    BITWISEAND #(.width(16)) bitwiseand_5921 (
        .y(_T_1167),
        .a(_T_1165),
        .b(_T_1166)
    );
    wire [15:0] _T_1168;
    BITWISEOR #(.width(16)) bitwiseor_5922 (
        .y(_T_1168),
        .a(_T_1163),
        .b(_T_1167)
    );
    wire [11:0] _T_1169;
    assign _T_1169 = 12'hFF;
    wire [15:0] _T_1170;
    assign _T_1170 = 16'hFF0;
    wire [15:0] _T_1171;
    assign _T_1171 = 16'hF0F;
    wire [11:0] _T_1172;
    SHR_UNSIGNED #(.width(16), .n(4)) u_shr_5923 (
        .y(_T_1172),
        .in(_T_1168)
    );
    wire [15:0] _T_1173;
    wire [15:0] _WTEMP_847;
    PAD_UNSIGNED #(.width(12), .n(16)) u_pad_5924 (
        .y(_WTEMP_847),
        .in(_T_1172)
    );
    BITWISEAND #(.width(16)) bitwiseand_5925 (
        .y(_T_1173),
        .a(_WTEMP_847),
        .b(_T_1171)
    );
    wire [11:0] _T_1174;
    BITS #(.width(16), .high(11), .low(0)) bits_5926 (
        .y(_T_1174),
        .in(_T_1168)
    );
    wire [15:0] _T_1175;
    SHL_UNSIGNED #(.width(12), .n(4)) u_shl_5927 (
        .y(_T_1175),
        .in(_T_1174)
    );
    wire [15:0] _T_1176;
    assign _T_1176 = 16'hF0F0;
    wire [15:0] _T_1177;
    BITWISEAND #(.width(16)) bitwiseand_5928 (
        .y(_T_1177),
        .a(_T_1175),
        .b(_T_1176)
    );
    wire [15:0] _T_1178;
    BITWISEOR #(.width(16)) bitwiseor_5929 (
        .y(_T_1178),
        .a(_T_1173),
        .b(_T_1177)
    );
    wire [13:0] _T_1179;
    assign _T_1179 = 14'hF0F;
    wire [15:0] _T_1180;
    assign _T_1180 = 16'h3C3C;
    wire [15:0] _T_1181;
    assign _T_1181 = 16'h3333;
    wire [13:0] _T_1182;
    SHR_UNSIGNED #(.width(16), .n(2)) u_shr_5930 (
        .y(_T_1182),
        .in(_T_1178)
    );
    wire [15:0] _T_1183;
    wire [15:0] _WTEMP_848;
    PAD_UNSIGNED #(.width(14), .n(16)) u_pad_5931 (
        .y(_WTEMP_848),
        .in(_T_1182)
    );
    BITWISEAND #(.width(16)) bitwiseand_5932 (
        .y(_T_1183),
        .a(_WTEMP_848),
        .b(_T_1181)
    );
    wire [13:0] _T_1184;
    BITS #(.width(16), .high(13), .low(0)) bits_5933 (
        .y(_T_1184),
        .in(_T_1178)
    );
    wire [15:0] _T_1185;
    SHL_UNSIGNED #(.width(14), .n(2)) u_shl_5934 (
        .y(_T_1185),
        .in(_T_1184)
    );
    wire [15:0] _T_1186;
    assign _T_1186 = 16'hCCCC;
    wire [15:0] _T_1187;
    BITWISEAND #(.width(16)) bitwiseand_5935 (
        .y(_T_1187),
        .a(_T_1185),
        .b(_T_1186)
    );
    wire [15:0] _T_1188;
    BITWISEOR #(.width(16)) bitwiseor_5936 (
        .y(_T_1188),
        .a(_T_1183),
        .b(_T_1187)
    );
    wire [14:0] _T_1189;
    assign _T_1189 = 15'h3333;
    wire [15:0] _T_1190;
    assign _T_1190 = 16'h6666;
    wire [15:0] _T_1191;
    assign _T_1191 = 16'h5555;
    wire [14:0] _T_1192;
    SHR_UNSIGNED #(.width(16), .n(1)) u_shr_5937 (
        .y(_T_1192),
        .in(_T_1188)
    );
    wire [15:0] _T_1193;
    wire [15:0] _WTEMP_849;
    PAD_UNSIGNED #(.width(15), .n(16)) u_pad_5938 (
        .y(_WTEMP_849),
        .in(_T_1192)
    );
    BITWISEAND #(.width(16)) bitwiseand_5939 (
        .y(_T_1193),
        .a(_WTEMP_849),
        .b(_T_1191)
    );
    wire [14:0] _T_1194;
    BITS #(.width(16), .high(14), .low(0)) bits_5940 (
        .y(_T_1194),
        .in(_T_1188)
    );
    wire [15:0] _T_1195;
    SHL_UNSIGNED #(.width(15), .n(1)) u_shl_5941 (
        .y(_T_1195),
        .in(_T_1194)
    );
    wire [15:0] _T_1196;
    assign _T_1196 = 16'hAAAA;
    wire [15:0] _T_1197;
    BITWISEAND #(.width(16)) bitwiseand_5942 (
        .y(_T_1197),
        .a(_T_1195),
        .b(_T_1196)
    );
    wire [15:0] _T_1198;
    BITWISEOR #(.width(16)) bitwiseor_5943 (
        .y(_T_1198),
        .a(_T_1193),
        .b(_T_1197)
    );
    wire [1:0] _T_1199;
    BITS #(.width(18), .high(17), .low(16)) bits_5944 (
        .y(_T_1199),
        .in(_T_1156)
    );
    wire _T_1200;
    BITS #(.width(2), .high(0), .low(0)) bits_5945 (
        .y(_T_1200),
        .in(_T_1199)
    );
    wire _T_1201;
    BITS #(.width(2), .high(1), .low(1)) bits_5946 (
        .y(_T_1201),
        .in(_T_1199)
    );
    wire [1:0] _T_1202;
    CAT #(.width_a(1), .width_b(1)) cat_5947 (
        .y(_T_1202),
        .a(_T_1200),
        .b(_T_1201)
    );
    wire [17:0] _T_1203;
    CAT #(.width_a(16), .width_b(2)) cat_5948 (
        .y(_T_1203),
        .a(_T_1198),
        .b(_T_1202)
    );
    wire [49:0] _T_1204;
    CAT #(.width_a(32), .width_b(18)) cat_5949 (
        .y(_T_1204),
        .a(_T_1155),
        .b(_T_1203)
    );
    wire [49:0] _T_1205;
    BITWISENOT #(.width(50)) bitwisenot_5950 (
        .y(_T_1205),
        .in(_T_1204)
    );
    wire [49:0] _T_1206;
    wire [49:0] _WTEMP_850;
    PAD_UNSIGNED #(.width(1), .n(50)) u_pad_5951 (
        .y(_WTEMP_850),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(50)) u_mux_5952 (
        .y(_T_1206),
        .sel(_T_1098),
        .a(_WTEMP_850),
        .b(_T_1205)
    );
    wire [49:0] _T_1207;
    BITWISENOT #(.width(50)) bitwisenot_5953 (
        .y(_T_1207),
        .in(_T_1206)
    );
    wire [49:0] _T_1208;
    BITWISENOT #(.width(50)) bitwisenot_5954 (
        .y(_T_1208),
        .in(_T_1207)
    );
    wire [49:0] _T_1209;
    wire [49:0] _WTEMP_851;
    PAD_UNSIGNED #(.width(1), .n(50)) u_pad_5955 (
        .y(_WTEMP_851),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(50)) u_mux_5956 (
        .y(_T_1209),
        .sel(_T_1095),
        .a(_WTEMP_851),
        .b(_T_1208)
    );
    wire [49:0] _T_1210;
    BITWISENOT #(.width(50)) bitwisenot_5957 (
        .y(_T_1210),
        .in(_T_1209)
    );
    wire [49:0] _T_1211;
    BITWISENOT #(.width(50)) bitwisenot_5958 (
        .y(_T_1211),
        .in(_T_1210)
    );
    wire [49:0] _T_1212;
    wire [49:0] _WTEMP_852;
    PAD_UNSIGNED #(.width(1), .n(50)) u_pad_5959 (
        .y(_WTEMP_852),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(50)) u_mux_5960 (
        .y(_T_1212),
        .sel(_T_1092),
        .a(_WTEMP_852),
        .b(_T_1211)
    );
    wire [49:0] _T_1213;
    BITWISENOT #(.width(50)) bitwisenot_5961 (
        .y(_T_1213),
        .in(_T_1212)
    );
    wire [49:0] _T_1214;
    BITWISENOT #(.width(50)) bitwisenot_5962 (
        .y(_T_1214),
        .in(_T_1213)
    );
    wire [49:0] _T_1215;
    wire [49:0] _WTEMP_853;
    PAD_UNSIGNED #(.width(1), .n(50)) u_pad_5963 (
        .y(_WTEMP_853),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(50)) u_mux_5964 (
        .y(_T_1215),
        .sel(_T_1089),
        .a(_WTEMP_853),
        .b(_T_1214)
    );
    wire [49:0] _T_1216;
    BITWISENOT #(.width(50)) bitwisenot_5965 (
        .y(_T_1216),
        .in(_T_1215)
    );
    wire [52:0] _T_1218;
    CAT #(.width_a(50), .width_b(3)) cat_5966 (
        .y(_T_1218),
        .a(_T_1216),
        .b(3'h7)
    );
    wire _T_1219;
    BITS #(.width(10), .high(9), .low(9)) bits_5967 (
        .y(_T_1219),
        .in(_T_1088)
    );
    wire [8:0] _T_1220;
    BITS #(.width(10), .high(8), .low(0)) bits_5968 (
        .y(_T_1220),
        .in(_T_1088)
    );
    wire _T_1221;
    BITS #(.width(9), .high(8), .low(8)) bits_5969 (
        .y(_T_1221),
        .in(_T_1220)
    );
    wire [7:0] _T_1222;
    BITS #(.width(9), .high(7), .low(0)) bits_5970 (
        .y(_T_1222),
        .in(_T_1220)
    );
    wire _T_1223;
    BITS #(.width(8), .high(7), .low(7)) bits_5971 (
        .y(_T_1223),
        .in(_T_1222)
    );
    wire [6:0] _T_1224;
    BITS #(.width(8), .high(6), .low(0)) bits_5972 (
        .y(_T_1224),
        .in(_T_1222)
    );
    wire _T_1225;
    BITS #(.width(7), .high(6), .low(6)) bits_5973 (
        .y(_T_1225),
        .in(_T_1224)
    );
    wire [5:0] _T_1226;
    BITS #(.width(7), .high(5), .low(0)) bits_5974 (
        .y(_T_1226),
        .in(_T_1224)
    );
    wire [64:0] _T_1228;
    DSHR_SIGNED #(.width_in(65), .width_n(6)) s_dshr_5975 (
        .y(_T_1228),
        .in(-65'sh10000000000000000),
        .n(_T_1226)
    );
    wire [2:0] _T_1229;
    BITS #(.width(65), .high(2), .low(0)) bits_5976 (
        .y(_T_1229),
        .in(_T_1228)
    );
    wire [1:0] _T_1230;
    BITS #(.width(3), .high(1), .low(0)) bits_5977 (
        .y(_T_1230),
        .in(_T_1229)
    );
    wire _T_1231;
    BITS #(.width(2), .high(0), .low(0)) bits_5978 (
        .y(_T_1231),
        .in(_T_1230)
    );
    wire _T_1232;
    BITS #(.width(2), .high(1), .low(1)) bits_5979 (
        .y(_T_1232),
        .in(_T_1230)
    );
    wire [1:0] _T_1233;
    CAT #(.width_a(1), .width_b(1)) cat_5980 (
        .y(_T_1233),
        .a(_T_1231),
        .b(_T_1232)
    );
    wire _T_1234;
    BITS #(.width(3), .high(2), .low(2)) bits_5981 (
        .y(_T_1234),
        .in(_T_1229)
    );
    wire [2:0] _T_1235;
    CAT #(.width_a(2), .width_b(1)) cat_5982 (
        .y(_T_1235),
        .a(_T_1233),
        .b(_T_1234)
    );
    wire [2:0] _T_1237;
    wire [2:0] _WTEMP_854;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_5983 (
        .y(_WTEMP_854),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(3)) u_mux_5984 (
        .y(_T_1237),
        .sel(_T_1225),
        .a(_T_1235),
        .b(_WTEMP_854)
    );
    wire [2:0] _T_1239;
    wire [2:0] _WTEMP_855;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_5985 (
        .y(_WTEMP_855),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(3)) u_mux_5986 (
        .y(_T_1239),
        .sel(_T_1223),
        .a(_T_1237),
        .b(_WTEMP_855)
    );
    wire [2:0] _T_1241;
    wire [2:0] _WTEMP_856;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_5987 (
        .y(_WTEMP_856),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(3)) u_mux_5988 (
        .y(_T_1241),
        .sel(_T_1221),
        .a(_T_1239),
        .b(_WTEMP_856)
    );
    wire [2:0] _T_1243;
    wire [2:0] _WTEMP_857;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_5989 (
        .y(_WTEMP_857),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(3)) u_mux_5990 (
        .y(_T_1243),
        .sel(_T_1219),
        .a(_T_1241),
        .b(_WTEMP_857)
    );
    wire [52:0] _T_1244;
    wire [52:0] _WTEMP_858;
    PAD_UNSIGNED #(.width(3), .n(53)) u_pad_5991 (
        .y(_WTEMP_858),
        .in(_T_1243)
    );
    MUX_UNSIGNED #(.width(53)) u_mux_5992 (
        .y(_T_1244),
        .sel(_T_1087),
        .a(_T_1218),
        .b(_WTEMP_858)
    );
    wire [52:0] _T_1246;
    wire [52:0] _WTEMP_859;
    PAD_UNSIGNED #(.width(1), .n(53)) u_pad_5993 (
        .y(_WTEMP_859),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(53)) u_mux_5994 (
        .y(_T_1246),
        .sel(_T_1085),
        .a(_T_1244),
        .b(_WTEMP_859)
    );
    wire [52:0] roundMask_E;
    wire [52:0] _WTEMP_860;
    PAD_UNSIGNED #(.width(1), .n(53)) u_pad_5995 (
        .y(_WTEMP_860),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(53)) u_mux_5996 (
        .y(roundMask_E),
        .sel(_T_1083),
        .a(_T_1246),
        .b(_WTEMP_860)
    );
    wire [53:0] _T_1249;
    CAT #(.width_a(1), .width_b(53)) cat_5997 (
        .y(_T_1249),
        .a(1'h0),
        .b(roundMask_E)
    );
    wire [53:0] _T_1250;
    BITWISENOT #(.width(54)) bitwisenot_5998 (
        .y(_T_1250),
        .in(_T_1249)
    );
    wire [53:0] _T_1252;
    CAT #(.width_a(53), .width_b(1)) cat_5999 (
        .y(_T_1252),
        .a(roundMask_E),
        .b(1'h1)
    );
    wire [53:0] incrPosMask_E;
    BITWISEAND #(.width(54)) bitwiseand_6000 (
        .y(incrPosMask_E),
        .a(_T_1250),
        .b(_T_1252)
    );
    wire [52:0] _T_1253;
    SHR_UNSIGNED #(.width(54), .n(1)) u_shr_6001 (
        .y(_T_1253),
        .in(incrPosMask_E)
    );
    wire [52:0] _T_1254;
    BITWISEAND #(.width(53)) bitwiseand_6002 (
        .y(_T_1254),
        .a(_sigT_E__q),
        .b(_T_1253)
    );
    wire hiRoundPosBitT_E;
    wire [52:0] _WTEMP_861;
    PAD_UNSIGNED #(.width(1), .n(53)) u_pad_6003 (
        .y(_WTEMP_861),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(53)) u_neq_6004 (
        .y(hiRoundPosBitT_E),
        .a(_T_1254),
        .b(_WTEMP_861)
    );
    wire [51:0] _T_1256;
    SHR_UNSIGNED #(.width(53), .n(1)) u_shr_6005 (
        .y(_T_1256),
        .in(roundMask_E)
    );
    wire [52:0] _T_1257;
    wire [52:0] _WTEMP_862;
    PAD_UNSIGNED #(.width(52), .n(53)) u_pad_6006 (
        .y(_WTEMP_862),
        .in(_T_1256)
    );
    BITWISEAND #(.width(53)) bitwiseand_6007 (
        .y(_T_1257),
        .a(_sigT_E__q),
        .b(_WTEMP_862)
    );
    wire all0sHiRoundExtraT_E;
    wire [52:0] _WTEMP_863;
    PAD_UNSIGNED #(.width(1), .n(53)) u_pad_6008 (
        .y(_WTEMP_863),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(53)) u_eq_6009 (
        .y(all0sHiRoundExtraT_E),
        .a(_T_1257),
        .b(_WTEMP_863)
    );
    wire [52:0] _T_1259;
    BITWISENOT #(.width(53)) bitwisenot_6010 (
        .y(_T_1259),
        .in(_sigT_E__q)
    );
    wire [51:0] _T_1260;
    SHR_UNSIGNED #(.width(53), .n(1)) u_shr_6011 (
        .y(_T_1260),
        .in(roundMask_E)
    );
    wire [52:0] _T_1261;
    wire [52:0] _WTEMP_864;
    PAD_UNSIGNED #(.width(52), .n(53)) u_pad_6012 (
        .y(_WTEMP_864),
        .in(_T_1260)
    );
    BITWISEAND #(.width(53)) bitwiseand_6013 (
        .y(_T_1261),
        .a(_T_1259),
        .b(_WTEMP_864)
    );
    wire all1sHiRoundExtraT_E;
    wire [52:0] _WTEMP_865;
    PAD_UNSIGNED #(.width(1), .n(53)) u_pad_6014 (
        .y(_WTEMP_865),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(53)) u_eq_6015 (
        .y(all1sHiRoundExtraT_E),
        .a(_T_1261),
        .b(_WTEMP_865)
    );
    wire _T_1263;
    BITS #(.width(53), .high(0), .low(0)) bits_6016 (
        .y(_T_1263),
        .in(roundMask_E)
    );
    wire _T_1265;
    EQ_UNSIGNED #(.width(1)) u_eq_6017 (
        .y(_T_1265),
        .a(_T_1263),
        .b(1'h0)
    );
    wire _T_1266;
    BITWISEOR #(.width(1)) bitwiseor_6018 (
        .y(_T_1266),
        .a(_T_1265),
        .b(hiRoundPosBitT_E)
    );
    wire all1sHiRoundT_E;
    BITWISEAND #(.width(1)) bitwiseand_6019 (
        .y(all1sHiRoundT_E),
        .a(_T_1266),
        .b(all1sHiRoundExtraT_E)
    );
    wire [54:0] _T_1268;
    wire [53:0] _WTEMP_866;
    PAD_UNSIGNED #(.width(53), .n(54)) u_pad_6020 (
        .y(_WTEMP_866),
        .in(_sigT_E__q)
    );
    ADD_UNSIGNED #(.width(54)) u_add_6021 (
        .y(_T_1268),
        .a(54'h0),
        .b(_WTEMP_866)
    );
    wire [53:0] _T_1269;
    TAIL #(.width(55), .n(1)) tail_6022 (
        .y(_T_1269),
        .in(_T_1268)
    );
    wire [54:0] _T_1270;
    wire [53:0] _WTEMP_867;
    PAD_UNSIGNED #(.width(1), .n(54)) u_pad_6023 (
        .y(_WTEMP_867),
        .in(roundMagUp_PC)
    );
    ADD_UNSIGNED #(.width(54)) u_add_6024 (
        .y(_T_1270),
        .a(_T_1269),
        .b(_WTEMP_867)
    );
    wire [53:0] sigAdjT_E;
    TAIL #(.width(55), .n(1)) tail_6025 (
        .y(sigAdjT_E),
        .in(_T_1270)
    );
    wire [52:0] _T_1272;
    BITWISENOT #(.width(53)) bitwisenot_6026 (
        .y(_T_1272),
        .in(roundMask_E)
    );
    wire [53:0] _T_1273;
    CAT #(.width_a(1), .width_b(53)) cat_6027 (
        .y(_T_1273),
        .a(1'h1),
        .b(_T_1272)
    );
    wire [53:0] sigY0_E;
    BITWISEAND #(.width(54)) bitwiseand_6028 (
        .y(sigY0_E),
        .a(sigAdjT_E),
        .b(_T_1273)
    );
    wire [53:0] _T_1275;
    CAT #(.width_a(1), .width_b(53)) cat_6029 (
        .y(_T_1275),
        .a(1'h0),
        .b(roundMask_E)
    );
    wire [53:0] _T_1276;
    BITWISEOR #(.width(54)) bitwiseor_6030 (
        .y(_T_1276),
        .a(sigAdjT_E),
        .b(_T_1275)
    );
    wire [54:0] _T_1278;
    wire [53:0] _WTEMP_868;
    PAD_UNSIGNED #(.width(1), .n(54)) u_pad_6031 (
        .y(_WTEMP_868),
        .in(1'h1)
    );
    ADD_UNSIGNED #(.width(54)) u_add_6032 (
        .y(_T_1278),
        .a(_T_1276),
        .b(_WTEMP_868)
    );
    wire [53:0] sigY1_E;
    TAIL #(.width(55), .n(1)) tail_6033 (
        .y(sigY1_E),
        .in(_T_1278)
    );
    wire _T_1280;
    EQ_UNSIGNED #(.width(1)) u_eq_6034 (
        .y(_T_1280),
        .a(_isNegRemT_E__q),
        .b(1'h0)
    );
    wire _T_1282;
    EQ_UNSIGNED #(.width(1)) u_eq_6035 (
        .y(_T_1282),
        .a(_isZeroRemT_E__q),
        .b(1'h0)
    );
    wire _T_1283;
    BITWISEAND #(.width(1)) bitwiseand_6036 (
        .y(_T_1283),
        .a(_T_1280),
        .b(_T_1282)
    );
    wire trueLtX_E1;
    MUX_UNSIGNED #(.width(1)) u_mux_6037 (
        .y(trueLtX_E1),
        .sel(_sqrtOp_PC__q),
        .a(_T_1283),
        .b(_isNegRemT_E__q)
    );
    wire _T_1284;
    BITS #(.width(53), .high(0), .low(0)) bits_6038 (
        .y(_T_1284),
        .in(roundMask_E)
    );
    wire _T_1286;
    EQ_UNSIGNED #(.width(1)) u_eq_6039 (
        .y(_T_1286),
        .a(trueLtX_E1),
        .b(1'h0)
    );
    wire _T_1287;
    BITWISEAND #(.width(1)) bitwiseand_6040 (
        .y(_T_1287),
        .a(_T_1284),
        .b(_T_1286)
    );
    wire _T_1288;
    BITWISEAND #(.width(1)) bitwiseand_6041 (
        .y(_T_1288),
        .a(_T_1287),
        .b(all1sHiRoundExtraT_E)
    );
    wire _T_1289;
    BITWISEAND #(.width(1)) bitwiseand_6042 (
        .y(_T_1289),
        .a(_T_1288),
        .b(_extraT_E__q)
    );
    wire hiRoundPosBit_E1;
    BITWISEXOR #(.width(1)) bitwisexor_6043 (
        .y(hiRoundPosBit_E1),
        .a(hiRoundPosBitT_E),
        .b(_T_1289)
    );
    wire _T_1291;
    EQ_UNSIGNED #(.width(1)) u_eq_6044 (
        .y(_T_1291),
        .a(_isZeroRemT_E__q),
        .b(1'h0)
    );
    wire _T_1293;
    EQ_UNSIGNED #(.width(1)) u_eq_6045 (
        .y(_T_1293),
        .a(_extraT_E__q),
        .b(1'h0)
    );
    wire _T_1294;
    BITWISEOR #(.width(1)) bitwiseor_6046 (
        .y(_T_1294),
        .a(_T_1291),
        .b(_T_1293)
    );
    wire _T_1296;
    EQ_UNSIGNED #(.width(1)) u_eq_6047 (
        .y(_T_1296),
        .a(all1sHiRoundExtraT_E),
        .b(1'h0)
    );
    wire anyRoundExtra_E1;
    BITWISEOR #(.width(1)) bitwiseor_6048 (
        .y(anyRoundExtra_E1),
        .a(_T_1294),
        .b(_T_1296)
    );
    wire _T_1297;
    BITWISEAND #(.width(1)) bitwiseand_6049 (
        .y(_T_1297),
        .a(roundingMode_near_even_PC),
        .b(hiRoundPosBit_E1)
    );
    wire _T_1299;
    EQ_UNSIGNED #(.width(1)) u_eq_6050 (
        .y(_T_1299),
        .a(anyRoundExtra_E1),
        .b(1'h0)
    );
    wire _T_1300;
    BITWISEAND #(.width(1)) bitwiseand_6051 (
        .y(_T_1300),
        .a(_T_1297),
        .b(_T_1299)
    );
    wire [53:0] roundEvenMask_E1;
    wire [53:0] _WTEMP_869;
    PAD_UNSIGNED #(.width(1), .n(54)) u_pad_6052 (
        .y(_WTEMP_869),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(54)) u_mux_6053 (
        .y(roundEvenMask_E1),
        .sel(_T_1300),
        .a(incrPosMask_E),
        .b(_WTEMP_869)
    );
    wire _T_1302;
    BITWISEAND #(.width(1)) bitwiseand_6054 (
        .y(_T_1302),
        .a(roundMagDown_PC),
        .b(_extraT_E__q)
    );
    wire _T_1304;
    EQ_UNSIGNED #(.width(1)) u_eq_6055 (
        .y(_T_1304),
        .a(trueLtX_E1),
        .b(1'h0)
    );
    wire _T_1305;
    BITWISEAND #(.width(1)) bitwiseand_6056 (
        .y(_T_1305),
        .a(_T_1302),
        .b(_T_1304)
    );
    wire _T_1306;
    BITWISEAND #(.width(1)) bitwiseand_6057 (
        .y(_T_1306),
        .a(_T_1305),
        .b(all1sHiRoundT_E)
    );
    wire _T_1308;
    EQ_UNSIGNED #(.width(1)) u_eq_6058 (
        .y(_T_1308),
        .a(trueLtX_E1),
        .b(1'h0)
    );
    wire _T_1309;
    BITWISEAND #(.width(1)) bitwiseand_6059 (
        .y(_T_1309),
        .a(_extraT_E__q),
        .b(_T_1308)
    );
    wire _T_1311;
    EQ_UNSIGNED #(.width(1)) u_eq_6060 (
        .y(_T_1311),
        .a(_isZeroRemT_E__q),
        .b(1'h0)
    );
    wire _T_1312;
    BITWISEAND #(.width(1)) bitwiseand_6061 (
        .y(_T_1312),
        .a(_T_1309),
        .b(_T_1311)
    );
    wire _T_1314;
    EQ_UNSIGNED #(.width(1)) u_eq_6062 (
        .y(_T_1314),
        .a(all1sHiRoundT_E),
        .b(1'h0)
    );
    wire _T_1315;
    BITWISEOR #(.width(1)) bitwiseor_6063 (
        .y(_T_1315),
        .a(_T_1312),
        .b(_T_1314)
    );
    wire _T_1316;
    BITWISEAND #(.width(1)) bitwiseand_6064 (
        .y(_T_1316),
        .a(roundMagUp_PC),
        .b(_T_1315)
    );
    wire _T_1317;
    BITWISEOR #(.width(1)) bitwiseor_6065 (
        .y(_T_1317),
        .a(_T_1306),
        .b(_T_1316)
    );
    wire _T_1319;
    EQ_UNSIGNED #(.width(1)) u_eq_6066 (
        .y(_T_1319),
        .a(trueLtX_E1),
        .b(1'h0)
    );
    wire _T_1320;
    BITWISEOR #(.width(1)) bitwiseor_6067 (
        .y(_T_1320),
        .a(_extraT_E__q),
        .b(_T_1319)
    );
    wire _T_1321;
    BITS #(.width(53), .high(0), .low(0)) bits_6068 (
        .y(_T_1321),
        .in(roundMask_E)
    );
    wire _T_1323;
    EQ_UNSIGNED #(.width(1)) u_eq_6069 (
        .y(_T_1323),
        .a(_T_1321),
        .b(1'h0)
    );
    wire _T_1324;
    BITWISEAND #(.width(1)) bitwiseand_6070 (
        .y(_T_1324),
        .a(_T_1320),
        .b(_T_1323)
    );
    wire _T_1325;
    BITWISEOR #(.width(1)) bitwiseor_6071 (
        .y(_T_1325),
        .a(hiRoundPosBitT_E),
        .b(_T_1324)
    );
    wire _T_1327;
    EQ_UNSIGNED #(.width(1)) u_eq_6072 (
        .y(_T_1327),
        .a(trueLtX_E1),
        .b(1'h0)
    );
    wire _T_1328;
    BITWISEAND #(.width(1)) bitwiseand_6073 (
        .y(_T_1328),
        .a(_extraT_E__q),
        .b(_T_1327)
    );
    wire _T_1329;
    BITWISEAND #(.width(1)) bitwiseand_6074 (
        .y(_T_1329),
        .a(_T_1328),
        .b(all1sHiRoundExtraT_E)
    );
    wire _T_1330;
    BITWISEOR #(.width(1)) bitwiseor_6075 (
        .y(_T_1330),
        .a(_T_1325),
        .b(_T_1329)
    );
    wire _T_1331;
    BITWISEAND #(.width(1)) bitwiseand_6076 (
        .y(_T_1331),
        .a(roundingMode_near_even_PC),
        .b(_T_1330)
    );
    wire _T_1332;
    BITWISEOR #(.width(1)) bitwiseor_6077 (
        .y(_T_1332),
        .a(_T_1317),
        .b(_T_1331)
    );
    wire [53:0] _T_1333;
    MUX_UNSIGNED #(.width(54)) u_mux_6078 (
        .y(_T_1333),
        .sel(_T_1332),
        .a(sigY1_E),
        .b(sigY0_E)
    );
    wire [53:0] _T_1334;
    BITWISENOT #(.width(54)) bitwisenot_6079 (
        .y(_T_1334),
        .in(roundEvenMask_E1)
    );
    wire [53:0] sigY_E1;
    BITWISEAND #(.width(54)) bitwiseand_6080 (
        .y(sigY_E1),
        .a(_T_1333),
        .b(_T_1334)
    );
    wire [51:0] fractY_E1;
    BITS #(.width(54), .high(51), .low(0)) bits_6081 (
        .y(fractY_E1),
        .in(sigY_E1)
    );
    wire inexactY_E1;
    BITWISEOR #(.width(1)) bitwiseor_6082 (
        .y(inexactY_E1),
        .a(hiRoundPosBit_E1),
        .b(anyRoundExtra_E1)
    );
    wire _T_1335;
    BITS #(.width(54), .high(53), .low(53)) bits_6083 (
        .y(_T_1335),
        .in(sigY_E1)
    );
    wire _T_1337;
    EQ_UNSIGNED #(.width(1)) u_eq_6084 (
        .y(_T_1337),
        .a(_T_1335),
        .b(1'h0)
    );
    wire [13:0] _T_1339;
    wire [13:0] _WTEMP_870;
    PAD_UNSIGNED #(.width(1), .n(14)) u_pad_6085 (
        .y(_WTEMP_870),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(14)) u_mux_6086 (
        .y(_T_1339),
        .sel(_T_1337),
        .a(sExpX_E),
        .b(_WTEMP_870)
    );
    wire _T_1340;
    BITS #(.width(54), .high(53), .low(53)) bits_6087 (
        .y(_T_1340),
        .in(sigY_E1)
    );
    wire _T_1342;
    EQ_UNSIGNED #(.width(1)) u_eq_6088 (
        .y(_T_1342),
        .a(_sqrtOp_PC__q),
        .b(1'h0)
    );
    wire _T_1343;
    BITWISEAND #(.width(1)) bitwiseand_6089 (
        .y(_T_1343),
        .a(_T_1340),
        .b(_T_1342)
    );
    wire _T_1344;
    BITWISEAND #(.width(1)) bitwiseand_6090 (
        .y(_T_1344),
        .a(_T_1343),
        .b(_E_E_div__q)
    );
    wire [13:0] _T_1346;
    wire [13:0] _WTEMP_871;
    PAD_UNSIGNED #(.width(1), .n(14)) u_pad_6091 (
        .y(_WTEMP_871),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(14)) u_mux_6092 (
        .y(_T_1346),
        .sel(_T_1344),
        .a(expP1_PC),
        .b(_WTEMP_871)
    );
    wire [13:0] _T_1347;
    BITWISEOR #(.width(14)) bitwiseor_6093 (
        .y(_T_1347),
        .a(_T_1339),
        .b(_T_1346)
    );
    wire _T_1348;
    BITS #(.width(54), .high(53), .low(53)) bits_6094 (
        .y(_T_1348),
        .in(sigY_E1)
    );
    wire _T_1350;
    EQ_UNSIGNED #(.width(1)) u_eq_6095 (
        .y(_T_1350),
        .a(_sqrtOp_PC__q),
        .b(1'h0)
    );
    wire _T_1351;
    BITWISEAND #(.width(1)) bitwiseand_6096 (
        .y(_T_1351),
        .a(_T_1348),
        .b(_T_1350)
    );
    wire _T_1353;
    EQ_UNSIGNED #(.width(1)) u_eq_6097 (
        .y(_T_1353),
        .a(_E_E_div__q),
        .b(1'h0)
    );
    wire _T_1354;
    BITWISEAND #(.width(1)) bitwiseand_6098 (
        .y(_T_1354),
        .a(_T_1351),
        .b(_T_1353)
    );
    wire [13:0] _T_1356;
    wire [13:0] _WTEMP_872;
    PAD_UNSIGNED #(.width(1), .n(14)) u_pad_6099 (
        .y(_WTEMP_872),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(14)) u_mux_6100 (
        .y(_T_1356),
        .sel(_T_1354),
        .a(expP2_PC),
        .b(_WTEMP_872)
    );
    wire [13:0] _T_1357;
    BITWISEOR #(.width(14)) bitwiseor_6101 (
        .y(_T_1357),
        .a(_T_1347),
        .b(_T_1356)
    );
    wire _T_1358;
    BITS #(.width(54), .high(53), .low(53)) bits_6102 (
        .y(_T_1358),
        .in(sigY_E1)
    );
    wire _T_1359;
    BITWISEAND #(.width(1)) bitwiseand_6103 (
        .y(_T_1359),
        .a(_T_1358),
        .b(_sqrtOp_PC__q)
    );
    wire [12:0] _T_1360;
    SHR_UNSIGNED #(.width(14), .n(1)) u_shr_6104 (
        .y(_T_1360),
        .in(expP2_PC)
    );
    wire [13:0] _T_1362;
    wire [12:0] _WTEMP_873;
    PAD_UNSIGNED #(.width(12), .n(13)) u_pad_6105 (
        .y(_WTEMP_873),
        .in(12'h400)
    );
    ADD_UNSIGNED #(.width(13)) u_add_6106 (
        .y(_T_1362),
        .a(_T_1360),
        .b(_WTEMP_873)
    );
    wire [12:0] _T_1363;
    TAIL #(.width(14), .n(1)) tail_6107 (
        .y(_T_1363),
        .in(_T_1362)
    );
    wire [12:0] _T_1365;
    wire [12:0] _WTEMP_874;
    PAD_UNSIGNED #(.width(1), .n(13)) u_pad_6108 (
        .y(_WTEMP_874),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(13)) u_mux_6109 (
        .y(_T_1365),
        .sel(_T_1359),
        .a(_T_1363),
        .b(_WTEMP_874)
    );
    wire [13:0] sExpY_E1;
    wire [13:0] _WTEMP_875;
    PAD_UNSIGNED #(.width(13), .n(14)) u_pad_6110 (
        .y(_WTEMP_875),
        .in(_T_1365)
    );
    BITWISEOR #(.width(14)) bitwiseor_6111 (
        .y(sExpY_E1),
        .a(_T_1357),
        .b(_WTEMP_875)
    );
    wire [11:0] expY_E1;
    BITS #(.width(14), .high(11), .low(0)) bits_6112 (
        .y(expY_E1),
        .in(sExpY_E1)
    );
    wire _T_1366;
    BITS #(.width(14), .high(13), .low(13)) bits_6113 (
        .y(_T_1366),
        .in(sExpY_E1)
    );
    wire _T_1368;
    EQ_UNSIGNED #(.width(1)) u_eq_6114 (
        .y(_T_1368),
        .a(_T_1366),
        .b(1'h0)
    );
    wire [2:0] _T_1370;
    BITS #(.width(14), .high(12), .low(10)) bits_6115 (
        .y(_T_1370),
        .in(sExpY_E1)
    );
    wire _T_1371;
    LEQ_UNSIGNED #(.width(3)) u_leq_6116 (
        .y(_T_1371),
        .a(3'h3),
        .b(_T_1370)
    );
    wire overflowY_E1;
    BITWISEAND #(.width(1)) bitwiseand_6117 (
        .y(overflowY_E1),
        .a(_T_1368),
        .b(_T_1371)
    );
    wire _T_1372;
    BITS #(.width(14), .high(13), .low(13)) bits_6118 (
        .y(_T_1372),
        .in(sExpY_E1)
    );
    wire [12:0] _T_1373;
    BITS #(.width(14), .high(12), .low(0)) bits_6119 (
        .y(_T_1373),
        .in(sExpY_E1)
    );
    wire _T_1375;
    LT_UNSIGNED #(.width(13)) u_lt_6120 (
        .y(_T_1375),
        .a(_T_1373),
        .b(13'h3CE)
    );
    wire totalUnderflowY_E1;
    BITWISEOR #(.width(1)) bitwiseor_6121 (
        .y(totalUnderflowY_E1),
        .a(_T_1372),
        .b(_T_1375)
    );
    wire _T_1377;
    LEQ_UNSIGNED #(.width(13)) u_leq_6122 (
        .y(_T_1377),
        .a(posExpX_E),
        .b(13'h401)
    );
    wire _T_1378;
    BITWISEAND #(.width(1)) bitwiseand_6123 (
        .y(_T_1378),
        .a(_T_1377),
        .b(inexactY_E1)
    );
    wire underflowY_E1;
    BITWISEOR #(.width(1)) bitwiseor_6124 (
        .y(underflowY_E1),
        .a(totalUnderflowY_E1),
        .b(_T_1378)
    );
    wire _T_1380;
    EQ_UNSIGNED #(.width(1)) u_eq_6125 (
        .y(_T_1380),
        .a(isNaNB_PC),
        .b(1'h0)
    );
    wire _T_1382;
    EQ_UNSIGNED #(.width(1)) u_eq_6126 (
        .y(_T_1382),
        .a(isZeroB_PC),
        .b(1'h0)
    );
    wire _T_1383;
    BITWISEAND #(.width(1)) bitwiseand_6127 (
        .y(_T_1383),
        .a(_T_1380),
        .b(_T_1382)
    );
    wire _T_1384;
    BITWISEAND #(.width(1)) bitwiseand_6128 (
        .y(_T_1384),
        .a(_T_1383),
        .b(_sign_PC__q)
    );
    wire _T_1385;
    BITWISEAND #(.width(1)) bitwiseand_6129 (
        .y(_T_1385),
        .a(isZeroA_PC),
        .b(isZeroB_PC)
    );
    wire _T_1386;
    BITWISEAND #(.width(1)) bitwiseand_6130 (
        .y(_T_1386),
        .a(isInfA_PC),
        .b(isInfB_PC)
    );
    wire _T_1387;
    BITWISEOR #(.width(1)) bitwiseor_6131 (
        .y(_T_1387),
        .a(_T_1385),
        .b(_T_1386)
    );
    wire notSigNaN_invalid_PC;
    MUX_UNSIGNED #(.width(1)) u_mux_6132 (
        .y(notSigNaN_invalid_PC),
        .sel(_sqrtOp_PC__q),
        .a(_T_1384),
        .b(_T_1387)
    );
    wire _T_1389;
    EQ_UNSIGNED #(.width(1)) u_eq_6133 (
        .y(_T_1389),
        .a(_sqrtOp_PC__q),
        .b(1'h0)
    );
    wire _T_1390;
    BITWISEAND #(.width(1)) bitwiseand_6134 (
        .y(_T_1390),
        .a(_T_1389),
        .b(isSigNaNA_PC)
    );
    wire _T_1391;
    BITWISEOR #(.width(1)) bitwiseor_6135 (
        .y(_T_1391),
        .a(_T_1390),
        .b(isSigNaNB_PC)
    );
    wire invalid_PC;
    BITWISEOR #(.width(1)) bitwiseor_6136 (
        .y(invalid_PC),
        .a(_T_1391),
        .b(notSigNaN_invalid_PC)
    );
    wire _T_1393;
    EQ_UNSIGNED #(.width(1)) u_eq_6137 (
        .y(_T_1393),
        .a(_sqrtOp_PC__q),
        .b(1'h0)
    );
    wire _T_1395;
    EQ_UNSIGNED #(.width(1)) u_eq_6138 (
        .y(_T_1395),
        .a(isSpecialA_PC),
        .b(1'h0)
    );
    wire _T_1396;
    BITWISEAND #(.width(1)) bitwiseand_6139 (
        .y(_T_1396),
        .a(_T_1393),
        .b(_T_1395)
    );
    wire _T_1398;
    EQ_UNSIGNED #(.width(1)) u_eq_6140 (
        .y(_T_1398),
        .a(isZeroA_PC),
        .b(1'h0)
    );
    wire _T_1399;
    BITWISEAND #(.width(1)) bitwiseand_6141 (
        .y(_T_1399),
        .a(_T_1396),
        .b(_T_1398)
    );
    wire infinity_PC;
    BITWISEAND #(.width(1)) bitwiseand_6142 (
        .y(infinity_PC),
        .a(_T_1399),
        .b(isZeroB_PC)
    );
    wire overflow_E1;
    BITWISEAND #(.width(1)) bitwiseand_6143 (
        .y(overflow_E1),
        .a(normalCase_PC),
        .b(overflowY_E1)
    );
    wire underflow_E1;
    BITWISEAND #(.width(1)) bitwiseand_6144 (
        .y(underflow_E1),
        .a(normalCase_PC),
        .b(underflowY_E1)
    );
    wire _T_1400;
    BITWISEOR #(.width(1)) bitwiseor_6145 (
        .y(_T_1400),
        .a(overflow_E1),
        .b(underflow_E1)
    );
    wire _T_1401;
    BITWISEAND #(.width(1)) bitwiseand_6146 (
        .y(_T_1401),
        .a(normalCase_PC),
        .b(inexactY_E1)
    );
    wire inexact_E1;
    BITWISEOR #(.width(1)) bitwiseor_6147 (
        .y(inexact_E1),
        .a(_T_1400),
        .b(_T_1401)
    );
    wire _T_1402;
    BITWISEOR #(.width(1)) bitwiseor_6148 (
        .y(_T_1402),
        .a(isZeroA_PC),
        .b(isInfB_PC)
    );
    wire _T_1404;
    EQ_UNSIGNED #(.width(1)) u_eq_6149 (
        .y(_T_1404),
        .a(roundMagUp_PC),
        .b(1'h0)
    );
    wire _T_1405;
    BITWISEAND #(.width(1)) bitwiseand_6150 (
        .y(_T_1405),
        .a(totalUnderflowY_E1),
        .b(_T_1404)
    );
    wire _T_1406;
    BITWISEOR #(.width(1)) bitwiseor_6151 (
        .y(_T_1406),
        .a(_T_1402),
        .b(_T_1405)
    );
    wire notSpecial_isZeroOut_E1;
    MUX_UNSIGNED #(.width(1)) u_mux_6152 (
        .y(notSpecial_isZeroOut_E1),
        .sel(_sqrtOp_PC__q),
        .a(isZeroB_PC),
        .b(_T_1406)
    );
    wire _T_1407;
    BITWISEAND #(.width(1)) bitwiseand_6153 (
        .y(_T_1407),
        .a(normalCase_PC),
        .b(totalUnderflowY_E1)
    );
    wire pegMinFiniteMagOut_E1;
    BITWISEAND #(.width(1)) bitwiseand_6154 (
        .y(pegMinFiniteMagOut_E1),
        .a(_T_1407),
        .b(roundMagUp_PC)
    );
    wire _T_1409;
    EQ_UNSIGNED #(.width(1)) u_eq_6155 (
        .y(_T_1409),
        .a(overflowY_roundMagUp_PC),
        .b(1'h0)
    );
    wire pegMaxFiniteMagOut_E1;
    BITWISEAND #(.width(1)) bitwiseand_6156 (
        .y(pegMaxFiniteMagOut_E1),
        .a(overflow_E1),
        .b(_T_1409)
    );
    wire _T_1410;
    BITWISEOR #(.width(1)) bitwiseor_6157 (
        .y(_T_1410),
        .a(isInfA_PC),
        .b(isZeroB_PC)
    );
    wire _T_1411;
    BITWISEAND #(.width(1)) bitwiseand_6158 (
        .y(_T_1411),
        .a(overflow_E1),
        .b(overflowY_roundMagUp_PC)
    );
    wire _T_1412;
    BITWISEOR #(.width(1)) bitwiseor_6159 (
        .y(_T_1412),
        .a(_T_1410),
        .b(_T_1411)
    );
    wire notNaN_isInfOut_E1;
    MUX_UNSIGNED #(.width(1)) u_mux_6160 (
        .y(notNaN_isInfOut_E1),
        .sel(_sqrtOp_PC__q),
        .a(isInfB_PC),
        .b(_T_1412)
    );
    wire _T_1414;
    EQ_UNSIGNED #(.width(1)) u_eq_6161 (
        .y(_T_1414),
        .a(_sqrtOp_PC__q),
        .b(1'h0)
    );
    wire _T_1415;
    BITWISEAND #(.width(1)) bitwiseand_6162 (
        .y(_T_1415),
        .a(_T_1414),
        .b(isNaNA_PC)
    );
    wire _T_1416;
    BITWISEOR #(.width(1)) bitwiseor_6163 (
        .y(_T_1416),
        .a(_T_1415),
        .b(isNaNB_PC)
    );
    wire isNaNOut_PC;
    BITWISEOR #(.width(1)) bitwiseor_6164 (
        .y(isNaNOut_PC),
        .a(_T_1416),
        .b(notSigNaN_invalid_PC)
    );
    wire _T_1418;
    EQ_UNSIGNED #(.width(1)) u_eq_6165 (
        .y(_T_1418),
        .a(isNaNOut_PC),
        .b(1'h0)
    );
    wire _T_1419;
    BITWISEAND #(.width(1)) bitwiseand_6166 (
        .y(_T_1419),
        .a(isZeroB_PC),
        .b(_sign_PC__q)
    );
    wire _T_1420;
    MUX_UNSIGNED #(.width(1)) u_mux_6167 (
        .y(_T_1420),
        .sel(_sqrtOp_PC__q),
        .a(_T_1419),
        .b(_sign_PC__q)
    );
    wire signOut_PC;
    BITWISEAND #(.width(1)) bitwiseand_6168 (
        .y(signOut_PC),
        .a(_T_1418),
        .b(_T_1420)
    );
    wire [11:0] _T_1422;
    assign _T_1422 = 12'hE00;
    wire [11:0] _T_1424;
    wire [11:0] _WTEMP_876;
    PAD_UNSIGNED #(.width(1), .n(12)) u_pad_6169 (
        .y(_WTEMP_876),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(12)) u_mux_6170 (
        .y(_T_1424),
        .sel(notSpecial_isZeroOut_E1),
        .a(_T_1422),
        .b(_WTEMP_876)
    );
    wire [11:0] _T_1425;
    BITWISENOT #(.width(12)) bitwisenot_6171 (
        .y(_T_1425),
        .in(_T_1424)
    );
    wire [11:0] _T_1426;
    BITWISEAND #(.width(12)) bitwiseand_6172 (
        .y(_T_1426),
        .a(expY_E1),
        .b(_T_1425)
    );
    wire [11:0] _T_1428;
    assign _T_1428 = 12'hC31;
    wire [11:0] _T_1430;
    wire [11:0] _WTEMP_877;
    PAD_UNSIGNED #(.width(1), .n(12)) u_pad_6173 (
        .y(_WTEMP_877),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(12)) u_mux_6174 (
        .y(_T_1430),
        .sel(pegMinFiniteMagOut_E1),
        .a(_T_1428),
        .b(_WTEMP_877)
    );
    wire [11:0] _T_1431;
    BITWISENOT #(.width(12)) bitwisenot_6175 (
        .y(_T_1431),
        .in(_T_1430)
    );
    wire [11:0] _T_1432;
    BITWISEAND #(.width(12)) bitwiseand_6176 (
        .y(_T_1432),
        .a(_T_1426),
        .b(_T_1431)
    );
    wire [11:0] _T_1434;
    assign _T_1434 = 12'h400;
    wire [11:0] _T_1436;
    wire [11:0] _WTEMP_878;
    PAD_UNSIGNED #(.width(1), .n(12)) u_pad_6177 (
        .y(_WTEMP_878),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(12)) u_mux_6178 (
        .y(_T_1436),
        .sel(pegMaxFiniteMagOut_E1),
        .a(_T_1434),
        .b(_WTEMP_878)
    );
    wire [11:0] _T_1437;
    BITWISENOT #(.width(12)) bitwisenot_6179 (
        .y(_T_1437),
        .in(_T_1436)
    );
    wire [11:0] _T_1438;
    BITWISEAND #(.width(12)) bitwiseand_6180 (
        .y(_T_1438),
        .a(_T_1432),
        .b(_T_1437)
    );
    wire [11:0] _T_1440;
    assign _T_1440 = 12'h200;
    wire [11:0] _T_1442;
    wire [11:0] _WTEMP_879;
    PAD_UNSIGNED #(.width(1), .n(12)) u_pad_6181 (
        .y(_WTEMP_879),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(12)) u_mux_6182 (
        .y(_T_1442),
        .sel(notNaN_isInfOut_E1),
        .a(_T_1440),
        .b(_WTEMP_879)
    );
    wire [11:0] _T_1443;
    BITWISENOT #(.width(12)) bitwisenot_6183 (
        .y(_T_1443),
        .in(_T_1442)
    );
    wire [11:0] _T_1444;
    BITWISEAND #(.width(12)) bitwiseand_6184 (
        .y(_T_1444),
        .a(_T_1438),
        .b(_T_1443)
    );
    wire [11:0] _T_1447;
    wire [11:0] _WTEMP_880;
    PAD_UNSIGNED #(.width(1), .n(12)) u_pad_6185 (
        .y(_WTEMP_880),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(12)) u_mux_6186 (
        .y(_T_1447),
        .sel(pegMinFiniteMagOut_E1),
        .a(12'h3CE),
        .b(_WTEMP_880)
    );
    wire [11:0] _T_1448;
    BITWISEOR #(.width(12)) bitwiseor_6187 (
        .y(_T_1448),
        .a(_T_1444),
        .b(_T_1447)
    );
    wire [11:0] _T_1451;
    wire [11:0] _WTEMP_881;
    PAD_UNSIGNED #(.width(1), .n(12)) u_pad_6188 (
        .y(_WTEMP_881),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(12)) u_mux_6189 (
        .y(_T_1451),
        .sel(pegMaxFiniteMagOut_E1),
        .a(12'hBFF),
        .b(_WTEMP_881)
    );
    wire [11:0] _T_1452;
    BITWISEOR #(.width(12)) bitwiseor_6190 (
        .y(_T_1452),
        .a(_T_1448),
        .b(_T_1451)
    );
    wire [11:0] _T_1455;
    wire [11:0] _WTEMP_882;
    PAD_UNSIGNED #(.width(1), .n(12)) u_pad_6191 (
        .y(_WTEMP_882),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(12)) u_mux_6192 (
        .y(_T_1455),
        .sel(notNaN_isInfOut_E1),
        .a(12'hC00),
        .b(_WTEMP_882)
    );
    wire [11:0] _T_1456;
    BITWISEOR #(.width(12)) bitwiseor_6193 (
        .y(_T_1456),
        .a(_T_1452),
        .b(_T_1455)
    );
    wire [11:0] _T_1459;
    wire [11:0] _WTEMP_883;
    PAD_UNSIGNED #(.width(1), .n(12)) u_pad_6194 (
        .y(_WTEMP_883),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(12)) u_mux_6195 (
        .y(_T_1459),
        .sel(isNaNOut_PC),
        .a(12'hE00),
        .b(_WTEMP_883)
    );
    wire [11:0] expOut_E1;
    BITWISEOR #(.width(12)) bitwiseor_6196 (
        .y(expOut_E1),
        .a(_T_1456),
        .b(_T_1459)
    );
    wire _T_1460;
    BITWISEOR #(.width(1)) bitwiseor_6197 (
        .y(_T_1460),
        .a(notSpecial_isZeroOut_E1),
        .b(totalUnderflowY_E1)
    );
    wire _T_1461;
    BITWISEOR #(.width(1)) bitwiseor_6198 (
        .y(_T_1461),
        .a(_T_1460),
        .b(isNaNOut_PC)
    );
    wire [51:0] _T_1463;
    assign _T_1463 = 52'h8000000000000;
    wire [51:0] _T_1465;
    wire [51:0] _WTEMP_884;
    PAD_UNSIGNED #(.width(1), .n(52)) u_pad_6199 (
        .y(_WTEMP_884),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(52)) u_mux_6200 (
        .y(_T_1465),
        .sel(isNaNOut_PC),
        .a(_T_1463),
        .b(_WTEMP_884)
    );
    wire [51:0] _T_1466;
    MUX_UNSIGNED #(.width(52)) u_mux_6201 (
        .y(_T_1466),
        .sel(_T_1461),
        .a(_T_1465),
        .b(fractY_E1)
    );
    wire _T_1467;
    BITS #(.width(1), .high(0), .low(0)) bits_6202 (
        .y(_T_1467),
        .in(pegMaxFiniteMagOut_E1)
    );
    wire [51:0] _T_1470;
    MUX_UNSIGNED #(.width(52)) u_mux_6203 (
        .y(_T_1470),
        .sel(_T_1467),
        .a(52'hFFFFFFFFFFFFF),
        .b(52'h0)
    );
    wire [51:0] fractOut_E1;
    BITWISEOR #(.width(52)) bitwiseor_6204 (
        .y(fractOut_E1),
        .a(_T_1466),
        .b(_T_1470)
    );
    wire [12:0] _T_1471;
    CAT #(.width_a(1), .width_b(12)) cat_6205 (
        .y(_T_1471),
        .a(signOut_PC),
        .b(expOut_E1)
    );
    wire [64:0] _T_1472;
    CAT #(.width_a(13), .width_b(52)) cat_6206 (
        .y(_T_1472),
        .a(_T_1471),
        .b(fractOut_E1)
    );
    wire [1:0] _T_1473;
    CAT #(.width_a(1), .width_b(1)) cat_6207 (
        .y(_T_1473),
        .a(underflow_E1),
        .b(inexact_E1)
    );
    wire [1:0] _T_1474;
    CAT #(.width_a(1), .width_b(1)) cat_6208 (
        .y(_T_1474),
        .a(invalid_PC),
        .b(infinity_PC)
    );
    wire [2:0] _T_1475;
    CAT #(.width_a(2), .width_b(1)) cat_6209 (
        .y(_T_1475),
        .a(_T_1474),
        .b(overflow_E1)
    );
    wire [4:0] _T_1476;
    CAT #(.width_a(3), .width_b(2)) cat_6210 (
        .y(_T_1476),
        .a(_T_1475),
        .b(_T_1473)
    );
    MUX_UNSIGNED #(.width(17)) u_mux_6211 (
        .y(_ER1_B_sqrt__d),
        .sel(cyc_A1_sqrt),
        .a(ER1_A1_sqrt),
        .b(_ER1_B_sqrt__q)
    );
    MUX_UNSIGNED #(.width(32)) u_mux_6212 (
        .y(_ESqrR1_B_sqrt__d),
        .sel(cyc_B8_sqrt),
        .a(ESqrR1_B8_sqrt),
        .b(_ESqrR1_B_sqrt__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6213 (
        .y(_E_E_div__d),
        .sel(cyc_C1),
        .a(E_C1_div),
        .b(_E_E_div__q)
    );
    assign cyc_B1 = _T_454;
    assign cyc_B10_sqrt = _T_436;
    assign cyc_B1_div = _T_475;
    assign cyc_B1_sqrt = _T_484;
    assign cyc_B2 = _T_452;
    assign cyc_B2_div = _T_472;
    assign cyc_B2_sqrt = _T_483;
    assign cyc_B3 = _T_450;
    assign cyc_B3_div = _T_469;
    assign cyc_B3_sqrt = _T_482;
    assign cyc_B4 = _T_448;
    assign cyc_B4_div = _T_466;
    assign cyc_B4_sqrt = _T_481;
    assign cyc_B5 = _T_446;
    assign cyc_B5_div = _T_462;
    assign cyc_B5_sqrt = _T_479;
    assign cyc_B6 = _T_444;
    assign cyc_B6_div = _T_458;
    assign cyc_B6_sqrt = _T_477;
    assign cyc_B7_sqrt = _T_442;
    assign cyc_B8_sqrt = _T_440;
    assign cyc_B9_sqrt = _T_438;
    assign cyc_C1 = _T_506;
    assign cyc_C2 = _T_504;
    assign cyc_C3 = _T_502;
    assign cyc_C4 = _T_500;
    assign cyc_C5 = _T_498;
    assign cyc_E1 = _T_533;
    assign cyc_E2 = _T_531;
    assign cyc_E3 = _T_529;
    assign cyc_E4 = _T_527;
    MUX_UNSIGNED #(.width(3)) u_mux_6214 (
        .y(_WTEMP_694),
        .sel(_T_395),
        .a(_T_411),
        .b(_cycleNum_A__q)
    );
    MUX_UNSIGNED #(.width(4)) u_mux_6215 (
        .y(_WTEMP_695),
        .sel(_T_426),
        .a(_T_434),
        .b(_cycleNum_B__q)
    );
    MUX_UNSIGNED #(.width(3)) u_mux_6216 (
        .y(_WTEMP_696),
        .sel(_T_487),
        .a(_T_495),
        .b(_cycleNum_C__q)
    );
    MUX_UNSIGNED #(.width(3)) u_mux_6217 (
        .y(_WTEMP_697),
        .sel(_T_519),
        .a(_T_525),
        .b(_cycleNum_E__q)
    );
    MUX_UNSIGNED #(.width(14)) u_mux_6218 (
        .y(_exp_PA__d),
        .sel(entering_PA_normalCase),
        .a(_T_243),
        .b(_exp_PA__q)
    );
    MUX_UNSIGNED #(.width(14)) u_mux_6219 (
        .y(_exp_PB__d),
        .sel(entering_PB_normalCase),
        .a(_exp_PA__q),
        .b(_exp_PB__q)
    );
    MUX_UNSIGNED #(.width(14)) u_mux_6220 (
        .y(_exp_PC__d),
        .sel(entering_PC_normalCase),
        .a(_exp_PB__q),
        .b(_exp_PC__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6221 (
        .y(_extraT_E__d),
        .sel(cyc_C1),
        .a(_T_1049),
        .b(_extraT_E__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6222 (
        .y(_fractA_0_PB__d),
        .sel(entering_PB_normalCase),
        .a(_T_290),
        .b(_fractA_0_PB__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6223 (
        .y(_fractA_0_PC__d),
        .sel(entering_PC_normalCase),
        .a(_fractA_0_PB__q),
        .b(_fractA_0_PC__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6224 (
        .y(_fractA_51_PA__d),
        .sel(_T_231),
        .a(_T_232),
        .b(_fractA_51_PA__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6225 (
        .y(_fractA_51_PB__d),
        .sel(entering_PB),
        .a(_T_285),
        .b(_fractA_51_PB__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6226 (
        .y(_fractA_51_PC__d),
        .sel(entering_PC),
        .a(_T_326),
        .b(_fractA_51_PC__q)
    );
    MUX_UNSIGNED #(.width(51)) u_mux_6227 (
        .y(_fractA_other_PA__d),
        .sel(cyc_A4_div),
        .a(_T_245),
        .b(_fractA_other_PA__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6228 (
        .y(_fractB_51_PA__d),
        .sel(entering_PA),
        .a(_T_228),
        .b(_fractB_51_PA__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6229 (
        .y(_fractB_51_PB__d),
        .sel(entering_PB),
        .a(_T_288),
        .b(_fractB_51_PB__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6230 (
        .y(_fractB_51_PC__d),
        .sel(entering_PC),
        .a(_T_329),
        .b(_fractB_51_PC__q)
    );
    MUX_UNSIGNED #(.width(51)) u_mux_6231 (
        .y(_fractB_other_PA__d),
        .sel(entering_PA_normalCase),
        .a(_T_244),
        .b(_fractB_other_PA__q)
    );
    MUX_UNSIGNED #(.width(51)) u_mux_6232 (
        .y(_fractB_other_PB__d),
        .sel(entering_PB_normalCase),
        .a(_fractB_other_PA__q),
        .b(_fractB_other_PB__q)
    );
    MUX_UNSIGNED #(.width(51)) u_mux_6233 (
        .y(_fractB_other_PC__d),
        .sel(entering_PC_normalCase),
        .a(_fractB_other_PB__q),
        .b(_fractB_other_PC__q)
    );
    MUX_UNSIGNED #(.width(9)) u_mux_6234 (
        .y(_fractR0_A__d),
        .sel(_T_832),
        .a(_T_833),
        .b(_fractR0_A__q)
    );
    wire [15:0] _WTEMP_885;
    BITS #(.width(16), .high(9), .low(0)) bits_6235 (
        .y(_hiSqrR0_A_sqrt__d),
        .in(_WTEMP_885)
    );
    wire [15:0] _WTEMP_886;
    PAD_UNSIGNED #(.width(10), .n(16)) u_pad_6236 (
        .y(_WTEMP_886),
        .in(_hiSqrR0_A_sqrt__q)
    );
    MUX_UNSIGNED #(.width(16)) u_mux_6237 (
        .y(_WTEMP_885),
        .sel(cyc_A5_sqrt),
        .a(_T_834),
        .b(_WTEMP_886)
    );
    assign io_exceptionFlags = _T_1476;
    assign io_inReady_div = _T_158;
    assign io_inReady_sqrt = _T_173;
    assign io_latchMulAddA_0 = _T_888;
    assign io_latchMulAddB_0 = _T_924;
    assign io_mulAddA_0 = _T_918;
    assign io_mulAddB_0 = _T_944;
    assign io_mulAddC_2 = _T_1017;
    assign io_out = _T_1472;
    assign io_outValid_div = _T_391;
    assign io_outValid_sqrt = _T_392;
    assign io_usingMulAdd = _T_979;
    MUX_UNSIGNED #(.width(1)) u_mux_6238 (
        .y(_isNegRemT_E__d),
        .sel(cyc_E2),
        .a(_T_1052),
        .b(_isNegRemT_E__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6239 (
        .y(_isZeroRemT_E__d),
        .sel(cyc_E2),
        .a(_T_1062),
        .b(_isZeroRemT_E__q)
    );
    assign leaving_PA = _T_275;
    assign leaving_PB = _T_316;
    assign leaving_PC = _T_385;
    wire [13:0] _WTEMP_887;
    BITS #(.width(14), .high(8), .low(0)) bits_6240 (
        .y(_nextMulAdd9A_A__d),
        .in(_WTEMP_887)
    );
    wire [13:0] _WTEMP_888;
    PAD_UNSIGNED #(.width(9), .n(14)) u_pad_6241 (
        .y(_WTEMP_888),
        .in(_nextMulAdd9A_A__q)
    );
    MUX_UNSIGNED #(.width(14)) u_mux_6242 (
        .y(_WTEMP_887),
        .sel(_T_843),
        .a(_T_860),
        .b(_WTEMP_888)
    );
    MUX_UNSIGNED #(.width(9)) u_mux_6243 (
        .y(_nextMulAdd9B_A__d),
        .sel(_T_864),
        .a(_T_881),
        .b(_nextMulAdd9B_A__q)
    );
    MUX_UNSIGNED #(.width(21)) u_mux_6244 (
        .y(_partNegSigma0_A__d),
        .sel(_T_835),
        .a(_T_838),
        .b(_partNegSigma0_A__q)
    );
    assign ready_PA = _T_278;
    assign ready_PB = _T_319;
    assign ready_PC = _T_388;
    MUX_UNSIGNED #(.width(2)) u_mux_6245 (
        .y(_roundingMode_PA__d),
        .sel(entering_PA),
        .a(io_roundingMode),
        .b(_roundingMode_PA__q)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_6246 (
        .y(_roundingMode_PB__d),
        .sel(entering_PB),
        .a(_T_289),
        .b(_roundingMode_PB__q)
    );
    MUX_UNSIGNED #(.width(2)) u_mux_6247 (
        .y(_roundingMode_PC__d),
        .sel(entering_PC),
        .a(_T_330),
        .b(_roundingMode_PC__q)
    );
    MUX_UNSIGNED #(.width(53)) u_mux_6248 (
        .y(_sigT_E__d),
        .sel(cyc_C1),
        .a(_T_1048),
        .b(_sigT_E__q)
    );
    MUX_UNSIGNED #(.width(58)) u_mux_6249 (
        .y(_sigX1_B__d),
        .sel(cyc_B3),
        .a(sigXNU_B3_CX),
        .b(_sigX1_B__q)
    );
    assign sigXNU_B3_CX = _T_1022;
    MUX_UNSIGNED #(.width(58)) u_mux_6250 (
        .y(_sigXN_C__d),
        .sel(_T_1046),
        .a(sigXNU_B3_CX),
        .b(_sigXN_C__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6251 (
        .y(_sign_PA__d),
        .sel(entering_PA),
        .a(sign_S),
        .b(_sign_PA__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6252 (
        .y(_sign_PB__d),
        .sel(entering_PB),
        .a(_T_282),
        .b(_sign_PB__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6253 (
        .y(_sign_PC__d),
        .sel(entering_PC),
        .a(_T_323),
        .b(_sign_PC__q)
    );
    MUX_UNSIGNED #(.width(3)) u_mux_6254 (
        .y(_specialCodeA_PA__d),
        .sel(_T_231),
        .a(specialCodeA_S),
        .b(_specialCodeA_PA__q)
    );
    MUX_UNSIGNED #(.width(3)) u_mux_6255 (
        .y(_specialCodeA_PB__d),
        .sel(entering_PB),
        .a(_T_283),
        .b(_specialCodeA_PB__q)
    );
    MUX_UNSIGNED #(.width(3)) u_mux_6256 (
        .y(_specialCodeA_PC__d),
        .sel(entering_PC),
        .a(_T_324),
        .b(_specialCodeA_PC__q)
    );
    MUX_UNSIGNED #(.width(3)) u_mux_6257 (
        .y(_specialCodeB_PA__d),
        .sel(entering_PA),
        .a(specialCodeB_S),
        .b(_specialCodeB_PA__q)
    );
    MUX_UNSIGNED #(.width(3)) u_mux_6258 (
        .y(_specialCodeB_PB__d),
        .sel(entering_PB),
        .a(_T_286),
        .b(_specialCodeB_PB__q)
    );
    MUX_UNSIGNED #(.width(3)) u_mux_6259 (
        .y(_specialCodeB_PC__d),
        .sel(entering_PC),
        .a(_T_327),
        .b(_specialCodeB_PC__q)
    );
    MUX_UNSIGNED #(.width(33)) u_mux_6260 (
        .y(_sqrSigma1_C__d),
        .sel(cyc_B1),
        .a(sqrSigma1_B1),
        .b(_sqrSigma1_C__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6261 (
        .y(_sqrtOp_PA__d),
        .sel(entering_PA),
        .a(io_sqrtOp),
        .b(_sqrtOp_PA__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6262 (
        .y(_sqrtOp_PB__d),
        .sel(entering_PB),
        .a(_T_281),
        .b(_sqrtOp_PB__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6263 (
        .y(_sqrtOp_PC__d),
        .sel(entering_PC),
        .a(_T_322),
        .b(_sqrtOp_PC__q)
    );
    MUX_UNSIGNED #(.width(31)) u_mux_6264 (
        .y(_u_C_sqrt__d),
        .sel(cyc_C5_sqrt),
        .a(_T_1047),
        .b(_u_C_sqrt__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6265 (
        .y(_WTEMP_691),
        .sel(_T_227),
        .a(entering_PA),
        .b(_valid_PA__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6266 (
        .y(_WTEMP_692),
        .sel(_T_280),
        .a(entering_PB),
        .b(_valid_PB__q)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_6267 (
        .y(_WTEMP_693),
        .sel(_T_321),
        .a(entering_PC),
        .b(_valid_PC__q)
    );
    assign zComplSigT_C1 = _T_1040;
    assign zComplSigT_C1_sqrt = _T_1044;
    assign zSigma1_B4 = _T_1021;
endmodule //DivSqrtRecF64_mulAddZ31
module Mul54(
    input clock,
    input reset,
    input io_val_s0,
    input io_latch_a_s0,
    input [53:0] io_a_s0,
    input io_latch_b_s0,
    input [53:0] io_b_s0,
    input [104:0] io_c_s2,
    output [104:0] io_result_s3
);
    wire _val_s1__q;
    wire _val_s1__d;
    DFF_POSCLK #(.width(1)) val_s1 (
        .q(_val_s1__q),
        .d(_val_s1__d),
        .clk(clock)
    );
    wire _val_s2__q;
    wire _val_s2__d;
    DFF_POSCLK #(.width(1)) val_s2 (
        .q(_val_s2__q),
        .d(_val_s2__d),
        .clk(clock)
    );
    wire [53:0] _reg_a_s1__q;
    wire [53:0] _reg_a_s1__d;
    DFF_POSCLK #(.width(54)) reg_a_s1 (
        .q(_reg_a_s1__q),
        .d(_reg_a_s1__d),
        .clk(clock)
    );
    wire [53:0] _reg_b_s1__q;
    wire [53:0] _reg_b_s1__d;
    DFF_POSCLK #(.width(54)) reg_b_s1 (
        .q(_reg_b_s1__q),
        .d(_reg_b_s1__d),
        .clk(clock)
    );
    wire [53:0] _reg_a_s2__q;
    wire [53:0] _reg_a_s2__d;
    DFF_POSCLK #(.width(54)) reg_a_s2 (
        .q(_reg_a_s2__q),
        .d(_reg_a_s2__d),
        .clk(clock)
    );
    wire [53:0] _reg_b_s2__q;
    wire [53:0] _reg_b_s2__d;
    DFF_POSCLK #(.width(54)) reg_b_s2 (
        .q(_reg_b_s2__q),
        .d(_reg_b_s2__d),
        .clk(clock)
    );
    wire [104:0] _reg_result_s3__q;
    wire [104:0] _reg_result_s3__d;
    DFF_POSCLK #(.width(105)) reg_result_s3 (
        .q(_reg_result_s3__q),
        .d(_reg_result_s3__d),
        .clk(clock)
    );
    wire [53:0] _node_71;
    MUX_UNSIGNED #(.width(54)) u_mux_6268 (
        .y(_node_71),
        .sel(io_latch_a_s0),
        .a(io_a_s0),
        .b(_reg_a_s1__q)
    );
    wire [53:0] _node_72;
    MUX_UNSIGNED #(.width(54)) u_mux_6269 (
        .y(_node_72),
        .sel(io_latch_b_s0),
        .a(io_b_s0),
        .b(_reg_b_s1__q)
    );
    wire [107:0] _T_23;
    MUL2_UNSIGNED #(.width_a(54), .width_b(54)) u_mul2_6270 (
        .y(_T_23),
        .a(_reg_a_s2__q),
        .b(_reg_b_s2__q)
    );
    wire [104:0] _T_24;
    BITS #(.width(108), .high(104), .low(0)) bits_6271 (
        .y(_T_24),
        .in(_T_23)
    );
    wire [105:0] _T_25;
    ADD_UNSIGNED #(.width(105)) u_add_6272 (
        .y(_T_25),
        .a(_T_24),
        .b(io_c_s2)
    );
    wire [104:0] _T_26;
    TAIL #(.width(106), .n(1)) tail_6273 (
        .y(_T_26),
        .in(_T_25)
    );
    assign io_result_s3 = _reg_result_s3__q;
    MUX_UNSIGNED #(.width(54)) u_mux_6274 (
        .y(_reg_a_s1__d),
        .sel(io_val_s0),
        .a(_node_71),
        .b(_reg_a_s1__q)
    );
    MUX_UNSIGNED #(.width(54)) u_mux_6275 (
        .y(_reg_a_s2__d),
        .sel(_val_s1__q),
        .a(_reg_a_s1__q),
        .b(_reg_a_s2__q)
    );
    MUX_UNSIGNED #(.width(54)) u_mux_6276 (
        .y(_reg_b_s1__d),
        .sel(io_val_s0),
        .a(_node_72),
        .b(_reg_b_s1__q)
    );
    MUX_UNSIGNED #(.width(54)) u_mux_6277 (
        .y(_reg_b_s2__d),
        .sel(_val_s1__q),
        .a(_reg_b_s1__q),
        .b(_reg_b_s2__q)
    );
    MUX_UNSIGNED #(.width(105)) u_mux_6278 (
        .y(_reg_result_s3__d),
        .sel(_val_s2__q),
        .a(_T_26),
        .b(_reg_result_s3__q)
    );
    assign _val_s1__d = io_val_s0;
    assign _val_s2__d = _val_s1__q;
endmodule //Mul54
module RecFNToRecFN_2(
    input clock,
    input reset,
    input [64:0] io_in,
    input [1:0] io_roundingMode,
    output [32:0] io_out,
    output [4:0] io_exceptionFlags
);
    wire [11:0] _T_10;
    BITS #(.width(65), .high(63), .low(52)) bits_6290 (
        .y(_T_10),
        .in(io_in)
    );
    wire [2:0] _T_11;
    BITS #(.width(12), .high(11), .low(9)) bits_6291 (
        .y(_T_11),
        .in(_T_10)
    );
    wire _T_13;
    wire [2:0] _WTEMP_889;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_6292 (
        .y(_WTEMP_889),
        .in(1'h0)
    );
    EQ_UNSIGNED #(.width(3)) u_eq_6293 (
        .y(_T_13),
        .a(_T_11),
        .b(_WTEMP_889)
    );
    wire [1:0] _T_14;
    BITS #(.width(12), .high(11), .low(10)) bits_6294 (
        .y(_T_14),
        .in(_T_10)
    );
    wire _T_16;
    EQ_UNSIGNED #(.width(2)) u_eq_6295 (
        .y(_T_16),
        .a(_T_14),
        .b(2'h3)
    );
    wire _T_24_sign;
    wire _T_24_isNaN;
    wire _T_24_isInf;
    wire _T_24_isZero;
    wire [12:0] _T_24_sExp;
    wire [55:0] _T_24_sig;
    wire _T_31;
    BITS #(.width(65), .high(64), .low(64)) bits_6296 (
        .y(_T_31),
        .in(io_in)
    );
    wire _T_32;
    BITS #(.width(12), .high(9), .low(9)) bits_6297 (
        .y(_T_32),
        .in(_T_10)
    );
    wire _T_33;
    BITWISEAND #(.width(1)) bitwiseand_6298 (
        .y(_T_33),
        .a(_T_16),
        .b(_T_32)
    );
    wire _T_34;
    BITS #(.width(12), .high(9), .low(9)) bits_6299 (
        .y(_T_34),
        .in(_T_10)
    );
    wire _T_36;
    EQ_UNSIGNED #(.width(1)) u_eq_6300 (
        .y(_T_36),
        .a(_T_34),
        .b(1'h0)
    );
    wire _T_37;
    BITWISEAND #(.width(1)) bitwiseand_6301 (
        .y(_T_37),
        .a(_T_16),
        .b(_T_36)
    );
    wire [12:0] _T_38;
    CVT_UNSIGNED #(.width(12)) u_cvt_6302 (
        .y(_T_38),
        .in(_T_10)
    );
    wire _T_41;
    EQ_UNSIGNED #(.width(1)) u_eq_6303 (
        .y(_T_41),
        .a(_T_13),
        .b(1'h0)
    );
    wire [51:0] _T_42;
    BITS #(.width(65), .high(51), .low(0)) bits_6304 (
        .y(_T_42),
        .in(io_in)
    );
    wire [53:0] _T_44;
    CAT #(.width_a(52), .width_b(2)) cat_6305 (
        .y(_T_44),
        .a(_T_42),
        .b(2'h0)
    );
    wire [1:0] _T_45;
    CAT #(.width_a(1), .width_b(1)) cat_6306 (
        .y(_T_45),
        .a(1'h0),
        .b(_T_41)
    );
    wire [55:0] _T_46;
    CAT #(.width_a(2), .width_b(54)) cat_6307 (
        .y(_T_46),
        .a(_T_45),
        .b(_T_44)
    );
    wire [13:0] _T_48;
    wire [12:0] _WTEMP_890;
    PAD_SIGNED #(.width(12), .n(13)) s_pad_6308 (
        .y(_WTEMP_890),
        .in(-12'sh700)
    );
    ADD_SIGNED #(.width(13)) s_add_6309 (
        .y(_T_48),
        .a(_T_24_sExp),
        .b(_WTEMP_890)
    );
    wire outRawFloat_sign;
    wire outRawFloat_isNaN;
    wire outRawFloat_isInf;
    wire outRawFloat_isZero;
    wire [9:0] outRawFloat_sExp;
    wire [26:0] outRawFloat_sig;
    wire _T_63;
    wire [13:0] _WTEMP_891;
    PAD_SIGNED #(.width(1), .n(14)) s_pad_6310 (
        .y(_WTEMP_891),
        .in(1'sh0)
    );
    LT_SIGNED #(.width(14)) s_lt_6311 (
        .y(_T_63),
        .a(_T_48),
        .b(_WTEMP_891)
    );
    wire [3:0] _T_64;
    BITS #(.width(14), .high(12), .low(9)) bits_6312 (
        .y(_T_64),
        .in(_T_48)
    );
    wire _T_66;
    wire [3:0] _WTEMP_892;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_6313 (
        .y(_WTEMP_892),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(4)) u_neq_6314 (
        .y(_T_66),
        .a(_T_64),
        .b(_WTEMP_892)
    );
    wire [6:0] _T_71;
    assign _T_71 = 7'h7F;
    wire [8:0] _T_73;
    assign _T_73 = 9'h1FC;
    wire [8:0] _T_74;
    BITS #(.width(14), .high(8), .low(0)) bits_6315 (
        .y(_T_74),
        .in(_T_48)
    );
    wire [8:0] _T_75;
    MUX_UNSIGNED #(.width(9)) u_mux_6316 (
        .y(_T_75),
        .sel(_T_66),
        .a(_T_73),
        .b(_T_74)
    );
    wire [9:0] _T_76;
    CAT #(.width_a(1), .width_b(9)) cat_6317 (
        .y(_T_76),
        .a(_T_63),
        .b(_T_75)
    );
    wire [9:0] _T_77;
    ASSINT #(.width(10)) assint_6318 (
        .y(_T_77),
        .in(_T_76)
    );
    wire [25:0] _T_78;
    BITS #(.width(56), .high(55), .low(30)) bits_6319 (
        .y(_T_78),
        .in(_T_24_sig)
    );
    wire [29:0] _T_79;
    BITS #(.width(56), .high(29), .low(0)) bits_6320 (
        .y(_T_79),
        .in(_T_24_sig)
    );
    wire _T_81;
    wire [29:0] _WTEMP_893;
    PAD_UNSIGNED #(.width(1), .n(30)) u_pad_6321 (
        .y(_WTEMP_893),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(30)) u_neq_6322 (
        .y(_T_81),
        .a(_T_79),
        .b(_WTEMP_893)
    );
    wire [26:0] _T_82;
    CAT #(.width_a(26), .width_b(1)) cat_6323 (
        .y(_T_82),
        .a(_T_78),
        .b(_T_81)
    );
    wire _T_83;
    BITS #(.width(27), .high(24), .low(24)) bits_6324 (
        .y(_T_83),
        .in(outRawFloat_sig)
    );
    wire _T_85;
    EQ_UNSIGNED #(.width(1)) u_eq_6325 (
        .y(_T_85),
        .a(_T_83),
        .b(1'h0)
    );
    wire invalidExc;
    BITWISEAND #(.width(1)) bitwiseand_6326 (
        .y(invalidExc),
        .a(outRawFloat_isNaN),
        .b(_T_85)
    );
    wire _RoundRawFNToRecFN__clock;
    wire _RoundRawFNToRecFN__reset;
    wire _RoundRawFNToRecFN__io_invalidExc;
    wire _RoundRawFNToRecFN__io_infiniteExc;
    wire _RoundRawFNToRecFN__io_in_sign;
    wire _RoundRawFNToRecFN__io_in_isNaN;
    wire _RoundRawFNToRecFN__io_in_isInf;
    wire _RoundRawFNToRecFN__io_in_isZero;
    wire [9:0] _RoundRawFNToRecFN__io_in_sExp;
    wire [26:0] _RoundRawFNToRecFN__io_in_sig;
    wire [1:0] _RoundRawFNToRecFN__io_roundingMode;
    wire [32:0] _RoundRawFNToRecFN__io_out;
    wire [4:0] _RoundRawFNToRecFN__io_exceptionFlags;
    RoundRawFNToRecFN_1 RoundRawFNToRecFN (
        .clock(_RoundRawFNToRecFN__clock),
        .reset(_RoundRawFNToRecFN__reset),
        .io_invalidExc(_RoundRawFNToRecFN__io_invalidExc),
        .io_infiniteExc(_RoundRawFNToRecFN__io_infiniteExc),
        .io_in_sign(_RoundRawFNToRecFN__io_in_sign),
        .io_in_isNaN(_RoundRawFNToRecFN__io_in_isNaN),
        .io_in_isInf(_RoundRawFNToRecFN__io_in_isInf),
        .io_in_isZero(_RoundRawFNToRecFN__io_in_isZero),
        .io_in_sExp(_RoundRawFNToRecFN__io_in_sExp),
        .io_in_sig(_RoundRawFNToRecFN__io_in_sig),
        .io_roundingMode(_RoundRawFNToRecFN__io_roundingMode),
        .io_out(_RoundRawFNToRecFN__io_out),
        .io_exceptionFlags(_RoundRawFNToRecFN__io_exceptionFlags)
    );
    assign _RoundRawFNToRecFN__clock = clock;
    assign _RoundRawFNToRecFN__io_in_isInf = outRawFloat_isInf;
    assign _RoundRawFNToRecFN__io_in_isNaN = outRawFloat_isNaN;
    assign _RoundRawFNToRecFN__io_in_isZero = outRawFloat_isZero;
    assign _RoundRawFNToRecFN__io_in_sExp = outRawFloat_sExp;
    assign _RoundRawFNToRecFN__io_in_sig = outRawFloat_sig;
    assign _RoundRawFNToRecFN__io_in_sign = outRawFloat_sign;
    assign _RoundRawFNToRecFN__io_infiniteExc = 1'h0;
    assign _RoundRawFNToRecFN__io_invalidExc = invalidExc;
    assign _RoundRawFNToRecFN__io_roundingMode = io_roundingMode;
    assign _RoundRawFNToRecFN__reset = reset;
    assign _T_24_isInf = _T_37;
    assign _T_24_isNaN = _T_33;
    assign _T_24_isZero = _T_13;
    assign _T_24_sExp = _T_38;
    assign _T_24_sig = _T_46;
    assign _T_24_sign = _T_31;
    assign io_exceptionFlags = _RoundRawFNToRecFN__io_exceptionFlags;
    assign io_out = _RoundRawFNToRecFN__io_out;
    assign outRawFloat_isInf = _T_24_isInf;
    assign outRawFloat_isNaN = _T_24_isNaN;
    assign outRawFloat_isZero = _T_24_isZero;
    assign outRawFloat_sExp = _T_77;
    assign outRawFloat_sig = _T_82;
    assign outRawFloat_sign = _T_24_sign;
endmodule //RecFNToRecFN_2
module RoundRawFNToRecFN_1(
    input clock,
    input reset,
    input io_invalidExc,
    input io_infiniteExc,
    input io_in_sign,
    input io_in_isNaN,
    input io_in_isInf,
    input io_in_isZero,
    input [9:0] io_in_sExp,
    input [26:0] io_in_sig,
    input [1:0] io_roundingMode,
    output [32:0] io_out,
    output [4:0] io_exceptionFlags
);
    wire roundingMode_nearest_even;
    EQ_UNSIGNED #(.width(2)) u_eq_6327 (
        .y(roundingMode_nearest_even),
        .a(io_roundingMode),
        .b(2'h0)
    );
    wire roundingMode_minMag;
    EQ_UNSIGNED #(.width(2)) u_eq_6328 (
        .y(roundingMode_minMag),
        .a(io_roundingMode),
        .b(2'h1)
    );
    wire roundingMode_min;
    EQ_UNSIGNED #(.width(2)) u_eq_6329 (
        .y(roundingMode_min),
        .a(io_roundingMode),
        .b(2'h2)
    );
    wire roundingMode_max;
    EQ_UNSIGNED #(.width(2)) u_eq_6330 (
        .y(roundingMode_max),
        .a(io_roundingMode),
        .b(2'h3)
    );
    wire _T_26;
    BITWISEAND #(.width(1)) bitwiseand_6331 (
        .y(_T_26),
        .a(roundingMode_min),
        .b(io_in_sign)
    );
    wire _T_28;
    EQ_UNSIGNED #(.width(1)) u_eq_6332 (
        .y(_T_28),
        .a(io_in_sign),
        .b(1'h0)
    );
    wire _T_29;
    BITWISEAND #(.width(1)) bitwiseand_6333 (
        .y(_T_29),
        .a(roundingMode_max),
        .b(_T_28)
    );
    wire roundMagUp;
    BITWISEOR #(.width(1)) bitwiseor_6334 (
        .y(roundMagUp),
        .a(_T_26),
        .b(_T_29)
    );
    wire doShiftSigDown1;
    BITS #(.width(27), .high(26), .low(26)) bits_6335 (
        .y(doShiftSigDown1),
        .in(io_in_sig)
    );
    wire isNegExp;
    wire [9:0] _WTEMP_894;
    PAD_SIGNED #(.width(1), .n(10)) s_pad_6336 (
        .y(_WTEMP_894),
        .in(1'sh0)
    );
    LT_SIGNED #(.width(10)) s_lt_6337 (
        .y(isNegExp),
        .a(io_in_sExp),
        .b(_WTEMP_894)
    );
    wire _T_31;
    BITS #(.width(1), .high(0), .low(0)) bits_6338 (
        .y(_T_31),
        .in(isNegExp)
    );
    wire [24:0] _T_34;
    MUX_UNSIGNED #(.width(25)) u_mux_6339 (
        .y(_T_34),
        .sel(_T_31),
        .a(25'h1FFFFFF),
        .b(25'h0)
    );
    wire [8:0] _T_35;
    BITS #(.width(10), .high(8), .low(0)) bits_6340 (
        .y(_T_35),
        .in(io_in_sExp)
    );
    wire [8:0] _T_36;
    BITWISENOT #(.width(9)) bitwisenot_6341 (
        .y(_T_36),
        .in(_T_35)
    );
    wire _T_37;
    BITS #(.width(9), .high(8), .low(8)) bits_6342 (
        .y(_T_37),
        .in(_T_36)
    );
    wire [7:0] _T_38;
    BITS #(.width(9), .high(7), .low(0)) bits_6343 (
        .y(_T_38),
        .in(_T_36)
    );
    wire _T_39;
    BITS #(.width(8), .high(7), .low(7)) bits_6344 (
        .y(_T_39),
        .in(_T_38)
    );
    wire [6:0] _T_40;
    BITS #(.width(8), .high(6), .low(0)) bits_6345 (
        .y(_T_40),
        .in(_T_38)
    );
    wire _T_41;
    BITS #(.width(7), .high(6), .low(6)) bits_6346 (
        .y(_T_41),
        .in(_T_40)
    );
    wire [5:0] _T_42;
    BITS #(.width(7), .high(5), .low(0)) bits_6347 (
        .y(_T_42),
        .in(_T_40)
    );
    wire [64:0] _T_45;
    DSHR_SIGNED #(.width_in(65), .width_n(6)) s_dshr_6348 (
        .y(_T_45),
        .in(-65'sh10000000000000000),
        .n(_T_42)
    );
    wire [21:0] _T_46;
    BITS #(.width(65), .high(63), .low(42)) bits_6349 (
        .y(_T_46),
        .in(_T_45)
    );
    wire [15:0] _T_47;
    BITS #(.width(22), .high(15), .low(0)) bits_6350 (
        .y(_T_47),
        .in(_T_46)
    );
    wire [15:0] _T_50;
    assign _T_50 = 16'hFF00;
    wire [15:0] _T_51;
    assign _T_51 = 16'hFF;
    wire [7:0] _T_52;
    SHR_UNSIGNED #(.width(16), .n(8)) u_shr_6351 (
        .y(_T_52),
        .in(_T_47)
    );
    wire [15:0] _T_53;
    wire [15:0] _WTEMP_895;
    PAD_UNSIGNED #(.width(8), .n(16)) u_pad_6352 (
        .y(_WTEMP_895),
        .in(_T_52)
    );
    BITWISEAND #(.width(16)) bitwiseand_6353 (
        .y(_T_53),
        .a(_WTEMP_895),
        .b(_T_51)
    );
    wire [7:0] _T_54;
    BITS #(.width(16), .high(7), .low(0)) bits_6354 (
        .y(_T_54),
        .in(_T_47)
    );
    wire [15:0] _T_55;
    SHL_UNSIGNED #(.width(8), .n(8)) u_shl_6355 (
        .y(_T_55),
        .in(_T_54)
    );
    wire [15:0] _T_56;
    assign _T_56 = 16'hFF00;
    wire [15:0] _T_57;
    BITWISEAND #(.width(16)) bitwiseand_6356 (
        .y(_T_57),
        .a(_T_55),
        .b(_T_56)
    );
    wire [15:0] _T_58;
    BITWISEOR #(.width(16)) bitwiseor_6357 (
        .y(_T_58),
        .a(_T_53),
        .b(_T_57)
    );
    wire [11:0] _T_59;
    assign _T_59 = 12'hFF;
    wire [15:0] _T_60;
    assign _T_60 = 16'hFF0;
    wire [15:0] _T_61;
    assign _T_61 = 16'hF0F;
    wire [11:0] _T_62;
    SHR_UNSIGNED #(.width(16), .n(4)) u_shr_6358 (
        .y(_T_62),
        .in(_T_58)
    );
    wire [15:0] _T_63;
    wire [15:0] _WTEMP_896;
    PAD_UNSIGNED #(.width(12), .n(16)) u_pad_6359 (
        .y(_WTEMP_896),
        .in(_T_62)
    );
    BITWISEAND #(.width(16)) bitwiseand_6360 (
        .y(_T_63),
        .a(_WTEMP_896),
        .b(_T_61)
    );
    wire [11:0] _T_64;
    BITS #(.width(16), .high(11), .low(0)) bits_6361 (
        .y(_T_64),
        .in(_T_58)
    );
    wire [15:0] _T_65;
    SHL_UNSIGNED #(.width(12), .n(4)) u_shl_6362 (
        .y(_T_65),
        .in(_T_64)
    );
    wire [15:0] _T_66;
    assign _T_66 = 16'hF0F0;
    wire [15:0] _T_67;
    BITWISEAND #(.width(16)) bitwiseand_6363 (
        .y(_T_67),
        .a(_T_65),
        .b(_T_66)
    );
    wire [15:0] _T_68;
    BITWISEOR #(.width(16)) bitwiseor_6364 (
        .y(_T_68),
        .a(_T_63),
        .b(_T_67)
    );
    wire [13:0] _T_69;
    assign _T_69 = 14'hF0F;
    wire [15:0] _T_70;
    assign _T_70 = 16'h3C3C;
    wire [15:0] _T_71;
    assign _T_71 = 16'h3333;
    wire [13:0] _T_72;
    SHR_UNSIGNED #(.width(16), .n(2)) u_shr_6365 (
        .y(_T_72),
        .in(_T_68)
    );
    wire [15:0] _T_73;
    wire [15:0] _WTEMP_897;
    PAD_UNSIGNED #(.width(14), .n(16)) u_pad_6366 (
        .y(_WTEMP_897),
        .in(_T_72)
    );
    BITWISEAND #(.width(16)) bitwiseand_6367 (
        .y(_T_73),
        .a(_WTEMP_897),
        .b(_T_71)
    );
    wire [13:0] _T_74;
    BITS #(.width(16), .high(13), .low(0)) bits_6368 (
        .y(_T_74),
        .in(_T_68)
    );
    wire [15:0] _T_75;
    SHL_UNSIGNED #(.width(14), .n(2)) u_shl_6369 (
        .y(_T_75),
        .in(_T_74)
    );
    wire [15:0] _T_76;
    assign _T_76 = 16'hCCCC;
    wire [15:0] _T_77;
    BITWISEAND #(.width(16)) bitwiseand_6370 (
        .y(_T_77),
        .a(_T_75),
        .b(_T_76)
    );
    wire [15:0] _T_78;
    BITWISEOR #(.width(16)) bitwiseor_6371 (
        .y(_T_78),
        .a(_T_73),
        .b(_T_77)
    );
    wire [14:0] _T_79;
    assign _T_79 = 15'h3333;
    wire [15:0] _T_80;
    assign _T_80 = 16'h6666;
    wire [15:0] _T_81;
    assign _T_81 = 16'h5555;
    wire [14:0] _T_82;
    SHR_UNSIGNED #(.width(16), .n(1)) u_shr_6372 (
        .y(_T_82),
        .in(_T_78)
    );
    wire [15:0] _T_83;
    wire [15:0] _WTEMP_898;
    PAD_UNSIGNED #(.width(15), .n(16)) u_pad_6373 (
        .y(_WTEMP_898),
        .in(_T_82)
    );
    BITWISEAND #(.width(16)) bitwiseand_6374 (
        .y(_T_83),
        .a(_WTEMP_898),
        .b(_T_81)
    );
    wire [14:0] _T_84;
    BITS #(.width(16), .high(14), .low(0)) bits_6375 (
        .y(_T_84),
        .in(_T_78)
    );
    wire [15:0] _T_85;
    SHL_UNSIGNED #(.width(15), .n(1)) u_shl_6376 (
        .y(_T_85),
        .in(_T_84)
    );
    wire [15:0] _T_86;
    assign _T_86 = 16'hAAAA;
    wire [15:0] _T_87;
    BITWISEAND #(.width(16)) bitwiseand_6377 (
        .y(_T_87),
        .a(_T_85),
        .b(_T_86)
    );
    wire [15:0] _T_88;
    BITWISEOR #(.width(16)) bitwiseor_6378 (
        .y(_T_88),
        .a(_T_83),
        .b(_T_87)
    );
    wire [5:0] _T_89;
    BITS #(.width(22), .high(21), .low(16)) bits_6379 (
        .y(_T_89),
        .in(_T_46)
    );
    wire [3:0] _T_90;
    BITS #(.width(6), .high(3), .low(0)) bits_6380 (
        .y(_T_90),
        .in(_T_89)
    );
    wire [1:0] _T_91;
    BITS #(.width(4), .high(1), .low(0)) bits_6381 (
        .y(_T_91),
        .in(_T_90)
    );
    wire _T_92;
    BITS #(.width(2), .high(0), .low(0)) bits_6382 (
        .y(_T_92),
        .in(_T_91)
    );
    wire _T_93;
    BITS #(.width(2), .high(1), .low(1)) bits_6383 (
        .y(_T_93),
        .in(_T_91)
    );
    wire [1:0] _T_94;
    CAT #(.width_a(1), .width_b(1)) cat_6384 (
        .y(_T_94),
        .a(_T_92),
        .b(_T_93)
    );
    wire [1:0] _T_95;
    BITS #(.width(4), .high(3), .low(2)) bits_6385 (
        .y(_T_95),
        .in(_T_90)
    );
    wire _T_96;
    BITS #(.width(2), .high(0), .low(0)) bits_6386 (
        .y(_T_96),
        .in(_T_95)
    );
    wire _T_97;
    BITS #(.width(2), .high(1), .low(1)) bits_6387 (
        .y(_T_97),
        .in(_T_95)
    );
    wire [1:0] _T_98;
    CAT #(.width_a(1), .width_b(1)) cat_6388 (
        .y(_T_98),
        .a(_T_96),
        .b(_T_97)
    );
    wire [3:0] _T_99;
    CAT #(.width_a(2), .width_b(2)) cat_6389 (
        .y(_T_99),
        .a(_T_94),
        .b(_T_98)
    );
    wire [1:0] _T_100;
    BITS #(.width(6), .high(5), .low(4)) bits_6390 (
        .y(_T_100),
        .in(_T_89)
    );
    wire _T_101;
    BITS #(.width(2), .high(0), .low(0)) bits_6391 (
        .y(_T_101),
        .in(_T_100)
    );
    wire _T_102;
    BITS #(.width(2), .high(1), .low(1)) bits_6392 (
        .y(_T_102),
        .in(_T_100)
    );
    wire [1:0] _T_103;
    CAT #(.width_a(1), .width_b(1)) cat_6393 (
        .y(_T_103),
        .a(_T_101),
        .b(_T_102)
    );
    wire [5:0] _T_104;
    CAT #(.width_a(4), .width_b(2)) cat_6394 (
        .y(_T_104),
        .a(_T_99),
        .b(_T_103)
    );
    wire [21:0] _T_105;
    CAT #(.width_a(16), .width_b(6)) cat_6395 (
        .y(_T_105),
        .a(_T_88),
        .b(_T_104)
    );
    wire [21:0] _T_106;
    BITWISENOT #(.width(22)) bitwisenot_6396 (
        .y(_T_106),
        .in(_T_105)
    );
    wire [21:0] _T_107;
    wire [21:0] _WTEMP_899;
    PAD_UNSIGNED #(.width(1), .n(22)) u_pad_6397 (
        .y(_WTEMP_899),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(22)) u_mux_6398 (
        .y(_T_107),
        .sel(_T_41),
        .a(_WTEMP_899),
        .b(_T_106)
    );
    wire [21:0] _T_108;
    BITWISENOT #(.width(22)) bitwisenot_6399 (
        .y(_T_108),
        .in(_T_107)
    );
    wire [24:0] _T_110;
    CAT #(.width_a(22), .width_b(3)) cat_6400 (
        .y(_T_110),
        .a(_T_108),
        .b(3'h7)
    );
    wire _T_111;
    BITS #(.width(7), .high(6), .low(6)) bits_6401 (
        .y(_T_111),
        .in(_T_40)
    );
    wire [5:0] _T_112;
    BITS #(.width(7), .high(5), .low(0)) bits_6402 (
        .y(_T_112),
        .in(_T_40)
    );
    wire [64:0] _T_114;
    DSHR_SIGNED #(.width_in(65), .width_n(6)) s_dshr_6403 (
        .y(_T_114),
        .in(-65'sh10000000000000000),
        .n(_T_112)
    );
    wire [2:0] _T_115;
    BITS #(.width(65), .high(2), .low(0)) bits_6404 (
        .y(_T_115),
        .in(_T_114)
    );
    wire [1:0] _T_116;
    BITS #(.width(3), .high(1), .low(0)) bits_6405 (
        .y(_T_116),
        .in(_T_115)
    );
    wire _T_117;
    BITS #(.width(2), .high(0), .low(0)) bits_6406 (
        .y(_T_117),
        .in(_T_116)
    );
    wire _T_118;
    BITS #(.width(2), .high(1), .low(1)) bits_6407 (
        .y(_T_118),
        .in(_T_116)
    );
    wire [1:0] _T_119;
    CAT #(.width_a(1), .width_b(1)) cat_6408 (
        .y(_T_119),
        .a(_T_117),
        .b(_T_118)
    );
    wire _T_120;
    BITS #(.width(3), .high(2), .low(2)) bits_6409 (
        .y(_T_120),
        .in(_T_115)
    );
    wire [2:0] _T_121;
    CAT #(.width_a(2), .width_b(1)) cat_6410 (
        .y(_T_121),
        .a(_T_119),
        .b(_T_120)
    );
    wire [2:0] _T_123;
    wire [2:0] _WTEMP_900;
    PAD_UNSIGNED #(.width(1), .n(3)) u_pad_6411 (
        .y(_WTEMP_900),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(3)) u_mux_6412 (
        .y(_T_123),
        .sel(_T_111),
        .a(_T_121),
        .b(_WTEMP_900)
    );
    wire [24:0] _T_124;
    wire [24:0] _WTEMP_901;
    PAD_UNSIGNED #(.width(3), .n(25)) u_pad_6413 (
        .y(_WTEMP_901),
        .in(_T_123)
    );
    MUX_UNSIGNED #(.width(25)) u_mux_6414 (
        .y(_T_124),
        .sel(_T_39),
        .a(_T_110),
        .b(_WTEMP_901)
    );
    wire [24:0] _T_126;
    wire [24:0] _WTEMP_902;
    PAD_UNSIGNED #(.width(1), .n(25)) u_pad_6415 (
        .y(_WTEMP_902),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(25)) u_mux_6416 (
        .y(_T_126),
        .sel(_T_37),
        .a(_T_124),
        .b(_WTEMP_902)
    );
    wire [24:0] _T_127;
    BITWISEOR #(.width(25)) bitwiseor_6417 (
        .y(_T_127),
        .a(_T_34),
        .b(_T_126)
    );
    wire [24:0] _T_128;
    wire [24:0] _WTEMP_903;
    PAD_UNSIGNED #(.width(1), .n(25)) u_pad_6418 (
        .y(_WTEMP_903),
        .in(doShiftSigDown1)
    );
    BITWISEOR #(.width(25)) bitwiseor_6419 (
        .y(_T_128),
        .a(_T_127),
        .b(_WTEMP_903)
    );
    wire [26:0] roundMask;
    CAT #(.width_a(25), .width_b(2)) cat_6420 (
        .y(roundMask),
        .a(_T_128),
        .b(2'h3)
    );
    wire [27:0] _T_130;
    CAT #(.width_a(1), .width_b(27)) cat_6421 (
        .y(_T_130),
        .a(isNegExp),
        .b(roundMask)
    );
    wire [26:0] shiftedRoundMask;
    SHR_UNSIGNED #(.width(28), .n(1)) u_shr_6422 (
        .y(shiftedRoundMask),
        .in(_T_130)
    );
    wire [26:0] _T_131;
    BITWISENOT #(.width(27)) bitwisenot_6423 (
        .y(_T_131),
        .in(shiftedRoundMask)
    );
    wire [26:0] roundPosMask;
    BITWISEAND #(.width(27)) bitwiseand_6424 (
        .y(roundPosMask),
        .a(_T_131),
        .b(roundMask)
    );
    wire [26:0] _T_132;
    BITWISEAND #(.width(27)) bitwiseand_6425 (
        .y(_T_132),
        .a(io_in_sig),
        .b(roundPosMask)
    );
    wire roundPosBit;
    wire [26:0] _WTEMP_904;
    PAD_UNSIGNED #(.width(1), .n(27)) u_pad_6426 (
        .y(_WTEMP_904),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(27)) u_neq_6427 (
        .y(roundPosBit),
        .a(_T_132),
        .b(_WTEMP_904)
    );
    wire [26:0] _T_134;
    BITWISEAND #(.width(27)) bitwiseand_6428 (
        .y(_T_134),
        .a(io_in_sig),
        .b(shiftedRoundMask)
    );
    wire anyRoundExtra;
    wire [26:0] _WTEMP_905;
    PAD_UNSIGNED #(.width(1), .n(27)) u_pad_6429 (
        .y(_WTEMP_905),
        .in(1'h0)
    );
    NEQ_UNSIGNED #(.width(27)) u_neq_6430 (
        .y(anyRoundExtra),
        .a(_T_134),
        .b(_WTEMP_905)
    );
    wire anyRound;
    BITWISEOR #(.width(1)) bitwiseor_6431 (
        .y(anyRound),
        .a(roundPosBit),
        .b(anyRoundExtra)
    );
    wire _T_136;
    BITWISEAND #(.width(1)) bitwiseand_6432 (
        .y(_T_136),
        .a(roundingMode_nearest_even),
        .b(roundPosBit)
    );
    wire _T_137;
    BITWISEAND #(.width(1)) bitwiseand_6433 (
        .y(_T_137),
        .a(roundMagUp),
        .b(anyRound)
    );
    wire _T_138;
    BITWISEOR #(.width(1)) bitwiseor_6434 (
        .y(_T_138),
        .a(_T_136),
        .b(_T_137)
    );
    wire [26:0] _T_139;
    BITWISEOR #(.width(27)) bitwiseor_6435 (
        .y(_T_139),
        .a(io_in_sig),
        .b(roundMask)
    );
    wire [24:0] _T_140;
    SHR_UNSIGNED #(.width(27), .n(2)) u_shr_6436 (
        .y(_T_140),
        .in(_T_139)
    );
    wire [25:0] _T_142;
    wire [24:0] _WTEMP_906;
    PAD_UNSIGNED #(.width(1), .n(25)) u_pad_6437 (
        .y(_WTEMP_906),
        .in(1'h1)
    );
    ADD_UNSIGNED #(.width(25)) u_add_6438 (
        .y(_T_142),
        .a(_T_140),
        .b(_WTEMP_906)
    );
    wire _T_143;
    BITWISEAND #(.width(1)) bitwiseand_6439 (
        .y(_T_143),
        .a(roundingMode_nearest_even),
        .b(roundPosBit)
    );
    wire _T_145;
    EQ_UNSIGNED #(.width(1)) u_eq_6440 (
        .y(_T_145),
        .a(anyRoundExtra),
        .b(1'h0)
    );
    wire _T_146;
    BITWISEAND #(.width(1)) bitwiseand_6441 (
        .y(_T_146),
        .a(_T_143),
        .b(_T_145)
    );
    wire [25:0] _T_147;
    SHR_UNSIGNED #(.width(27), .n(1)) u_shr_6442 (
        .y(_T_147),
        .in(roundMask)
    );
    wire [25:0] _T_149;
    MUX_UNSIGNED #(.width(26)) u_mux_6443 (
        .y(_T_149),
        .sel(_T_146),
        .a(_T_147),
        .b(26'h0)
    );
    wire [25:0] _T_150;
    BITWISENOT #(.width(26)) bitwisenot_6444 (
        .y(_T_150),
        .in(_T_149)
    );
    wire [25:0] _T_151;
    BITWISEAND #(.width(26)) bitwiseand_6445 (
        .y(_T_151),
        .a(_T_142),
        .b(_T_150)
    );
    wire [26:0] _T_152;
    BITWISENOT #(.width(27)) bitwisenot_6446 (
        .y(_T_152),
        .in(roundMask)
    );
    wire [26:0] _T_153;
    BITWISEAND #(.width(27)) bitwiseand_6447 (
        .y(_T_153),
        .a(io_in_sig),
        .b(_T_152)
    );
    wire [24:0] _T_154;
    SHR_UNSIGNED #(.width(27), .n(2)) u_shr_6448 (
        .y(_T_154),
        .in(_T_153)
    );
    wire [25:0] roundedSig;
    wire [25:0] _WTEMP_907;
    PAD_UNSIGNED #(.width(25), .n(26)) u_pad_6449 (
        .y(_WTEMP_907),
        .in(_T_154)
    );
    MUX_UNSIGNED #(.width(26)) u_mux_6450 (
        .y(roundedSig),
        .sel(_T_138),
        .a(_T_151),
        .b(_WTEMP_907)
    );
    wire [1:0] _T_155;
    SHR_UNSIGNED #(.width(26), .n(24)) u_shr_6451 (
        .y(_T_155),
        .in(roundedSig)
    );
    wire [2:0] _T_156;
    CVT_UNSIGNED #(.width(2)) u_cvt_6452 (
        .y(_T_156),
        .in(_T_155)
    );
    wire [10:0] sRoundedExp;
    wire [9:0] _WTEMP_908;
    PAD_SIGNED #(.width(3), .n(10)) s_pad_6453 (
        .y(_WTEMP_908),
        .in(_T_156)
    );
    ADD_SIGNED #(.width(10)) s_add_6454 (
        .y(sRoundedExp),
        .a(io_in_sExp),
        .b(_WTEMP_908)
    );
    wire [8:0] common_expOut;
    BITS #(.width(11), .high(8), .low(0)) bits_6455 (
        .y(common_expOut),
        .in(sRoundedExp)
    );
    wire [22:0] _T_157;
    BITS #(.width(26), .high(23), .low(1)) bits_6456 (
        .y(_T_157),
        .in(roundedSig)
    );
    wire [22:0] _T_158;
    BITS #(.width(26), .high(22), .low(0)) bits_6457 (
        .y(_T_158),
        .in(roundedSig)
    );
    wire [22:0] common_fractOut;
    MUX_UNSIGNED #(.width(23)) u_mux_6458 (
        .y(common_fractOut),
        .sel(doShiftSigDown1),
        .a(_T_157),
        .b(_T_158)
    );
    wire [3:0] _T_159;
    SHR_SIGNED #(.width(11), .n(7)) s_shr_6459 (
        .y(_T_159),
        .in(sRoundedExp)
    );
    wire common_overflow;
    wire [3:0] _WTEMP_909;
    PAD_SIGNED #(.width(3), .n(4)) s_pad_6460 (
        .y(_WTEMP_909),
        .in(3'sh3)
    );
    GEQ_SIGNED #(.width(4)) s_geq_6461 (
        .y(common_overflow),
        .a(_T_159),
        .b(_WTEMP_909)
    );
    wire common_totalUnderflow;
    wire [10:0] _WTEMP_910;
    PAD_SIGNED #(.width(8), .n(11)) s_pad_6462 (
        .y(_WTEMP_910),
        .in(8'sh6B)
    );
    LT_SIGNED #(.width(11)) s_lt_6463 (
        .y(common_totalUnderflow),
        .a(sRoundedExp),
        .b(_WTEMP_910)
    );
    wire [8:0] _T_164;
    MUX_SIGNED #(.width(9)) s_mux_6464 (
        .y(_T_164),
        .sel(doShiftSigDown1),
        .a(9'sh81),
        .b(9'sh82)
    );
    wire _T_165;
    wire [9:0] _WTEMP_911;
    PAD_SIGNED #(.width(9), .n(10)) s_pad_6465 (
        .y(_WTEMP_911),
        .in(_T_164)
    );
    LT_SIGNED #(.width(10)) s_lt_6466 (
        .y(_T_165),
        .a(io_in_sExp),
        .b(_WTEMP_911)
    );
    wire common_underflow;
    BITWISEAND #(.width(1)) bitwiseand_6467 (
        .y(common_underflow),
        .a(anyRound),
        .b(_T_165)
    );
    wire isNaNOut;
    BITWISEOR #(.width(1)) bitwiseor_6468 (
        .y(isNaNOut),
        .a(io_invalidExc),
        .b(io_in_isNaN)
    );
    wire notNaN_isSpecialInfOut;
    BITWISEOR #(.width(1)) bitwiseor_6469 (
        .y(notNaN_isSpecialInfOut),
        .a(io_infiniteExc),
        .b(io_in_isInf)
    );
    wire _T_167;
    EQ_UNSIGNED #(.width(1)) u_eq_6470 (
        .y(_T_167),
        .a(isNaNOut),
        .b(1'h0)
    );
    wire _T_169;
    EQ_UNSIGNED #(.width(1)) u_eq_6471 (
        .y(_T_169),
        .a(notNaN_isSpecialInfOut),
        .b(1'h0)
    );
    wire _T_170;
    BITWISEAND #(.width(1)) bitwiseand_6472 (
        .y(_T_170),
        .a(_T_167),
        .b(_T_169)
    );
    wire _T_172;
    EQ_UNSIGNED #(.width(1)) u_eq_6473 (
        .y(_T_172),
        .a(io_in_isZero),
        .b(1'h0)
    );
    wire commonCase;
    BITWISEAND #(.width(1)) bitwiseand_6474 (
        .y(commonCase),
        .a(_T_170),
        .b(_T_172)
    );
    wire overflow;
    BITWISEAND #(.width(1)) bitwiseand_6475 (
        .y(overflow),
        .a(commonCase),
        .b(common_overflow)
    );
    wire underflow;
    BITWISEAND #(.width(1)) bitwiseand_6476 (
        .y(underflow),
        .a(commonCase),
        .b(common_underflow)
    );
    wire _T_173;
    BITWISEAND #(.width(1)) bitwiseand_6477 (
        .y(_T_173),
        .a(commonCase),
        .b(anyRound)
    );
    wire inexact;
    BITWISEOR #(.width(1)) bitwiseor_6478 (
        .y(inexact),
        .a(overflow),
        .b(_T_173)
    );
    wire overflow_roundMagUp;
    BITWISEOR #(.width(1)) bitwiseor_6479 (
        .y(overflow_roundMagUp),
        .a(roundingMode_nearest_even),
        .b(roundMagUp)
    );
    wire _T_174;
    BITWISEAND #(.width(1)) bitwiseand_6480 (
        .y(_T_174),
        .a(commonCase),
        .b(common_totalUnderflow)
    );
    wire pegMinNonzeroMagOut;
    BITWISEAND #(.width(1)) bitwiseand_6481 (
        .y(pegMinNonzeroMagOut),
        .a(_T_174),
        .b(roundMagUp)
    );
    wire _T_175;
    BITWISEAND #(.width(1)) bitwiseand_6482 (
        .y(_T_175),
        .a(commonCase),
        .b(overflow)
    );
    wire _T_177;
    EQ_UNSIGNED #(.width(1)) u_eq_6483 (
        .y(_T_177),
        .a(overflow_roundMagUp),
        .b(1'h0)
    );
    wire pegMaxFiniteMagOut;
    BITWISEAND #(.width(1)) bitwiseand_6484 (
        .y(pegMaxFiniteMagOut),
        .a(_T_175),
        .b(_T_177)
    );
    wire _T_178;
    BITWISEAND #(.width(1)) bitwiseand_6485 (
        .y(_T_178),
        .a(overflow),
        .b(overflow_roundMagUp)
    );
    wire notNaN_isInfOut;
    BITWISEOR #(.width(1)) bitwiseor_6486 (
        .y(notNaN_isInfOut),
        .a(notNaN_isSpecialInfOut),
        .b(_T_178)
    );
    wire signOut;
    MUX_UNSIGNED #(.width(1)) u_mux_6487 (
        .y(signOut),
        .sel(isNaNOut),
        .a(1'h0),
        .b(io_in_sign)
    );
    wire _T_180;
    BITWISEOR #(.width(1)) bitwiseor_6488 (
        .y(_T_180),
        .a(io_in_isZero),
        .b(common_totalUnderflow)
    );
    wire [8:0] _T_183;
    wire [8:0] _WTEMP_912;
    PAD_UNSIGNED #(.width(1), .n(9)) u_pad_6489 (
        .y(_WTEMP_912),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(9)) u_mux_6490 (
        .y(_T_183),
        .sel(_T_180),
        .a(9'h1C0),
        .b(_WTEMP_912)
    );
    wire [8:0] _T_184;
    BITWISENOT #(.width(9)) bitwisenot_6491 (
        .y(_T_184),
        .in(_T_183)
    );
    wire [8:0] _T_185;
    BITWISEAND #(.width(9)) bitwiseand_6492 (
        .y(_T_185),
        .a(common_expOut),
        .b(_T_184)
    );
    wire [8:0] _T_187;
    assign _T_187 = 9'h194;
    wire [8:0] _T_189;
    wire [8:0] _WTEMP_913;
    PAD_UNSIGNED #(.width(1), .n(9)) u_pad_6493 (
        .y(_WTEMP_913),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(9)) u_mux_6494 (
        .y(_T_189),
        .sel(pegMinNonzeroMagOut),
        .a(_T_187),
        .b(_WTEMP_913)
    );
    wire [8:0] _T_190;
    BITWISENOT #(.width(9)) bitwisenot_6495 (
        .y(_T_190),
        .in(_T_189)
    );
    wire [8:0] _T_191;
    BITWISEAND #(.width(9)) bitwiseand_6496 (
        .y(_T_191),
        .a(_T_185),
        .b(_T_190)
    );
    wire [8:0] _T_194;
    wire [8:0] _WTEMP_914;
    PAD_UNSIGNED #(.width(1), .n(9)) u_pad_6497 (
        .y(_WTEMP_914),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(9)) u_mux_6498 (
        .y(_T_194),
        .sel(pegMaxFiniteMagOut),
        .a(9'h80),
        .b(_WTEMP_914)
    );
    wire [8:0] _T_195;
    BITWISENOT #(.width(9)) bitwisenot_6499 (
        .y(_T_195),
        .in(_T_194)
    );
    wire [8:0] _T_196;
    BITWISEAND #(.width(9)) bitwiseand_6500 (
        .y(_T_196),
        .a(_T_191),
        .b(_T_195)
    );
    wire [8:0] _T_199;
    wire [8:0] _WTEMP_915;
    PAD_UNSIGNED #(.width(1), .n(9)) u_pad_6501 (
        .y(_WTEMP_915),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(9)) u_mux_6502 (
        .y(_T_199),
        .sel(notNaN_isInfOut),
        .a(9'h40),
        .b(_WTEMP_915)
    );
    wire [8:0] _T_200;
    BITWISENOT #(.width(9)) bitwisenot_6503 (
        .y(_T_200),
        .in(_T_199)
    );
    wire [8:0] _T_201;
    BITWISEAND #(.width(9)) bitwiseand_6504 (
        .y(_T_201),
        .a(_T_196),
        .b(_T_200)
    );
    wire [8:0] _T_204;
    wire [8:0] _WTEMP_916;
    PAD_UNSIGNED #(.width(1), .n(9)) u_pad_6505 (
        .y(_WTEMP_916),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(9)) u_mux_6506 (
        .y(_T_204),
        .sel(pegMinNonzeroMagOut),
        .a(9'h6B),
        .b(_WTEMP_916)
    );
    wire [8:0] _T_205;
    BITWISEOR #(.width(9)) bitwiseor_6507 (
        .y(_T_205),
        .a(_T_201),
        .b(_T_204)
    );
    wire [8:0] _T_208;
    wire [8:0] _WTEMP_917;
    PAD_UNSIGNED #(.width(1), .n(9)) u_pad_6508 (
        .y(_WTEMP_917),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(9)) u_mux_6509 (
        .y(_T_208),
        .sel(pegMaxFiniteMagOut),
        .a(9'h17F),
        .b(_WTEMP_917)
    );
    wire [8:0] _T_209;
    BITWISEOR #(.width(9)) bitwiseor_6510 (
        .y(_T_209),
        .a(_T_205),
        .b(_T_208)
    );
    wire [8:0] _T_212;
    wire [8:0] _WTEMP_918;
    PAD_UNSIGNED #(.width(1), .n(9)) u_pad_6511 (
        .y(_WTEMP_918),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(9)) u_mux_6512 (
        .y(_T_212),
        .sel(notNaN_isInfOut),
        .a(9'h180),
        .b(_WTEMP_918)
    );
    wire [8:0] _T_213;
    BITWISEOR #(.width(9)) bitwiseor_6513 (
        .y(_T_213),
        .a(_T_209),
        .b(_T_212)
    );
    wire [8:0] _T_216;
    wire [8:0] _WTEMP_919;
    PAD_UNSIGNED #(.width(1), .n(9)) u_pad_6514 (
        .y(_WTEMP_919),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(9)) u_mux_6515 (
        .y(_T_216),
        .sel(isNaNOut),
        .a(9'h1C0),
        .b(_WTEMP_919)
    );
    wire [8:0] expOut;
    BITWISEOR #(.width(9)) bitwiseor_6516 (
        .y(expOut),
        .a(_T_213),
        .b(_T_216)
    );
    wire _T_217;
    BITWISEOR #(.width(1)) bitwiseor_6517 (
        .y(_T_217),
        .a(common_totalUnderflow),
        .b(isNaNOut)
    );
    wire [22:0] _T_219;
    assign _T_219 = 23'h400000;
    wire [22:0] _T_221;
    wire [22:0] _WTEMP_920;
    PAD_UNSIGNED #(.width(1), .n(23)) u_pad_6518 (
        .y(_WTEMP_920),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(23)) u_mux_6519 (
        .y(_T_221),
        .sel(isNaNOut),
        .a(_T_219),
        .b(_WTEMP_920)
    );
    wire [22:0] _T_222;
    MUX_UNSIGNED #(.width(23)) u_mux_6520 (
        .y(_T_222),
        .sel(_T_217),
        .a(_T_221),
        .b(common_fractOut)
    );
    wire _T_223;
    BITS #(.width(1), .high(0), .low(0)) bits_6521 (
        .y(_T_223),
        .in(pegMaxFiniteMagOut)
    );
    wire [22:0] _T_226;
    MUX_UNSIGNED #(.width(23)) u_mux_6522 (
        .y(_T_226),
        .sel(_T_223),
        .a(23'h7FFFFF),
        .b(23'h0)
    );
    wire [22:0] fractOut;
    BITWISEOR #(.width(23)) bitwiseor_6523 (
        .y(fractOut),
        .a(_T_222),
        .b(_T_226)
    );
    wire [9:0] _T_227;
    CAT #(.width_a(1), .width_b(9)) cat_6524 (
        .y(_T_227),
        .a(signOut),
        .b(expOut)
    );
    wire [32:0] _T_228;
    CAT #(.width_a(10), .width_b(23)) cat_6525 (
        .y(_T_228),
        .a(_T_227),
        .b(fractOut)
    );
    wire [1:0] _T_229;
    CAT #(.width_a(1), .width_b(1)) cat_6526 (
        .y(_T_229),
        .a(underflow),
        .b(inexact)
    );
    wire [1:0] _T_230;
    CAT #(.width_a(1), .width_b(1)) cat_6527 (
        .y(_T_230),
        .a(io_invalidExc),
        .b(io_infiniteExc)
    );
    wire [2:0] _T_231;
    CAT #(.width_a(2), .width_b(1)) cat_6528 (
        .y(_T_231),
        .a(_T_230),
        .b(overflow)
    );
    wire [4:0] _T_232;
    CAT #(.width_a(3), .width_b(2)) cat_6529 (
        .y(_T_232),
        .a(_T_231),
        .b(_T_229)
    );
    assign io_exceptionFlags = _T_232;
    assign io_out = _T_228;
endmodule //RoundRawFNToRecFN_1
