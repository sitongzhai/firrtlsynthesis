module Console( // @[:@3.2]
  input        clock, // @[:@4.4]
  input        reset, // @[:@5.4]
  input        io_toggle, // @[:@6.4]
  output [7:0] io_character, // @[:@6.4]
  output [7:0] io_characterAvailable // @[:@6.4]
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  reg [8:0] pointer; // @[ConsoleTester.scala 26:24:@397.4]
  reg [8:0] arrivedPointer; // @[ConsoleTester.scala 27:31:@398.4]
  reg  lastToggle; // @[ConsoleTester.scala 28:27:@399.4]
  reg  characterArrived; // @[ConsoleTester.scala 29:33:@400.4]
  wire  gotToggle = io_toggle != lastToggle; // @[ConsoleTester.scala 31:29:@401.4]
  wire [8:0] _T_798 = 9'h184 - 9'h1; // @[ConsoleTester.scala 36:50:@407.6]
  wire  _T_799 = pointer == _T_798; // @[ConsoleTester.scala 36:28:@408.6]
  wire [8:0] _T_803 = pointer + 9'h1; // @[ConsoleTester.scala 36:70:@410.6]
  wire  _GEN_2 = gotToggle ? 1'h0 : characterArrived; // @[ConsoleTester.scala 33:3:@402.4]
  reg  _T_807; // @[Reg.scala 11:16:@415.4]
  reg  _T_809; // @[Reg.scala 11:16:@419.4]
  reg  _T_811; // @[Reg.scala 11:16:@423.4]
  reg  _T_813; // @[Reg.scala 11:16:@427.4]
  reg  _T_815; // @[Reg.scala 11:16:@431.4]
  wire  _GEN_10 = _T_815 | _GEN_2; // @[ConsoleTester.scala 41:3:@435.4]
  wire [7:0] _GEN_11 = 9'h1 == arrivedPointer ? 8'h65 : 8'h57; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_12 = 9'h2 == arrivedPointer ? 8'h20 : _GEN_11; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_13 = 9'h3 == arrivedPointer ? 8'h63 : _GEN_12; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_14 = 9'h4 == arrivedPointer ? 8'h68 : _GEN_13; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_15 = 9'h5 == arrivedPointer ? 8'h6f : _GEN_14; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_16 = 9'h6 == arrivedPointer ? 8'h6f : _GEN_15; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_17 = 9'h7 == arrivedPointer ? 8'h73 : _GEN_16; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_18 = 9'h8 == arrivedPointer ? 8'h65 : _GEN_17; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_19 = 9'h9 == arrivedPointer ? 8'h20 : _GEN_18; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_20 = 9'ha == arrivedPointer ? 8'h74 : _GEN_19; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_21 = 9'hb == arrivedPointer ? 8'h6f : _GEN_20; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_22 = 9'hc == arrivedPointer ? 8'h20 : _GEN_21; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_23 = 9'hd == arrivedPointer ? 8'h67 : _GEN_22; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_24 = 9'he == arrivedPointer ? 8'h6f : _GEN_23; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_25 = 9'hf == arrivedPointer ? 8'h20 : _GEN_24; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_26 = 9'h10 == arrivedPointer ? 8'h74 : _GEN_25; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_27 = 9'h11 == arrivedPointer ? 8'h6f : _GEN_26; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_28 = 9'h12 == arrivedPointer ? 8'h20 : _GEN_27; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_29 = 9'h13 == arrivedPointer ? 8'h74 : _GEN_28; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_30 = 9'h14 == arrivedPointer ? 8'h68 : _GEN_29; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_31 = 9'h15 == arrivedPointer ? 8'h65 : _GEN_30; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_32 = 9'h16 == arrivedPointer ? 8'h20 : _GEN_31; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_33 = 9'h17 == arrivedPointer ? 8'h6d : _GEN_32; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_34 = 9'h18 == arrivedPointer ? 8'h6f : _GEN_33; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_35 = 9'h19 == arrivedPointer ? 8'h6f : _GEN_34; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_36 = 9'h1a == arrivedPointer ? 8'h6e : _GEN_35; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_37 = 9'h1b == arrivedPointer ? 8'h2e : _GEN_36; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_38 = 9'h1c == arrivedPointer ? 8'h20 : _GEN_37; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_39 = 9'h1d == arrivedPointer ? 8'h57 : _GEN_38; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_40 = 9'h1e == arrivedPointer ? 8'h65 : _GEN_39; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_41 = 9'h1f == arrivedPointer ? 8'h20 : _GEN_40; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_42 = 9'h20 == arrivedPointer ? 8'h63 : _GEN_41; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_43 = 9'h21 == arrivedPointer ? 8'h68 : _GEN_42; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_44 = 9'h22 == arrivedPointer ? 8'h6f : _GEN_43; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_45 = 9'h23 == arrivedPointer ? 8'h6f : _GEN_44; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_46 = 9'h24 == arrivedPointer ? 8'h73 : _GEN_45; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_47 = 9'h25 == arrivedPointer ? 8'h65 : _GEN_46; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_48 = 9'h26 == arrivedPointer ? 8'h20 : _GEN_47; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_49 = 9'h27 == arrivedPointer ? 8'h74 : _GEN_48; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_50 = 9'h28 == arrivedPointer ? 8'h6f : _GEN_49; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_51 = 9'h29 == arrivedPointer ? 8'h20 : _GEN_50; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_52 = 9'h2a == arrivedPointer ? 8'h67 : _GEN_51; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_53 = 9'h2b == arrivedPointer ? 8'h6f : _GEN_52; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_54 = 9'h2c == arrivedPointer ? 8'h20 : _GEN_53; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_55 = 9'h2d == arrivedPointer ? 8'h74 : _GEN_54; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_56 = 9'h2e == arrivedPointer ? 8'h6f : _GEN_55; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_57 = 9'h2f == arrivedPointer ? 8'h20 : _GEN_56; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_58 = 9'h30 == arrivedPointer ? 8'h74 : _GEN_57; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_59 = 9'h31 == arrivedPointer ? 8'h68 : _GEN_58; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_60 = 9'h32 == arrivedPointer ? 8'h65 : _GEN_59; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_61 = 9'h33 == arrivedPointer ? 8'h20 : _GEN_60; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_62 = 9'h34 == arrivedPointer ? 8'h6d : _GEN_61; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_63 = 9'h35 == arrivedPointer ? 8'h6f : _GEN_62; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_64 = 9'h36 == arrivedPointer ? 8'h6f : _GEN_63; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_65 = 9'h37 == arrivedPointer ? 8'h6e : _GEN_64; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_66 = 9'h38 == arrivedPointer ? 8'h20 : _GEN_65; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_67 = 9'h39 == arrivedPointer ? 8'h69 : _GEN_66; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_68 = 9'h3a == arrivedPointer ? 8'h6e : _GEN_67; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_69 = 9'h3b == arrivedPointer ? 8'h20 : _GEN_68; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_70 = 9'h3c == arrivedPointer ? 8'h74 : _GEN_69; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_71 = 9'h3d == arrivedPointer ? 8'h68 : _GEN_70; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_72 = 9'h3e == arrivedPointer ? 8'h69 : _GEN_71; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_73 = 9'h3f == arrivedPointer ? 8'h73 : _GEN_72; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_74 = 9'h40 == arrivedPointer ? 8'h20 : _GEN_73; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_75 = 9'h41 == arrivedPointer ? 8'h64 : _GEN_74; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_76 = 9'h42 == arrivedPointer ? 8'h65 : _GEN_75; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_77 = 9'h43 == arrivedPointer ? 8'h63 : _GEN_76; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_78 = 9'h44 == arrivedPointer ? 8'h61 : _GEN_77; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_79 = 9'h45 == arrivedPointer ? 8'h64 : _GEN_78; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_80 = 9'h46 == arrivedPointer ? 8'h65 : _GEN_79; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_81 = 9'h47 == arrivedPointer ? 8'h20 : _GEN_80; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_82 = 9'h48 == arrivedPointer ? 8'h61 : _GEN_81; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_83 = 9'h49 == arrivedPointer ? 8'h6e : _GEN_82; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_84 = 9'h4a == arrivedPointer ? 8'h64 : _GEN_83; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_85 = 9'h4b == arrivedPointer ? 8'h20 : _GEN_84; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_86 = 9'h4c == arrivedPointer ? 8'h64 : _GEN_85; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_87 = 9'h4d == arrivedPointer ? 8'h6f : _GEN_86; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_88 = 9'h4e == arrivedPointer ? 8'h20 : _GEN_87; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_89 = 9'h4f == arrivedPointer ? 8'h74 : _GEN_88; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_90 = 9'h50 == arrivedPointer ? 8'h68 : _GEN_89; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_91 = 9'h51 == arrivedPointer ? 8'h65 : _GEN_90; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_92 = 9'h52 == arrivedPointer ? 8'h20 : _GEN_91; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_93 = 9'h53 == arrivedPointer ? 8'h6f : _GEN_92; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_94 = 9'h54 == arrivedPointer ? 8'h74 : _GEN_93; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_95 = 9'h55 == arrivedPointer ? 8'h68 : _GEN_94; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_96 = 9'h56 == arrivedPointer ? 8'h65 : _GEN_95; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_97 = 9'h57 == arrivedPointer ? 8'h72 : _GEN_96; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_98 = 9'h58 == arrivedPointer ? 8'h20 : _GEN_97; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_99 = 9'h59 == arrivedPointer ? 8'h74 : _GEN_98; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_100 = 9'h5a == arrivedPointer ? 8'h68 : _GEN_99; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_101 = 9'h5b == arrivedPointer ? 8'h69 : _GEN_100; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_102 = 9'h5c == arrivedPointer ? 8'h6e : _GEN_101; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_103 = 9'h5d == arrivedPointer ? 8'h67 : _GEN_102; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_104 = 9'h5e == arrivedPointer ? 8'h73 : _GEN_103; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_105 = 9'h5f == arrivedPointer ? 8'h2c : _GEN_104; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_106 = 9'h60 == arrivedPointer ? 8'h20 : _GEN_105; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_107 = 9'h61 == arrivedPointer ? 8'h6e : _GEN_106; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_108 = 9'h62 == arrivedPointer ? 8'h6f : _GEN_107; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_109 = 9'h63 == arrivedPointer ? 8'h74 : _GEN_108; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_110 = 9'h64 == arrivedPointer ? 8'h20 : _GEN_109; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_111 = 9'h65 == arrivedPointer ? 8'h62 : _GEN_110; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_112 = 9'h66 == arrivedPointer ? 8'h65 : _GEN_111; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_113 = 9'h67 == arrivedPointer ? 8'h63 : _GEN_112; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_114 = 9'h68 == arrivedPointer ? 8'h61 : _GEN_113; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_115 = 9'h69 == arrivedPointer ? 8'h75 : _GEN_114; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_116 = 9'h6a == arrivedPointer ? 8'h73 : _GEN_115; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_117 = 9'h6b == arrivedPointer ? 8'h65 : _GEN_116; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_118 = 9'h6c == arrivedPointer ? 8'h20 : _GEN_117; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_119 = 9'h6d == arrivedPointer ? 8'h74 : _GEN_118; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_120 = 9'h6e == arrivedPointer ? 8'h68 : _GEN_119; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_121 = 9'h6f == arrivedPointer ? 8'h65 : _GEN_120; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_122 = 9'h70 == arrivedPointer ? 8'h79 : _GEN_121; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_123 = 9'h71 == arrivedPointer ? 8'h20 : _GEN_122; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_124 = 9'h72 == arrivedPointer ? 8'h61 : _GEN_123; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_125 = 9'h73 == arrivedPointer ? 8'h72 : _GEN_124; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_126 = 9'h74 == arrivedPointer ? 8'h65 : _GEN_125; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_127 = 9'h75 == arrivedPointer ? 8'h20 : _GEN_126; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_128 = 9'h76 == arrivedPointer ? 8'h65 : _GEN_127; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_129 = 9'h77 == arrivedPointer ? 8'h61 : _GEN_128; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_130 = 9'h78 == arrivedPointer ? 8'h73 : _GEN_129; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_131 = 9'h79 == arrivedPointer ? 8'h79 : _GEN_130; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_132 = 9'h7a == arrivedPointer ? 8'h2c : _GEN_131; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_133 = 9'h7b == arrivedPointer ? 8'h20 : _GEN_132; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_134 = 9'h7c == arrivedPointer ? 8'h62 : _GEN_133; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_135 = 9'h7d == arrivedPointer ? 8'h75 : _GEN_134; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_136 = 9'h7e == arrivedPointer ? 8'h74 : _GEN_135; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_137 = 9'h7f == arrivedPointer ? 8'h20 : _GEN_136; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_138 = 9'h80 == arrivedPointer ? 8'h62 : _GEN_137; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_139 = 9'h81 == arrivedPointer ? 8'h65 : _GEN_138; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_140 = 9'h82 == arrivedPointer ? 8'h63 : _GEN_139; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_141 = 9'h83 == arrivedPointer ? 8'h61 : _GEN_140; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_142 = 9'h84 == arrivedPointer ? 8'h75 : _GEN_141; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_143 = 9'h85 == arrivedPointer ? 8'h73 : _GEN_142; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_144 = 9'h86 == arrivedPointer ? 8'h65 : _GEN_143; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_145 = 9'h87 == arrivedPointer ? 8'h20 : _GEN_144; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_146 = 9'h88 == arrivedPointer ? 8'h74 : _GEN_145; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_147 = 9'h89 == arrivedPointer ? 8'h68 : _GEN_146; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_148 = 9'h8a == arrivedPointer ? 8'h65 : _GEN_147; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_149 = 9'h8b == arrivedPointer ? 8'h79 : _GEN_148; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_150 = 9'h8c == arrivedPointer ? 8'h20 : _GEN_149; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_151 = 9'h8d == arrivedPointer ? 8'h61 : _GEN_150; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_152 = 9'h8e == arrivedPointer ? 8'h72 : _GEN_151; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_153 = 9'h8f == arrivedPointer ? 8'h65 : _GEN_152; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_154 = 9'h90 == arrivedPointer ? 8'h20 : _GEN_153; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_155 = 9'h91 == arrivedPointer ? 8'h68 : _GEN_154; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_156 = 9'h92 == arrivedPointer ? 8'h61 : _GEN_155; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_157 = 9'h93 == arrivedPointer ? 8'h72 : _GEN_156; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_158 = 9'h94 == arrivedPointer ? 8'h64 : _GEN_157; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_159 = 9'h95 == arrivedPointer ? 8'h2c : _GEN_158; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_160 = 9'h96 == arrivedPointer ? 8'h20 : _GEN_159; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_161 = 9'h97 == arrivedPointer ? 8'h62 : _GEN_160; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_162 = 9'h98 == arrivedPointer ? 8'h65 : _GEN_161; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_163 = 9'h99 == arrivedPointer ? 8'h63 : _GEN_162; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_164 = 9'h9a == arrivedPointer ? 8'h61 : _GEN_163; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_165 = 9'h9b == arrivedPointer ? 8'h75 : _GEN_164; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_166 = 9'h9c == arrivedPointer ? 8'h73 : _GEN_165; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_167 = 9'h9d == arrivedPointer ? 8'h65 : _GEN_166; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_168 = 9'h9e == arrivedPointer ? 8'h20 : _GEN_167; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_169 = 9'h9f == arrivedPointer ? 8'h74 : _GEN_168; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_170 = 9'ha0 == arrivedPointer ? 8'h68 : _GEN_169; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_171 = 9'ha1 == arrivedPointer ? 8'h61 : _GEN_170; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_172 = 9'ha2 == arrivedPointer ? 8'h74 : _GEN_171; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_173 = 9'ha3 == arrivedPointer ? 8'h20 : _GEN_172; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_174 = 9'ha4 == arrivedPointer ? 8'h67 : _GEN_173; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_175 = 9'ha5 == arrivedPointer ? 8'h6f : _GEN_174; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_176 = 9'ha6 == arrivedPointer ? 8'h61 : _GEN_175; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_177 = 9'ha7 == arrivedPointer ? 8'h6c : _GEN_176; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_178 = 9'ha8 == arrivedPointer ? 8'h20 : _GEN_177; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_179 = 9'ha9 == arrivedPointer ? 8'h77 : _GEN_178; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_180 = 9'haa == arrivedPointer ? 8'h69 : _GEN_179; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_181 = 9'hab == arrivedPointer ? 8'h6c : _GEN_180; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_182 = 9'hac == arrivedPointer ? 8'h6c : _GEN_181; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_183 = 9'had == arrivedPointer ? 8'h20 : _GEN_182; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_184 = 9'hae == arrivedPointer ? 8'h73 : _GEN_183; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_185 = 9'haf == arrivedPointer ? 8'h65 : _GEN_184; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_186 = 9'hb0 == arrivedPointer ? 8'h72 : _GEN_185; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_187 = 9'hb1 == arrivedPointer ? 8'h76 : _GEN_186; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_188 = 9'hb2 == arrivedPointer ? 8'h65 : _GEN_187; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_189 = 9'hb3 == arrivedPointer ? 8'h20 : _GEN_188; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_190 = 9'hb4 == arrivedPointer ? 8'h74 : _GEN_189; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_191 = 9'hb5 == arrivedPointer ? 8'h6f : _GEN_190; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_192 = 9'hb6 == arrivedPointer ? 8'h20 : _GEN_191; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_193 = 9'hb7 == arrivedPointer ? 8'h6f : _GEN_192; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_194 = 9'hb8 == arrivedPointer ? 8'h72 : _GEN_193; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_195 = 9'hb9 == arrivedPointer ? 8'h67 : _GEN_194; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_196 = 9'hba == arrivedPointer ? 8'h61 : _GEN_195; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_197 = 9'hbb == arrivedPointer ? 8'h6e : _GEN_196; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_198 = 9'hbc == arrivedPointer ? 8'h69 : _GEN_197; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_199 = 9'hbd == arrivedPointer ? 8'h7a : _GEN_198; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_200 = 9'hbe == arrivedPointer ? 8'h65 : _GEN_199; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_201 = 9'hbf == arrivedPointer ? 8'h20 : _GEN_200; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_202 = 9'hc0 == arrivedPointer ? 8'h61 : _GEN_201; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_203 = 9'hc1 == arrivedPointer ? 8'h6e : _GEN_202; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_204 = 9'hc2 == arrivedPointer ? 8'h64 : _GEN_203; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_205 = 9'hc3 == arrivedPointer ? 8'h20 : _GEN_204; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_206 = 9'hc4 == arrivedPointer ? 8'h6d : _GEN_205; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_207 = 9'hc5 == arrivedPointer ? 8'h65 : _GEN_206; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_208 = 9'hc6 == arrivedPointer ? 8'h61 : _GEN_207; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_209 = 9'hc7 == arrivedPointer ? 8'h73 : _GEN_208; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_210 = 9'hc8 == arrivedPointer ? 8'h75 : _GEN_209; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_211 = 9'hc9 == arrivedPointer ? 8'h72 : _GEN_210; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_212 = 9'hca == arrivedPointer ? 8'h65 : _GEN_211; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_213 = 9'hcb == arrivedPointer ? 8'h20 : _GEN_212; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_214 = 9'hcc == arrivedPointer ? 8'h74 : _GEN_213; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_215 = 9'hcd == arrivedPointer ? 8'h68 : _GEN_214; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_216 = 9'hce == arrivedPointer ? 8'h65 : _GEN_215; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_217 = 9'hcf == arrivedPointer ? 8'h20 : _GEN_216; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_218 = 9'hd0 == arrivedPointer ? 8'h62 : _GEN_217; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_219 = 9'hd1 == arrivedPointer ? 8'h65 : _GEN_218; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_220 = 9'hd2 == arrivedPointer ? 8'h73 : _GEN_219; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_221 = 9'hd3 == arrivedPointer ? 8'h74 : _GEN_220; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_222 = 9'hd4 == arrivedPointer ? 8'h20 : _GEN_221; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_223 = 9'hd5 == arrivedPointer ? 8'h6f : _GEN_222; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_224 = 9'hd6 == arrivedPointer ? 8'h66 : _GEN_223; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_225 = 9'hd7 == arrivedPointer ? 8'h20 : _GEN_224; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_226 = 9'hd8 == arrivedPointer ? 8'h6f : _GEN_225; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_227 = 9'hd9 == arrivedPointer ? 8'h75 : _GEN_226; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_228 = 9'hda == arrivedPointer ? 8'h72 : _GEN_227; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_229 = 9'hdb == arrivedPointer ? 8'h20 : _GEN_228; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_230 = 9'hdc == arrivedPointer ? 8'h65 : _GEN_229; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_231 = 9'hdd == arrivedPointer ? 8'h6e : _GEN_230; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_232 = 9'hde == arrivedPointer ? 8'h65 : _GEN_231; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_233 = 9'hdf == arrivedPointer ? 8'h72 : _GEN_232; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_234 = 9'he0 == arrivedPointer ? 8'h67 : _GEN_233; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_235 = 9'he1 == arrivedPointer ? 8'h69 : _GEN_234; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_236 = 9'he2 == arrivedPointer ? 8'h65 : _GEN_235; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_237 = 9'he3 == arrivedPointer ? 8'h73 : _GEN_236; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_238 = 9'he4 == arrivedPointer ? 8'h20 : _GEN_237; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_239 = 9'he5 == arrivedPointer ? 8'h61 : _GEN_238; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_240 = 9'he6 == arrivedPointer ? 8'h6e : _GEN_239; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_241 = 9'he7 == arrivedPointer ? 8'h64 : _GEN_240; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_242 = 9'he8 == arrivedPointer ? 8'h20 : _GEN_241; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_243 = 9'he9 == arrivedPointer ? 8'h73 : _GEN_242; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_244 = 9'hea == arrivedPointer ? 8'h6b : _GEN_243; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_245 = 9'heb == arrivedPointer ? 8'h69 : _GEN_244; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_246 = 9'hec == arrivedPointer ? 8'h6c : _GEN_245; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_247 = 9'hed == arrivedPointer ? 8'h6c : _GEN_246; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_248 = 9'hee == arrivedPointer ? 8'h73 : _GEN_247; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_249 = 9'hef == arrivedPointer ? 8'h2c : _GEN_248; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_250 = 9'hf0 == arrivedPointer ? 8'h20 : _GEN_249; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_251 = 9'hf1 == arrivedPointer ? 8'h62 : _GEN_250; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_252 = 9'hf2 == arrivedPointer ? 8'h65 : _GEN_251; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_253 = 9'hf3 == arrivedPointer ? 8'h63 : _GEN_252; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_254 = 9'hf4 == arrivedPointer ? 8'h61 : _GEN_253; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_255 = 9'hf5 == arrivedPointer ? 8'h75 : _GEN_254; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_256 = 9'hf6 == arrivedPointer ? 8'h73 : _GEN_255; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_257 = 9'hf7 == arrivedPointer ? 8'h65 : _GEN_256; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_258 = 9'hf8 == arrivedPointer ? 8'h20 : _GEN_257; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_259 = 9'hf9 == arrivedPointer ? 8'h74 : _GEN_258; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_260 = 9'hfa == arrivedPointer ? 8'h68 : _GEN_259; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_261 = 9'hfb == arrivedPointer ? 8'h61 : _GEN_260; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_262 = 9'hfc == arrivedPointer ? 8'h74 : _GEN_261; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_263 = 9'hfd == arrivedPointer ? 8'h20 : _GEN_262; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_264 = 9'hfe == arrivedPointer ? 8'h63 : _GEN_263; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_265 = 9'hff == arrivedPointer ? 8'h68 : _GEN_264; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_266 = 9'h100 == arrivedPointer ? 8'h61 : _GEN_265; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_267 = 9'h101 == arrivedPointer ? 8'h6c : _GEN_266; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_268 = 9'h102 == arrivedPointer ? 8'h6c : _GEN_267; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_269 = 9'h103 == arrivedPointer ? 8'h65 : _GEN_268; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_270 = 9'h104 == arrivedPointer ? 8'h6e : _GEN_269; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_271 = 9'h105 == arrivedPointer ? 8'h67 : _GEN_270; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_272 = 9'h106 == arrivedPointer ? 8'h65 : _GEN_271; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_273 = 9'h107 == arrivedPointer ? 8'h20 : _GEN_272; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_274 = 9'h108 == arrivedPointer ? 8'h69 : _GEN_273; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_275 = 9'h109 == arrivedPointer ? 8'h73 : _GEN_274; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_276 = 9'h10a == arrivedPointer ? 8'h20 : _GEN_275; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_277 = 9'h10b == arrivedPointer ? 8'h6f : _GEN_276; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_278 = 9'h10c == arrivedPointer ? 8'h6e : _GEN_277; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_279 = 9'h10d == arrivedPointer ? 8'h65 : _GEN_278; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_280 = 9'h10e == arrivedPointer ? 8'h20 : _GEN_279; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_281 = 9'h10f == arrivedPointer ? 8'h74 : _GEN_280; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_282 = 9'h110 == arrivedPointer ? 8'h68 : _GEN_281; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_283 = 9'h111 == arrivedPointer ? 8'h61 : _GEN_282; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_284 = 9'h112 == arrivedPointer ? 8'h74 : _GEN_283; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_285 = 9'h113 == arrivedPointer ? 8'h20 : _GEN_284; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_286 = 9'h114 == arrivedPointer ? 8'h77 : _GEN_285; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_287 = 9'h115 == arrivedPointer ? 8'h65 : _GEN_286; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_288 = 9'h116 == arrivedPointer ? 8'h20 : _GEN_287; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_289 = 9'h117 == arrivedPointer ? 8'h61 : _GEN_288; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_290 = 9'h118 == arrivedPointer ? 8'h72 : _GEN_289; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_291 = 9'h119 == arrivedPointer ? 8'h65 : _GEN_290; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_292 = 9'h11a == arrivedPointer ? 8'h20 : _GEN_291; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_293 = 9'h11b == arrivedPointer ? 8'h77 : _GEN_292; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_294 = 9'h11c == arrivedPointer ? 8'h69 : _GEN_293; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_295 = 9'h11d == arrivedPointer ? 8'h6c : _GEN_294; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_296 = 9'h11e == arrivedPointer ? 8'h6c : _GEN_295; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_297 = 9'h11f == arrivedPointer ? 8'h69 : _GEN_296; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_298 = 9'h120 == arrivedPointer ? 8'h6e : _GEN_297; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_299 = 9'h121 == arrivedPointer ? 8'h67 : _GEN_298; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_300 = 9'h122 == arrivedPointer ? 8'h20 : _GEN_299; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_301 = 9'h123 == arrivedPointer ? 8'h74 : _GEN_300; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_302 = 9'h124 == arrivedPointer ? 8'h6f : _GEN_301; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_303 = 9'h125 == arrivedPointer ? 8'h20 : _GEN_302; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_304 = 9'h126 == arrivedPointer ? 8'h61 : _GEN_303; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_305 = 9'h127 == arrivedPointer ? 8'h63 : _GEN_304; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_306 = 9'h128 == arrivedPointer ? 8'h63 : _GEN_305; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_307 = 9'h129 == arrivedPointer ? 8'h65 : _GEN_306; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_308 = 9'h12a == arrivedPointer ? 8'h70 : _GEN_307; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_309 = 9'h12b == arrivedPointer ? 8'h74 : _GEN_308; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_310 = 9'h12c == arrivedPointer ? 8'h2c : _GEN_309; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_311 = 9'h12d == arrivedPointer ? 8'h20 : _GEN_310; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_312 = 9'h12e == arrivedPointer ? 8'h6f : _GEN_311; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_313 = 9'h12f == arrivedPointer ? 8'h6e : _GEN_312; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_314 = 9'h130 == arrivedPointer ? 8'h65 : _GEN_313; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_315 = 9'h131 == arrivedPointer ? 8'h20 : _GEN_314; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_316 = 9'h132 == arrivedPointer ? 8'h77 : _GEN_315; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_317 = 9'h133 == arrivedPointer ? 8'h65 : _GEN_316; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_318 = 9'h134 == arrivedPointer ? 8'h20 : _GEN_317; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_319 = 9'h135 == arrivedPointer ? 8'h61 : _GEN_318; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_320 = 9'h136 == arrivedPointer ? 8'h72 : _GEN_319; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_321 = 9'h137 == arrivedPointer ? 8'h65 : _GEN_320; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_322 = 9'h138 == arrivedPointer ? 8'h20 : _GEN_321; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_323 = 9'h139 == arrivedPointer ? 8'h75 : _GEN_322; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_324 = 9'h13a == arrivedPointer ? 8'h6e : _GEN_323; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_325 = 9'h13b == arrivedPointer ? 8'h77 : _GEN_324; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_326 = 9'h13c == arrivedPointer ? 8'h69 : _GEN_325; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_327 = 9'h13d == arrivedPointer ? 8'h6c : _GEN_326; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_328 = 9'h13e == arrivedPointer ? 8'h6c : _GEN_327; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_329 = 9'h13f == arrivedPointer ? 8'h69 : _GEN_328; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_330 = 9'h140 == arrivedPointer ? 8'h6e : _GEN_329; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_331 = 9'h141 == arrivedPointer ? 8'h67 : _GEN_330; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_332 = 9'h142 == arrivedPointer ? 8'h20 : _GEN_331; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_333 = 9'h143 == arrivedPointer ? 8'h74 : _GEN_332; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_334 = 9'h144 == arrivedPointer ? 8'h6f : _GEN_333; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_335 = 9'h145 == arrivedPointer ? 8'h20 : _GEN_334; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_336 = 9'h146 == arrivedPointer ? 8'h70 : _GEN_335; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_337 = 9'h147 == arrivedPointer ? 8'h6f : _GEN_336; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_338 = 9'h148 == arrivedPointer ? 8'h73 : _GEN_337; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_339 = 9'h149 == arrivedPointer ? 8'h74 : _GEN_338; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_340 = 9'h14a == arrivedPointer ? 8'h70 : _GEN_339; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_341 = 9'h14b == arrivedPointer ? 8'h6f : _GEN_340; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_342 = 9'h14c == arrivedPointer ? 8'h6e : _GEN_341; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_343 = 9'h14d == arrivedPointer ? 8'h65 : _GEN_342; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_344 = 9'h14e == arrivedPointer ? 8'h2c : _GEN_343; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_345 = 9'h14f == arrivedPointer ? 8'h20 : _GEN_344; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_346 = 9'h150 == arrivedPointer ? 8'h61 : _GEN_345; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_347 = 9'h151 == arrivedPointer ? 8'h6e : _GEN_346; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_348 = 9'h152 == arrivedPointer ? 8'h64 : _GEN_347; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_349 = 9'h153 == arrivedPointer ? 8'h20 : _GEN_348; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_350 = 9'h154 == arrivedPointer ? 8'h6f : _GEN_349; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_351 = 9'h155 == arrivedPointer ? 8'h6e : _GEN_350; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_352 = 9'h156 == arrivedPointer ? 8'h65 : _GEN_351; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_353 = 9'h157 == arrivedPointer ? 8'h20 : _GEN_352; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_354 = 9'h158 == arrivedPointer ? 8'h77 : _GEN_353; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_355 = 9'h159 == arrivedPointer ? 8'h68 : _GEN_354; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_356 = 9'h15a == arrivedPointer ? 8'h69 : _GEN_355; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_357 = 9'h15b == arrivedPointer ? 8'h63 : _GEN_356; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_358 = 9'h15c == arrivedPointer ? 8'h68 : _GEN_357; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_359 = 9'h15d == arrivedPointer ? 8'h20 : _GEN_358; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_360 = 9'h15e == arrivedPointer ? 8'h77 : _GEN_359; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_361 = 9'h15f == arrivedPointer ? 8'h65 : _GEN_360; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_362 = 9'h160 == arrivedPointer ? 8'h20 : _GEN_361; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_363 = 9'h161 == arrivedPointer ? 8'h69 : _GEN_362; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_364 = 9'h162 == arrivedPointer ? 8'h6e : _GEN_363; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_365 = 9'h163 == arrivedPointer ? 8'h74 : _GEN_364; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_366 = 9'h164 == arrivedPointer ? 8'h65 : _GEN_365; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_367 = 9'h165 == arrivedPointer ? 8'h6e : _GEN_366; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_368 = 9'h166 == arrivedPointer ? 8'h64 : _GEN_367; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_369 = 9'h167 == arrivedPointer ? 8'h20 : _GEN_368; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_370 = 9'h168 == arrivedPointer ? 8'h74 : _GEN_369; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_371 = 9'h169 == arrivedPointer ? 8'h6f : _GEN_370; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_372 = 9'h16a == arrivedPointer ? 8'h20 : _GEN_371; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_373 = 9'h16b == arrivedPointer ? 8'h77 : _GEN_372; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_374 = 9'h16c == arrivedPointer ? 8'h69 : _GEN_373; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_375 = 9'h16d == arrivedPointer ? 8'h6e : _GEN_374; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_376 = 9'h16e == arrivedPointer ? 8'h2c : _GEN_375; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_377 = 9'h16f == arrivedPointer ? 8'h20 : _GEN_376; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_378 = 9'h170 == arrivedPointer ? 8'h61 : _GEN_377; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_379 = 9'h171 == arrivedPointer ? 8'h6e : _GEN_378; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_380 = 9'h172 == arrivedPointer ? 8'h64 : _GEN_379; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_381 = 9'h173 == arrivedPointer ? 8'h20 : _GEN_380; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_382 = 9'h174 == arrivedPointer ? 8'h74 : _GEN_381; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_383 = 9'h175 == arrivedPointer ? 8'h68 : _GEN_382; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_384 = 9'h176 == arrivedPointer ? 8'h65 : _GEN_383; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_385 = 9'h177 == arrivedPointer ? 8'h20 : _GEN_384; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_386 = 9'h178 == arrivedPointer ? 8'h6f : _GEN_385; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_387 = 9'h179 == arrivedPointer ? 8'h74 : _GEN_386; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_388 = 9'h17a == arrivedPointer ? 8'h68 : _GEN_387; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_389 = 9'h17b == arrivedPointer ? 8'h65 : _GEN_388; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_390 = 9'h17c == arrivedPointer ? 8'h72 : _GEN_389; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_391 = 9'h17d == arrivedPointer ? 8'h73 : _GEN_390; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_392 = 9'h17e == arrivedPointer ? 8'h2c : _GEN_391; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_393 = 9'h17f == arrivedPointer ? 8'h20 : _GEN_392; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_394 = 9'h180 == arrivedPointer ? 8'h74 : _GEN_393; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_395 = 9'h181 == arrivedPointer ? 8'h6f : _GEN_394; // @[ConsoleTester.scala 45:16:@438.4]
  wire [7:0] _GEN_396 = 9'h182 == arrivedPointer ? 8'h6f : _GEN_395; // @[ConsoleTester.scala 45:16:@438.4]
  assign io_character = 9'h183 == arrivedPointer ? 8'h2e : _GEN_396; // @[ConsoleTester.scala 45:16:@438.4]
  assign io_characterAvailable = {{7'd0}, characterArrived};
  always @(posedge clock) begin
    if (reset) begin
      pointer <= 9'h0;
    end else if (gotToggle) begin // @[ConsoleTester.scala 33:3:@402.4]
      if (_T_799) begin // @[ConsoleTester.scala 36:19:@411.6]
        pointer <= 9'h0;
      end else begin
        pointer <= _T_803;
      end
    end
    if (reset) begin
      arrivedPointer <= 9'h0;
    end else if (gotToggle) begin // @[ConsoleTester.scala 33:3:@402.4]
      arrivedPointer <= pointer;
    end
    if (reset) begin
      lastToggle <= 1'h0;
    end else if (gotToggle) begin // @[ConsoleTester.scala 33:3:@402.4]
      lastToggle <= io_toggle;
    end
    if (reset) begin
      characterArrived <= 1'h0;
    end else begin
      characterArrived <= _GEN_10;
    end
    _T_807 <= io_toggle != lastToggle; // @[ConsoleTester.scala 31:29:@401.4]
    _T_809 <= _T_807; // @[Reg.scala 12:19:@420.4]
    _T_811 <= _T_809; // @[Reg.scala 12:19:@424.4]
    _T_813 <= _T_811; // @[Reg.scala 12:19:@428.4]
    _T_815 <= _T_813; // @[Reg.scala 12:19:@432.4]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pointer = _RAND_0[8:0];
  _RAND_1 = {1{`RANDOM}};
  arrivedPointer = _RAND_1[8:0];
  _RAND_2 = {1{`RANDOM}};
  lastToggle = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  characterArrived = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  _T_807 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  _T_809 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  _T_811 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  _T_813 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  _T_815 = _RAND_8[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
