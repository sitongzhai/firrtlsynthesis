module RouterUnitTester(
    input clock,
    input reset
);
    wire _c__clock;
    wire _c__reset;
    wire _c__io_read_routing_table_request_ready;
    wire _c__io_read_routing_table_request_valid;
    wire [31:0] _c__io_read_routing_table_request_bits_addr;
    wire _c__io_read_routing_table_response_ready;
    wire _c__io_read_routing_table_response_valid;
    wire [31:0] _c__io_read_routing_table_response_bits;
    wire _c__io_load_routing_table_request_ready;
    wire _c__io_load_routing_table_request_valid;
    wire [31:0] _c__io_load_routing_table_request_bits_addr;
    wire [31:0] _c__io_load_routing_table_request_bits_data;
    wire _c__io_in_ready;
    wire _c__io_in_valid;
    wire [7:0] _c__io_in_bits_header;
    wire [63:0] _c__io_in_bits_body;
    wire _c__io_outs_0_ready;
    wire _c__io_outs_0_valid;
    wire [7:0] _c__io_outs_0_bits_header;
    wire [63:0] _c__io_outs_0_bits_body;
    wire _c__io_outs_1_ready;
    wire _c__io_outs_1_valid;
    wire [7:0] _c__io_outs_1_bits_header;
    wire [63:0] _c__io_outs_1_bits_body;
    wire _c__io_outs_2_ready;
    wire _c__io_outs_2_valid;
    wire [7:0] _c__io_outs_2_bits_header;
    wire [63:0] _c__io_outs_2_bits_body;
    wire _c__io_outs_3_ready;
    wire _c__io_outs_3_valid;
    wire [7:0] _c__io_outs_3_bits_header;
    wire [63:0] _c__io_outs_3_bits_body;
    Router c (
        .clock(_c__clock),
        .reset(_c__reset),
        .io_read_routing_table_request_ready(_c__io_read_routing_table_request_ready),
        .io_read_routing_table_request_valid(_c__io_read_routing_table_request_valid),
        .io_read_routing_table_request_bits_addr(_c__io_read_routing_table_request_bits_addr),
        .io_read_routing_table_response_ready(_c__io_read_routing_table_response_ready),
        .io_read_routing_table_response_valid(_c__io_read_routing_table_response_valid),
        .io_read_routing_table_response_bits(_c__io_read_routing_table_response_bits),
        .io_load_routing_table_request_ready(_c__io_load_routing_table_request_ready),
        .io_load_routing_table_request_valid(_c__io_load_routing_table_request_valid),
        .io_load_routing_table_request_bits_addr(_c__io_load_routing_table_request_bits_addr),
        .io_load_routing_table_request_bits_data(_c__io_load_routing_table_request_bits_data),
        .io_in_ready(_c__io_in_ready),
        .io_in_valid(_c__io_in_valid),
        .io_in_bits_header(_c__io_in_bits_header),
        .io_in_bits_body(_c__io_in_bits_body),
        .io_outs_0_ready(_c__io_outs_0_ready),
        .io_outs_0_valid(_c__io_outs_0_valid),
        .io_outs_0_bits_header(_c__io_outs_0_bits_header),
        .io_outs_0_bits_body(_c__io_outs_0_bits_body),
        .io_outs_1_ready(_c__io_outs_1_ready),
        .io_outs_1_valid(_c__io_outs_1_valid),
        .io_outs_1_bits_header(_c__io_outs_1_bits_header),
        .io_outs_1_bits_body(_c__io_outs_1_bits_body),
        .io_outs_2_ready(_c__io_outs_2_ready),
        .io_outs_2_valid(_c__io_outs_2_valid),
        .io_outs_2_bits_header(_c__io_outs_2_bits_header),
        .io_outs_2_bits_body(_c__io_outs_2_bits_body),
        .io_outs_3_ready(_c__io_outs_3_ready),
        .io_outs_3_valid(_c__io_outs_3_valid),
        .io_outs_3_bits_header(_c__io_outs_3_bits_header),
        .io_outs_3_bits_body(_c__io_outs_3_bits_body)
    );
    wire [7:0] __T_4__q;
    wire [7:0] __T_4__d;
    DFF_POSCLK #(.width(8)) _T_4 (
        .q(__T_4__q),
        .d(__T_4__d),
        .clk(clock)
    );
    wire [7:0] _WTEMP_4;
    MUX_UNSIGNED #(.width(8)) u_mux_105 (
        .y(__T_4__d),
        .sel(reset),
        .a(8'h0),
        .b(_WTEMP_4)
    );
    wire __T_7__q;
    wire __T_7__d;
    DFF_POSCLK #(.width(1)) _T_7 (
        .q(__T_7__q),
        .d(__T_7__d),
        .clk(clock)
    );
    wire _WTEMP_5;
    MUX_UNSIGNED #(.width(1)) u_mux_106 (
        .y(__T_7__d),
        .sel(reset),
        .a(1'h0),
        .b(_WTEMP_5)
    );
    wire [7:0] __T_10__q;
    wire [7:0] __T_10__d;
    DFF_POSCLK #(.width(8)) _T_10 (
        .q(__T_10__q),
        .d(__T_10__d),
        .clk(clock)
    );
    wire [7:0] _WTEMP_6;
    MUX_UNSIGNED #(.width(8)) u_mux_107 (
        .y(__T_10__d),
        .sel(reset),
        .a(8'h0),
        .b(_WTEMP_6)
    );
    wire __T_13__q;
    wire __T_13__d;
    DFF_POSCLK #(.width(1)) _T_13 (
        .q(__T_13__q),
        .d(__T_13__d),
        .clk(clock)
    );
    wire _WTEMP_7;
    MUX_UNSIGNED #(.width(1)) u_mux_108 (
        .y(__T_13__d),
        .sel(reset),
        .a(1'h0),
        .b(_WTEMP_7)
    );
    wire _T_14;
    BITWISEAND #(.width(1)) bitwiseand_109 (
        .y(_T_14),
        .a(__T_7__q),
        .b(__T_13__q)
    );
    wire _T_16;
    EQ_UNSIGNED #(.width(1)) u_eq_110 (
        .y(_T_16),
        .a(reset),
        .b(1'h0)
    );
    wire _T_18;
    EQ_UNSIGNED #(.width(1)) u_eq_111 (
        .y(_T_18),
        .a(reset),
        .b(1'h0)
    );
    wire [13:0] __T_21__q;
    wire [13:0] __T_21__d;
    DFF_POSCLK #(.width(14)) _T_21 (
        .q(__T_21__q),
        .d(__T_21__d),
        .clk(clock)
    );
    wire [13:0] _WTEMP_8;
    MUX_UNSIGNED #(.width(14)) u_mux_112 (
        .y(__T_21__d),
        .sel(reset),
        .a(14'h0),
        .b(_WTEMP_8)
    );
    wire [14:0] _T_23;
    wire [13:0] _WTEMP_9;
    PAD_UNSIGNED #(.width(1), .n(14)) u_pad_113 (
        .y(_WTEMP_9),
        .in(1'h1)
    );
    ADD_UNSIGNED #(.width(14)) u_add_114 (
        .y(_T_23),
        .a(__T_21__q),
        .b(_WTEMP_9)
    );
    wire [13:0] _T_24;
    TAIL #(.width(15), .n(1)) tail_115 (
        .y(_T_24),
        .in(_T_23)
    );
    wire _T_26;
    GT_UNSIGNED #(.width(14)) u_gt_116 (
        .y(_T_26),
        .a(__T_21__q),
        .b(14'h2710)
    );
    wire _T_29;
    EQ_UNSIGNED #(.width(1)) u_eq_117 (
        .y(_T_29),
        .a(reset),
        .b(1'h0)
    );
    wire _T_31;
    EQ_UNSIGNED #(.width(1)) u_eq_118 (
        .y(_T_31),
        .a(reset),
        .b(1'h0)
    );
    wire _T_87_0;
    wire _T_87_1;
    wire _T_87_2;
    wire _T_87_3;
    wire _T_87_4;
    wire _T_87_5;
    wire _T_87_6;
    wire _T_87_7;
    wire _T_87_8;
    wire _T_87_9;
    wire _T_87_10;
    wire _T_87_11;
    wire _T_87_12;
    wire _T_87_13;
    wire _T_87_14;
    wire _T_87_15;
    wire _T_87_16;
    wire _T_87_17;
    wire _T_87_18;
    wire _T_87_19;
    wire _T_87_20;
    wire _T_87_21;
    wire _T_87_22;
    wire _T_87_23;
    wire _T_87_24;
    wire _T_87_25;
    wire _T_87_26;
    wire _T_87_27;
    wire _T_87_28;
    wire _T_87_29;
    wire _T_87_30;
    wire _T_87_31;
    wire _T_87_32;
    wire _T_87_33;
    wire _T_87_34;
    wire _T_87_35;
    wire _T_87_36;
    wire _T_87_37;
    wire _T_87_38;
    wire _T_87_39;
    wire _T_87_40;
    wire _T_87_41;
    wire _T_87_42;
    wire _T_87_43;
    wire _T_87_44;
    wire _T_87_45;
    wire _T_87_46;
    wire _T_87_47;
    wire _T_87_48;
    wire _T_87_49;
    wire _T_87_50;
    wire _T_87_51;
    wire _T_87_52;
    wire [3:0] _value__q;
    wire [3:0] _value__d;
    DFF_POSCLK #(.width(4)) value (
        .q(_value__q),
        .d(_value__d),
        .clk(clock)
    );
    wire [3:0] _WTEMP_10;
    MUX_UNSIGNED #(.width(4)) u_mux_119 (
        .y(_value__d),
        .sel(reset),
        .a(4'h0),
        .b(_WTEMP_10)
    );
    wire [1:0] _T_157_0;
    wire [1:0] _T_157_1;
    wire [1:0] _T_157_2;
    wire [1:0] _T_157_3;
    wire [1:0] _T_157_4;
    wire [1:0] _T_157_5;
    wire [1:0] _T_157_6;
    wire [1:0] _T_157_7;
    wire [1:0] _T_157_8;
    wire [1:0] _T_157_9;
    wire _node_105;
    EQ_UNSIGNED #(.width(4)) u_eq_120 (
        .y(_node_105),
        .a(4'd0),
        .b(_value__q)
    );
    wire [1:0] _node_106;
    assign _node_106 = _T_157_0;
    wire _node_107;
    EQ_UNSIGNED #(.width(4)) u_eq_121 (
        .y(_node_107),
        .a(4'd1),
        .b(_value__q)
    );
    wire [1:0] _node_108;
    MUX_UNSIGNED #(.width(2)) u_mux_122 (
        .y(_node_108),
        .sel(_node_107),
        .a(_T_157_1),
        .b(_node_106)
    );
    wire _node_109;
    EQ_UNSIGNED #(.width(4)) u_eq_123 (
        .y(_node_109),
        .a(4'd2),
        .b(_value__q)
    );
    wire [1:0] _node_110;
    MUX_UNSIGNED #(.width(2)) u_mux_124 (
        .y(_node_110),
        .sel(_node_109),
        .a(_T_157_2),
        .b(_node_108)
    );
    wire _node_111;
    EQ_UNSIGNED #(.width(4)) u_eq_125 (
        .y(_node_111),
        .a(4'd3),
        .b(_value__q)
    );
    wire [1:0] _node_112;
    MUX_UNSIGNED #(.width(2)) u_mux_126 (
        .y(_node_112),
        .sel(_node_111),
        .a(_T_157_3),
        .b(_node_110)
    );
    wire _node_113;
    EQ_UNSIGNED #(.width(4)) u_eq_127 (
        .y(_node_113),
        .a(4'd4),
        .b(_value__q)
    );
    wire [1:0] _node_114;
    MUX_UNSIGNED #(.width(2)) u_mux_128 (
        .y(_node_114),
        .sel(_node_113),
        .a(_T_157_4),
        .b(_node_112)
    );
    wire _node_115;
    EQ_UNSIGNED #(.width(4)) u_eq_129 (
        .y(_node_115),
        .a(4'd5),
        .b(_value__q)
    );
    wire [1:0] _node_116;
    MUX_UNSIGNED #(.width(2)) u_mux_130 (
        .y(_node_116),
        .sel(_node_115),
        .a(_T_157_5),
        .b(_node_114)
    );
    wire _node_117;
    EQ_UNSIGNED #(.width(4)) u_eq_131 (
        .y(_node_117),
        .a(4'd6),
        .b(_value__q)
    );
    wire [1:0] _node_118;
    MUX_UNSIGNED #(.width(2)) u_mux_132 (
        .y(_node_118),
        .sel(_node_117),
        .a(_T_157_6),
        .b(_node_116)
    );
    wire _node_119;
    EQ_UNSIGNED #(.width(4)) u_eq_133 (
        .y(_node_119),
        .a(4'd7),
        .b(_value__q)
    );
    wire [1:0] _node_120;
    MUX_UNSIGNED #(.width(2)) u_mux_134 (
        .y(_node_120),
        .sel(_node_119),
        .a(_T_157_7),
        .b(_node_118)
    );
    wire _node_121;
    EQ_UNSIGNED #(.width(4)) u_eq_135 (
        .y(_node_121),
        .a(4'd8),
        .b(_value__q)
    );
    wire [1:0] _node_122;
    MUX_UNSIGNED #(.width(2)) u_mux_136 (
        .y(_node_122),
        .sel(_node_121),
        .a(_T_157_8),
        .b(_node_120)
    );
    wire _node_123;
    EQ_UNSIGNED #(.width(4)) u_eq_137 (
        .y(_node_123),
        .a(4'd9),
        .b(_value__q)
    );
    wire [1:0] _node_124;
    MUX_UNSIGNED #(.width(2)) u_mux_138 (
        .y(_node_124),
        .sel(_node_123),
        .a(_T_157_9),
        .b(_node_122)
    );
    wire [5:0] _T_172;
    BITS #(.width(8), .high(5), .low(0)) bits_139 (
        .y(_T_172),
        .in(__T_4__q)
    );
    wire _node_125;
    EQ_UNSIGNED #(.width(6)) u_eq_140 (
        .y(_node_125),
        .a(6'd0),
        .b(_T_172)
    );
    wire _node_126;
    assign _node_126 = _T_87_0;
    wire _node_127;
    EQ_UNSIGNED #(.width(6)) u_eq_141 (
        .y(_node_127),
        .a(6'd1),
        .b(_T_172)
    );
    wire _node_128;
    MUX_UNSIGNED #(.width(1)) u_mux_142 (
        .y(_node_128),
        .sel(_node_127),
        .a(_T_87_1),
        .b(_node_126)
    );
    wire _node_129;
    EQ_UNSIGNED #(.width(6)) u_eq_143 (
        .y(_node_129),
        .a(6'd2),
        .b(_T_172)
    );
    wire _node_130;
    MUX_UNSIGNED #(.width(1)) u_mux_144 (
        .y(_node_130),
        .sel(_node_129),
        .a(_T_87_2),
        .b(_node_128)
    );
    wire _node_131;
    EQ_UNSIGNED #(.width(6)) u_eq_145 (
        .y(_node_131),
        .a(6'd3),
        .b(_T_172)
    );
    wire _node_132;
    MUX_UNSIGNED #(.width(1)) u_mux_146 (
        .y(_node_132),
        .sel(_node_131),
        .a(_T_87_3),
        .b(_node_130)
    );
    wire _node_133;
    EQ_UNSIGNED #(.width(6)) u_eq_147 (
        .y(_node_133),
        .a(6'd4),
        .b(_T_172)
    );
    wire _node_134;
    MUX_UNSIGNED #(.width(1)) u_mux_148 (
        .y(_node_134),
        .sel(_node_133),
        .a(_T_87_4),
        .b(_node_132)
    );
    wire _node_135;
    EQ_UNSIGNED #(.width(6)) u_eq_149 (
        .y(_node_135),
        .a(6'd5),
        .b(_T_172)
    );
    wire _node_136;
    MUX_UNSIGNED #(.width(1)) u_mux_150 (
        .y(_node_136),
        .sel(_node_135),
        .a(_T_87_5),
        .b(_node_134)
    );
    wire _node_137;
    EQ_UNSIGNED #(.width(6)) u_eq_151 (
        .y(_node_137),
        .a(6'd6),
        .b(_T_172)
    );
    wire _node_138;
    MUX_UNSIGNED #(.width(1)) u_mux_152 (
        .y(_node_138),
        .sel(_node_137),
        .a(_T_87_6),
        .b(_node_136)
    );
    wire _node_139;
    EQ_UNSIGNED #(.width(6)) u_eq_153 (
        .y(_node_139),
        .a(6'd7),
        .b(_T_172)
    );
    wire _node_140;
    MUX_UNSIGNED #(.width(1)) u_mux_154 (
        .y(_node_140),
        .sel(_node_139),
        .a(_T_87_7),
        .b(_node_138)
    );
    wire _node_141;
    EQ_UNSIGNED #(.width(6)) u_eq_155 (
        .y(_node_141),
        .a(6'd8),
        .b(_T_172)
    );
    wire _node_142;
    MUX_UNSIGNED #(.width(1)) u_mux_156 (
        .y(_node_142),
        .sel(_node_141),
        .a(_T_87_8),
        .b(_node_140)
    );
    wire _node_143;
    EQ_UNSIGNED #(.width(6)) u_eq_157 (
        .y(_node_143),
        .a(6'd9),
        .b(_T_172)
    );
    wire _node_144;
    MUX_UNSIGNED #(.width(1)) u_mux_158 (
        .y(_node_144),
        .sel(_node_143),
        .a(_T_87_9),
        .b(_node_142)
    );
    wire _node_145;
    EQ_UNSIGNED #(.width(6)) u_eq_159 (
        .y(_node_145),
        .a(6'd10),
        .b(_T_172)
    );
    wire _node_146;
    MUX_UNSIGNED #(.width(1)) u_mux_160 (
        .y(_node_146),
        .sel(_node_145),
        .a(_T_87_10),
        .b(_node_144)
    );
    wire _node_147;
    EQ_UNSIGNED #(.width(6)) u_eq_161 (
        .y(_node_147),
        .a(6'd11),
        .b(_T_172)
    );
    wire _node_148;
    MUX_UNSIGNED #(.width(1)) u_mux_162 (
        .y(_node_148),
        .sel(_node_147),
        .a(_T_87_11),
        .b(_node_146)
    );
    wire _node_149;
    EQ_UNSIGNED #(.width(6)) u_eq_163 (
        .y(_node_149),
        .a(6'd12),
        .b(_T_172)
    );
    wire _node_150;
    MUX_UNSIGNED #(.width(1)) u_mux_164 (
        .y(_node_150),
        .sel(_node_149),
        .a(_T_87_12),
        .b(_node_148)
    );
    wire _node_151;
    EQ_UNSIGNED #(.width(6)) u_eq_165 (
        .y(_node_151),
        .a(6'd13),
        .b(_T_172)
    );
    wire _node_152;
    MUX_UNSIGNED #(.width(1)) u_mux_166 (
        .y(_node_152),
        .sel(_node_151),
        .a(_T_87_13),
        .b(_node_150)
    );
    wire _node_153;
    EQ_UNSIGNED #(.width(6)) u_eq_167 (
        .y(_node_153),
        .a(6'd14),
        .b(_T_172)
    );
    wire _node_154;
    MUX_UNSIGNED #(.width(1)) u_mux_168 (
        .y(_node_154),
        .sel(_node_153),
        .a(_T_87_14),
        .b(_node_152)
    );
    wire _node_155;
    EQ_UNSIGNED #(.width(6)) u_eq_169 (
        .y(_node_155),
        .a(6'd15),
        .b(_T_172)
    );
    wire _node_156;
    MUX_UNSIGNED #(.width(1)) u_mux_170 (
        .y(_node_156),
        .sel(_node_155),
        .a(_T_87_15),
        .b(_node_154)
    );
    wire _node_157;
    EQ_UNSIGNED #(.width(6)) u_eq_171 (
        .y(_node_157),
        .a(6'd16),
        .b(_T_172)
    );
    wire _node_158;
    MUX_UNSIGNED #(.width(1)) u_mux_172 (
        .y(_node_158),
        .sel(_node_157),
        .a(_T_87_16),
        .b(_node_156)
    );
    wire _node_159;
    EQ_UNSIGNED #(.width(6)) u_eq_173 (
        .y(_node_159),
        .a(6'd17),
        .b(_T_172)
    );
    wire _node_160;
    MUX_UNSIGNED #(.width(1)) u_mux_174 (
        .y(_node_160),
        .sel(_node_159),
        .a(_T_87_17),
        .b(_node_158)
    );
    wire _node_161;
    EQ_UNSIGNED #(.width(6)) u_eq_175 (
        .y(_node_161),
        .a(6'd18),
        .b(_T_172)
    );
    wire _node_162;
    MUX_UNSIGNED #(.width(1)) u_mux_176 (
        .y(_node_162),
        .sel(_node_161),
        .a(_T_87_18),
        .b(_node_160)
    );
    wire _node_163;
    EQ_UNSIGNED #(.width(6)) u_eq_177 (
        .y(_node_163),
        .a(6'd19),
        .b(_T_172)
    );
    wire _node_164;
    MUX_UNSIGNED #(.width(1)) u_mux_178 (
        .y(_node_164),
        .sel(_node_163),
        .a(_T_87_19),
        .b(_node_162)
    );
    wire _node_165;
    EQ_UNSIGNED #(.width(6)) u_eq_179 (
        .y(_node_165),
        .a(6'd20),
        .b(_T_172)
    );
    wire _node_166;
    MUX_UNSIGNED #(.width(1)) u_mux_180 (
        .y(_node_166),
        .sel(_node_165),
        .a(_T_87_20),
        .b(_node_164)
    );
    wire _node_167;
    EQ_UNSIGNED #(.width(6)) u_eq_181 (
        .y(_node_167),
        .a(6'd21),
        .b(_T_172)
    );
    wire _node_168;
    MUX_UNSIGNED #(.width(1)) u_mux_182 (
        .y(_node_168),
        .sel(_node_167),
        .a(_T_87_21),
        .b(_node_166)
    );
    wire _node_169;
    EQ_UNSIGNED #(.width(6)) u_eq_183 (
        .y(_node_169),
        .a(6'd22),
        .b(_T_172)
    );
    wire _node_170;
    MUX_UNSIGNED #(.width(1)) u_mux_184 (
        .y(_node_170),
        .sel(_node_169),
        .a(_T_87_22),
        .b(_node_168)
    );
    wire _node_171;
    EQ_UNSIGNED #(.width(6)) u_eq_185 (
        .y(_node_171),
        .a(6'd23),
        .b(_T_172)
    );
    wire _node_172;
    MUX_UNSIGNED #(.width(1)) u_mux_186 (
        .y(_node_172),
        .sel(_node_171),
        .a(_T_87_23),
        .b(_node_170)
    );
    wire _node_173;
    EQ_UNSIGNED #(.width(6)) u_eq_187 (
        .y(_node_173),
        .a(6'd24),
        .b(_T_172)
    );
    wire _node_174;
    MUX_UNSIGNED #(.width(1)) u_mux_188 (
        .y(_node_174),
        .sel(_node_173),
        .a(_T_87_24),
        .b(_node_172)
    );
    wire _node_175;
    EQ_UNSIGNED #(.width(6)) u_eq_189 (
        .y(_node_175),
        .a(6'd25),
        .b(_T_172)
    );
    wire _node_176;
    MUX_UNSIGNED #(.width(1)) u_mux_190 (
        .y(_node_176),
        .sel(_node_175),
        .a(_T_87_25),
        .b(_node_174)
    );
    wire _node_177;
    EQ_UNSIGNED #(.width(6)) u_eq_191 (
        .y(_node_177),
        .a(6'd26),
        .b(_T_172)
    );
    wire _node_178;
    MUX_UNSIGNED #(.width(1)) u_mux_192 (
        .y(_node_178),
        .sel(_node_177),
        .a(_T_87_26),
        .b(_node_176)
    );
    wire _node_179;
    EQ_UNSIGNED #(.width(6)) u_eq_193 (
        .y(_node_179),
        .a(6'd27),
        .b(_T_172)
    );
    wire _node_180;
    MUX_UNSIGNED #(.width(1)) u_mux_194 (
        .y(_node_180),
        .sel(_node_179),
        .a(_T_87_27),
        .b(_node_178)
    );
    wire _node_181;
    EQ_UNSIGNED #(.width(6)) u_eq_195 (
        .y(_node_181),
        .a(6'd28),
        .b(_T_172)
    );
    wire _node_182;
    MUX_UNSIGNED #(.width(1)) u_mux_196 (
        .y(_node_182),
        .sel(_node_181),
        .a(_T_87_28),
        .b(_node_180)
    );
    wire _node_183;
    EQ_UNSIGNED #(.width(6)) u_eq_197 (
        .y(_node_183),
        .a(6'd29),
        .b(_T_172)
    );
    wire _node_184;
    MUX_UNSIGNED #(.width(1)) u_mux_198 (
        .y(_node_184),
        .sel(_node_183),
        .a(_T_87_29),
        .b(_node_182)
    );
    wire _node_185;
    EQ_UNSIGNED #(.width(6)) u_eq_199 (
        .y(_node_185),
        .a(6'd30),
        .b(_T_172)
    );
    wire _node_186;
    MUX_UNSIGNED #(.width(1)) u_mux_200 (
        .y(_node_186),
        .sel(_node_185),
        .a(_T_87_30),
        .b(_node_184)
    );
    wire _node_187;
    EQ_UNSIGNED #(.width(6)) u_eq_201 (
        .y(_node_187),
        .a(6'd31),
        .b(_T_172)
    );
    wire _node_188;
    MUX_UNSIGNED #(.width(1)) u_mux_202 (
        .y(_node_188),
        .sel(_node_187),
        .a(_T_87_31),
        .b(_node_186)
    );
    wire _node_189;
    EQ_UNSIGNED #(.width(6)) u_eq_203 (
        .y(_node_189),
        .a(6'd32),
        .b(_T_172)
    );
    wire _node_190;
    MUX_UNSIGNED #(.width(1)) u_mux_204 (
        .y(_node_190),
        .sel(_node_189),
        .a(_T_87_32),
        .b(_node_188)
    );
    wire _node_191;
    EQ_UNSIGNED #(.width(6)) u_eq_205 (
        .y(_node_191),
        .a(6'd33),
        .b(_T_172)
    );
    wire _node_192;
    MUX_UNSIGNED #(.width(1)) u_mux_206 (
        .y(_node_192),
        .sel(_node_191),
        .a(_T_87_33),
        .b(_node_190)
    );
    wire _node_193;
    EQ_UNSIGNED #(.width(6)) u_eq_207 (
        .y(_node_193),
        .a(6'd34),
        .b(_T_172)
    );
    wire _node_194;
    MUX_UNSIGNED #(.width(1)) u_mux_208 (
        .y(_node_194),
        .sel(_node_193),
        .a(_T_87_34),
        .b(_node_192)
    );
    wire _node_195;
    EQ_UNSIGNED #(.width(6)) u_eq_209 (
        .y(_node_195),
        .a(6'd35),
        .b(_T_172)
    );
    wire _node_196;
    MUX_UNSIGNED #(.width(1)) u_mux_210 (
        .y(_node_196),
        .sel(_node_195),
        .a(_T_87_35),
        .b(_node_194)
    );
    wire _node_197;
    EQ_UNSIGNED #(.width(6)) u_eq_211 (
        .y(_node_197),
        .a(6'd36),
        .b(_T_172)
    );
    wire _node_198;
    MUX_UNSIGNED #(.width(1)) u_mux_212 (
        .y(_node_198),
        .sel(_node_197),
        .a(_T_87_36),
        .b(_node_196)
    );
    wire _node_199;
    EQ_UNSIGNED #(.width(6)) u_eq_213 (
        .y(_node_199),
        .a(6'd37),
        .b(_T_172)
    );
    wire _node_200;
    MUX_UNSIGNED #(.width(1)) u_mux_214 (
        .y(_node_200),
        .sel(_node_199),
        .a(_T_87_37),
        .b(_node_198)
    );
    wire _node_201;
    EQ_UNSIGNED #(.width(6)) u_eq_215 (
        .y(_node_201),
        .a(6'd38),
        .b(_T_172)
    );
    wire _node_202;
    MUX_UNSIGNED #(.width(1)) u_mux_216 (
        .y(_node_202),
        .sel(_node_201),
        .a(_T_87_38),
        .b(_node_200)
    );
    wire _node_203;
    EQ_UNSIGNED #(.width(6)) u_eq_217 (
        .y(_node_203),
        .a(6'd39),
        .b(_T_172)
    );
    wire _node_204;
    MUX_UNSIGNED #(.width(1)) u_mux_218 (
        .y(_node_204),
        .sel(_node_203),
        .a(_T_87_39),
        .b(_node_202)
    );
    wire _node_205;
    EQ_UNSIGNED #(.width(6)) u_eq_219 (
        .y(_node_205),
        .a(6'd40),
        .b(_T_172)
    );
    wire _node_206;
    MUX_UNSIGNED #(.width(1)) u_mux_220 (
        .y(_node_206),
        .sel(_node_205),
        .a(_T_87_40),
        .b(_node_204)
    );
    wire _node_207;
    EQ_UNSIGNED #(.width(6)) u_eq_221 (
        .y(_node_207),
        .a(6'd41),
        .b(_T_172)
    );
    wire _node_208;
    MUX_UNSIGNED #(.width(1)) u_mux_222 (
        .y(_node_208),
        .sel(_node_207),
        .a(_T_87_41),
        .b(_node_206)
    );
    wire _node_209;
    EQ_UNSIGNED #(.width(6)) u_eq_223 (
        .y(_node_209),
        .a(6'd42),
        .b(_T_172)
    );
    wire _node_210;
    MUX_UNSIGNED #(.width(1)) u_mux_224 (
        .y(_node_210),
        .sel(_node_209),
        .a(_T_87_42),
        .b(_node_208)
    );
    wire _node_211;
    EQ_UNSIGNED #(.width(6)) u_eq_225 (
        .y(_node_211),
        .a(6'd43),
        .b(_T_172)
    );
    wire _node_212;
    MUX_UNSIGNED #(.width(1)) u_mux_226 (
        .y(_node_212),
        .sel(_node_211),
        .a(_T_87_43),
        .b(_node_210)
    );
    wire _node_213;
    EQ_UNSIGNED #(.width(6)) u_eq_227 (
        .y(_node_213),
        .a(6'd44),
        .b(_T_172)
    );
    wire _node_214;
    MUX_UNSIGNED #(.width(1)) u_mux_228 (
        .y(_node_214),
        .sel(_node_213),
        .a(_T_87_44),
        .b(_node_212)
    );
    wire _node_215;
    EQ_UNSIGNED #(.width(6)) u_eq_229 (
        .y(_node_215),
        .a(6'd45),
        .b(_T_172)
    );
    wire _node_216;
    MUX_UNSIGNED #(.width(1)) u_mux_230 (
        .y(_node_216),
        .sel(_node_215),
        .a(_T_87_45),
        .b(_node_214)
    );
    wire _node_217;
    EQ_UNSIGNED #(.width(6)) u_eq_231 (
        .y(_node_217),
        .a(6'd46),
        .b(_T_172)
    );
    wire _node_218;
    MUX_UNSIGNED #(.width(1)) u_mux_232 (
        .y(_node_218),
        .sel(_node_217),
        .a(_T_87_46),
        .b(_node_216)
    );
    wire _node_219;
    EQ_UNSIGNED #(.width(6)) u_eq_233 (
        .y(_node_219),
        .a(6'd47),
        .b(_T_172)
    );
    wire _node_220;
    MUX_UNSIGNED #(.width(1)) u_mux_234 (
        .y(_node_220),
        .sel(_node_219),
        .a(_T_87_47),
        .b(_node_218)
    );
    wire _node_221;
    EQ_UNSIGNED #(.width(6)) u_eq_235 (
        .y(_node_221),
        .a(6'd48),
        .b(_T_172)
    );
    wire _node_222;
    MUX_UNSIGNED #(.width(1)) u_mux_236 (
        .y(_node_222),
        .sel(_node_221),
        .a(_T_87_48),
        .b(_node_220)
    );
    wire _node_223;
    EQ_UNSIGNED #(.width(6)) u_eq_237 (
        .y(_node_223),
        .a(6'd49),
        .b(_T_172)
    );
    wire _node_224;
    MUX_UNSIGNED #(.width(1)) u_mux_238 (
        .y(_node_224),
        .sel(_node_223),
        .a(_T_87_49),
        .b(_node_222)
    );
    wire _node_225;
    EQ_UNSIGNED #(.width(6)) u_eq_239 (
        .y(_node_225),
        .a(6'd50),
        .b(_T_172)
    );
    wire _node_226;
    MUX_UNSIGNED #(.width(1)) u_mux_240 (
        .y(_node_226),
        .sel(_node_225),
        .a(_T_87_50),
        .b(_node_224)
    );
    wire _node_227;
    EQ_UNSIGNED #(.width(6)) u_eq_241 (
        .y(_node_227),
        .a(6'd51),
        .b(_T_172)
    );
    wire _node_228;
    MUX_UNSIGNED #(.width(1)) u_mux_242 (
        .y(_node_228),
        .sel(_node_227),
        .a(_T_87_51),
        .b(_node_226)
    );
    wire _node_229;
    EQ_UNSIGNED #(.width(6)) u_eq_243 (
        .y(_node_229),
        .a(6'd52),
        .b(_T_172)
    );
    wire _node_230;
    MUX_UNSIGNED #(.width(1)) u_mux_244 (
        .y(_node_230),
        .sel(_node_229),
        .a(_T_87_52),
        .b(_node_228)
    );
    wire _T_173;
    BITWISEAND #(.width(1)) bitwiseand_245 (
        .y(_T_173),
        .a(_c__io_read_routing_table_request_valid),
        .b(_c__io_read_routing_table_request_ready)
    );
    wire _T_175;
    EQ_UNSIGNED #(.width(4)) u_eq_246 (
        .y(_T_175),
        .a(_value__q),
        .b(4'h8)
    );
    wire [4:0] _T_177;
    wire [3:0] _WTEMP_11;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_247 (
        .y(_WTEMP_11),
        .in(1'h1)
    );
    ADD_UNSIGNED #(.width(4)) u_add_248 (
        .y(_T_177),
        .a(_value__q),
        .b(_WTEMP_11)
    );
    wire [3:0] _T_178;
    TAIL #(.width(5), .n(1)) tail_249 (
        .y(_T_178),
        .in(_T_177)
    );
    wire _T_181;
    EQ_UNSIGNED #(.width(1)) u_eq_250 (
        .y(_T_181),
        .a(__T_7__q),
        .b(1'h0)
    );
    wire _T_183;
    wire [7:0] _WTEMP_12;
    PAD_UNSIGNED #(.width(6), .n(8)) u_pad_251 (
        .y(_WTEMP_12),
        .in(6'h33)
    );
    EQ_UNSIGNED #(.width(8)) u_eq_252 (
        .y(_T_183),
        .a(__T_4__q),
        .b(_WTEMP_12)
    );
    wire [8:0] _T_186;
    wire [7:0] _WTEMP_13;
    PAD_UNSIGNED #(.width(1), .n(8)) u_pad_253 (
        .y(_WTEMP_13),
        .in(1'h1)
    );
    ADD_UNSIGNED #(.width(8)) u_add_254 (
        .y(_T_186),
        .a(__T_4__q),
        .b(_WTEMP_13)
    );
    wire [7:0] _T_187;
    TAIL #(.width(9), .n(1)) tail_255 (
        .y(_T_187),
        .in(_T_186)
    );
    wire _node_231;
    MUX_UNSIGNED #(.width(1)) u_mux_256 (
        .y(_node_231),
        .sel(_T_183),
        .a(1'h1),
        .b(__T_7__q)
    );
    wire [7:0] _node_232;
    MUX_UNSIGNED #(.width(8)) u_mux_257 (
        .y(_node_232),
        .sel(_T_181),
        .a(_T_187),
        .b(__T_4__q)
    );
    wire _node_233;
    MUX_UNSIGNED #(.width(1)) u_mux_258 (
        .y(_node_233),
        .sel(_T_181),
        .a(_node_231),
        .b(__T_7__q)
    );
    wire [3:0] _node_234;
    wire [3:0] _WTEMP_14;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_259 (
        .y(_WTEMP_14),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(4)) u_mux_260 (
        .y(_node_234),
        .sel(_T_175),
        .a(_WTEMP_14),
        .b(_T_178)
    );
    wire _T_243_0;
    wire _T_243_1;
    wire _T_243_2;
    wire _T_243_3;
    wire _T_243_4;
    wire _T_243_5;
    wire _T_243_6;
    wire _T_243_7;
    wire _T_243_8;
    wire _T_243_9;
    wire _T_243_10;
    wire _T_243_11;
    wire _T_243_12;
    wire _T_243_13;
    wire _T_243_14;
    wire _T_243_15;
    wire _T_243_16;
    wire _T_243_17;
    wire _T_243_18;
    wire _T_243_19;
    wire _T_243_20;
    wire _T_243_21;
    wire _T_243_22;
    wire _T_243_23;
    wire _T_243_24;
    wire _T_243_25;
    wire _T_243_26;
    wire _T_243_27;
    wire _T_243_28;
    wire _T_243_29;
    wire _T_243_30;
    wire _T_243_31;
    wire _T_243_32;
    wire _T_243_33;
    wire _T_243_34;
    wire _T_243_35;
    wire _T_243_36;
    wire _T_243_37;
    wire _T_243_38;
    wire _T_243_39;
    wire _T_243_40;
    wire _T_243_41;
    wire _T_243_42;
    wire _T_243_43;
    wire _T_243_44;
    wire _T_243_45;
    wire _T_243_46;
    wire _T_243_47;
    wire _T_243_48;
    wire _T_243_49;
    wire _T_243_50;
    wire _T_243_51;
    wire _T_243_52;
    wire [4:0] _value_1__q;
    wire [4:0] _value_1__d;
    DFF_POSCLK #(.width(5)) value_1 (
        .q(_value_1__q),
        .d(_value_1__d),
        .clk(clock)
    );
    wire [4:0] _WTEMP_15;
    MUX_UNSIGNED #(.width(5)) u_mux_261 (
        .y(_value_1__d),
        .sel(reset),
        .a(5'h0),
        .b(_WTEMP_15)
    );
    wire [3:0] _T_328_0;
    wire [3:0] _T_328_1;
    wire [3:0] _T_328_2;
    wire [3:0] _T_328_3;
    wire [3:0] _T_328_4;
    wire [3:0] _T_328_5;
    wire [3:0] _T_328_6;
    wire [3:0] _T_328_7;
    wire [3:0] _T_328_8;
    wire [3:0] _T_328_9;
    wire [3:0] _T_328_10;
    wire [3:0] _T_328_11;
    wire [3:0] _T_328_12;
    wire [3:0] _T_328_13;
    wire [3:0] _T_328_14;
    wire [3:0] _T_328_15;
    wire [3:0] _T_328_16;
    wire [3:0] _T_328_17;
    wire [3:0] _T_328_18;
    wire [3:0] _T_328_19;
    wire [3:0] _T_328_20;
    wire [3:0] _T_328_21;
    wire [3:0] _T_328_22;
    wire [3:0] _T_328_23;
    wire [3:0] _T_328_24;
    wire [30:0] _T_383_0;
    wire [30:0] _T_383_1;
    wire [30:0] _T_383_2;
    wire [30:0] _T_383_3;
    wire [30:0] _T_383_4;
    wire [30:0] _T_383_5;
    wire [30:0] _T_383_6;
    wire [30:0] _T_383_7;
    wire [30:0] _T_383_8;
    wire [30:0] _T_383_9;
    wire [30:0] _T_383_10;
    wire [30:0] _T_383_11;
    wire [30:0] _T_383_12;
    wire [30:0] _T_383_13;
    wire [30:0] _T_383_14;
    wire [30:0] _T_383_15;
    wire [30:0] _T_383_16;
    wire [30:0] _T_383_17;
    wire [30:0] _T_383_18;
    wire [30:0] _T_383_19;
    wire [30:0] _T_383_20;
    wire [30:0] _T_383_21;
    wire [30:0] _T_383_22;
    wire [30:0] _T_383_23;
    wire [30:0] _T_383_24;
    wire _node_235;
    EQ_UNSIGNED #(.width(5)) u_eq_262 (
        .y(_node_235),
        .a(5'd0),
        .b(_value_1__q)
    );
    wire [3:0] _node_236;
    assign _node_236 = _T_328_0;
    wire _node_237;
    EQ_UNSIGNED #(.width(5)) u_eq_263 (
        .y(_node_237),
        .a(5'd1),
        .b(_value_1__q)
    );
    wire [3:0] _node_238;
    MUX_UNSIGNED #(.width(4)) u_mux_264 (
        .y(_node_238),
        .sel(_node_237),
        .a(_T_328_1),
        .b(_node_236)
    );
    wire _node_239;
    EQ_UNSIGNED #(.width(5)) u_eq_265 (
        .y(_node_239),
        .a(5'd2),
        .b(_value_1__q)
    );
    wire [3:0] _node_240;
    MUX_UNSIGNED #(.width(4)) u_mux_266 (
        .y(_node_240),
        .sel(_node_239),
        .a(_T_328_2),
        .b(_node_238)
    );
    wire _node_241;
    EQ_UNSIGNED #(.width(5)) u_eq_267 (
        .y(_node_241),
        .a(5'd3),
        .b(_value_1__q)
    );
    wire [3:0] _node_242;
    MUX_UNSIGNED #(.width(4)) u_mux_268 (
        .y(_node_242),
        .sel(_node_241),
        .a(_T_328_3),
        .b(_node_240)
    );
    wire _node_243;
    EQ_UNSIGNED #(.width(5)) u_eq_269 (
        .y(_node_243),
        .a(5'd4),
        .b(_value_1__q)
    );
    wire [3:0] _node_244;
    MUX_UNSIGNED #(.width(4)) u_mux_270 (
        .y(_node_244),
        .sel(_node_243),
        .a(_T_328_4),
        .b(_node_242)
    );
    wire _node_245;
    EQ_UNSIGNED #(.width(5)) u_eq_271 (
        .y(_node_245),
        .a(5'd5),
        .b(_value_1__q)
    );
    wire [3:0] _node_246;
    MUX_UNSIGNED #(.width(4)) u_mux_272 (
        .y(_node_246),
        .sel(_node_245),
        .a(_T_328_5),
        .b(_node_244)
    );
    wire _node_247;
    EQ_UNSIGNED #(.width(5)) u_eq_273 (
        .y(_node_247),
        .a(5'd6),
        .b(_value_1__q)
    );
    wire [3:0] _node_248;
    MUX_UNSIGNED #(.width(4)) u_mux_274 (
        .y(_node_248),
        .sel(_node_247),
        .a(_T_328_6),
        .b(_node_246)
    );
    wire _node_249;
    EQ_UNSIGNED #(.width(5)) u_eq_275 (
        .y(_node_249),
        .a(5'd7),
        .b(_value_1__q)
    );
    wire [3:0] _node_250;
    MUX_UNSIGNED #(.width(4)) u_mux_276 (
        .y(_node_250),
        .sel(_node_249),
        .a(_T_328_7),
        .b(_node_248)
    );
    wire _node_251;
    EQ_UNSIGNED #(.width(5)) u_eq_277 (
        .y(_node_251),
        .a(5'd8),
        .b(_value_1__q)
    );
    wire [3:0] _node_252;
    MUX_UNSIGNED #(.width(4)) u_mux_278 (
        .y(_node_252),
        .sel(_node_251),
        .a(_T_328_8),
        .b(_node_250)
    );
    wire _node_253;
    EQ_UNSIGNED #(.width(5)) u_eq_279 (
        .y(_node_253),
        .a(5'd9),
        .b(_value_1__q)
    );
    wire [3:0] _node_254;
    MUX_UNSIGNED #(.width(4)) u_mux_280 (
        .y(_node_254),
        .sel(_node_253),
        .a(_T_328_9),
        .b(_node_252)
    );
    wire _node_255;
    EQ_UNSIGNED #(.width(5)) u_eq_281 (
        .y(_node_255),
        .a(5'd10),
        .b(_value_1__q)
    );
    wire [3:0] _node_256;
    MUX_UNSIGNED #(.width(4)) u_mux_282 (
        .y(_node_256),
        .sel(_node_255),
        .a(_T_328_10),
        .b(_node_254)
    );
    wire _node_257;
    EQ_UNSIGNED #(.width(5)) u_eq_283 (
        .y(_node_257),
        .a(5'd11),
        .b(_value_1__q)
    );
    wire [3:0] _node_258;
    MUX_UNSIGNED #(.width(4)) u_mux_284 (
        .y(_node_258),
        .sel(_node_257),
        .a(_T_328_11),
        .b(_node_256)
    );
    wire _node_259;
    EQ_UNSIGNED #(.width(5)) u_eq_285 (
        .y(_node_259),
        .a(5'd12),
        .b(_value_1__q)
    );
    wire [3:0] _node_260;
    MUX_UNSIGNED #(.width(4)) u_mux_286 (
        .y(_node_260),
        .sel(_node_259),
        .a(_T_328_12),
        .b(_node_258)
    );
    wire _node_261;
    EQ_UNSIGNED #(.width(5)) u_eq_287 (
        .y(_node_261),
        .a(5'd13),
        .b(_value_1__q)
    );
    wire [3:0] _node_262;
    MUX_UNSIGNED #(.width(4)) u_mux_288 (
        .y(_node_262),
        .sel(_node_261),
        .a(_T_328_13),
        .b(_node_260)
    );
    wire _node_263;
    EQ_UNSIGNED #(.width(5)) u_eq_289 (
        .y(_node_263),
        .a(5'd14),
        .b(_value_1__q)
    );
    wire [3:0] _node_264;
    MUX_UNSIGNED #(.width(4)) u_mux_290 (
        .y(_node_264),
        .sel(_node_263),
        .a(_T_328_14),
        .b(_node_262)
    );
    wire _node_265;
    EQ_UNSIGNED #(.width(5)) u_eq_291 (
        .y(_node_265),
        .a(5'd15),
        .b(_value_1__q)
    );
    wire [3:0] _node_266;
    MUX_UNSIGNED #(.width(4)) u_mux_292 (
        .y(_node_266),
        .sel(_node_265),
        .a(_T_328_15),
        .b(_node_264)
    );
    wire _node_267;
    EQ_UNSIGNED #(.width(5)) u_eq_293 (
        .y(_node_267),
        .a(5'd16),
        .b(_value_1__q)
    );
    wire [3:0] _node_268;
    MUX_UNSIGNED #(.width(4)) u_mux_294 (
        .y(_node_268),
        .sel(_node_267),
        .a(_T_328_16),
        .b(_node_266)
    );
    wire _node_269;
    EQ_UNSIGNED #(.width(5)) u_eq_295 (
        .y(_node_269),
        .a(5'd17),
        .b(_value_1__q)
    );
    wire [3:0] _node_270;
    MUX_UNSIGNED #(.width(4)) u_mux_296 (
        .y(_node_270),
        .sel(_node_269),
        .a(_T_328_17),
        .b(_node_268)
    );
    wire _node_271;
    EQ_UNSIGNED #(.width(5)) u_eq_297 (
        .y(_node_271),
        .a(5'd18),
        .b(_value_1__q)
    );
    wire [3:0] _node_272;
    MUX_UNSIGNED #(.width(4)) u_mux_298 (
        .y(_node_272),
        .sel(_node_271),
        .a(_T_328_18),
        .b(_node_270)
    );
    wire _node_273;
    EQ_UNSIGNED #(.width(5)) u_eq_299 (
        .y(_node_273),
        .a(5'd19),
        .b(_value_1__q)
    );
    wire [3:0] _node_274;
    MUX_UNSIGNED #(.width(4)) u_mux_300 (
        .y(_node_274),
        .sel(_node_273),
        .a(_T_328_19),
        .b(_node_272)
    );
    wire _node_275;
    EQ_UNSIGNED #(.width(5)) u_eq_301 (
        .y(_node_275),
        .a(5'd20),
        .b(_value_1__q)
    );
    wire [3:0] _node_276;
    MUX_UNSIGNED #(.width(4)) u_mux_302 (
        .y(_node_276),
        .sel(_node_275),
        .a(_T_328_20),
        .b(_node_274)
    );
    wire _node_277;
    EQ_UNSIGNED #(.width(5)) u_eq_303 (
        .y(_node_277),
        .a(5'd21),
        .b(_value_1__q)
    );
    wire [3:0] _node_278;
    MUX_UNSIGNED #(.width(4)) u_mux_304 (
        .y(_node_278),
        .sel(_node_277),
        .a(_T_328_21),
        .b(_node_276)
    );
    wire _node_279;
    EQ_UNSIGNED #(.width(5)) u_eq_305 (
        .y(_node_279),
        .a(5'd22),
        .b(_value_1__q)
    );
    wire [3:0] _node_280;
    MUX_UNSIGNED #(.width(4)) u_mux_306 (
        .y(_node_280),
        .sel(_node_279),
        .a(_T_328_22),
        .b(_node_278)
    );
    wire _node_281;
    EQ_UNSIGNED #(.width(5)) u_eq_307 (
        .y(_node_281),
        .a(5'd23),
        .b(_value_1__q)
    );
    wire [3:0] _node_282;
    MUX_UNSIGNED #(.width(4)) u_mux_308 (
        .y(_node_282),
        .sel(_node_281),
        .a(_T_328_23),
        .b(_node_280)
    );
    wire _node_283;
    EQ_UNSIGNED #(.width(5)) u_eq_309 (
        .y(_node_283),
        .a(5'd24),
        .b(_value_1__q)
    );
    wire [3:0] _node_284;
    MUX_UNSIGNED #(.width(4)) u_mux_310 (
        .y(_node_284),
        .sel(_node_283),
        .a(_T_328_24),
        .b(_node_282)
    );
    wire _node_285;
    EQ_UNSIGNED #(.width(5)) u_eq_311 (
        .y(_node_285),
        .a(5'd0),
        .b(_value_1__q)
    );
    wire [30:0] _node_286;
    assign _node_286 = _T_383_0;
    wire _node_287;
    EQ_UNSIGNED #(.width(5)) u_eq_312 (
        .y(_node_287),
        .a(5'd1),
        .b(_value_1__q)
    );
    wire [30:0] _node_288;
    MUX_UNSIGNED #(.width(31)) u_mux_313 (
        .y(_node_288),
        .sel(_node_287),
        .a(_T_383_1),
        .b(_node_286)
    );
    wire _node_289;
    EQ_UNSIGNED #(.width(5)) u_eq_314 (
        .y(_node_289),
        .a(5'd2),
        .b(_value_1__q)
    );
    wire [30:0] _node_290;
    MUX_UNSIGNED #(.width(31)) u_mux_315 (
        .y(_node_290),
        .sel(_node_289),
        .a(_T_383_2),
        .b(_node_288)
    );
    wire _node_291;
    EQ_UNSIGNED #(.width(5)) u_eq_316 (
        .y(_node_291),
        .a(5'd3),
        .b(_value_1__q)
    );
    wire [30:0] _node_292;
    MUX_UNSIGNED #(.width(31)) u_mux_317 (
        .y(_node_292),
        .sel(_node_291),
        .a(_T_383_3),
        .b(_node_290)
    );
    wire _node_293;
    EQ_UNSIGNED #(.width(5)) u_eq_318 (
        .y(_node_293),
        .a(5'd4),
        .b(_value_1__q)
    );
    wire [30:0] _node_294;
    MUX_UNSIGNED #(.width(31)) u_mux_319 (
        .y(_node_294),
        .sel(_node_293),
        .a(_T_383_4),
        .b(_node_292)
    );
    wire _node_295;
    EQ_UNSIGNED #(.width(5)) u_eq_320 (
        .y(_node_295),
        .a(5'd5),
        .b(_value_1__q)
    );
    wire [30:0] _node_296;
    MUX_UNSIGNED #(.width(31)) u_mux_321 (
        .y(_node_296),
        .sel(_node_295),
        .a(_T_383_5),
        .b(_node_294)
    );
    wire _node_297;
    EQ_UNSIGNED #(.width(5)) u_eq_322 (
        .y(_node_297),
        .a(5'd6),
        .b(_value_1__q)
    );
    wire [30:0] _node_298;
    MUX_UNSIGNED #(.width(31)) u_mux_323 (
        .y(_node_298),
        .sel(_node_297),
        .a(_T_383_6),
        .b(_node_296)
    );
    wire _node_299;
    EQ_UNSIGNED #(.width(5)) u_eq_324 (
        .y(_node_299),
        .a(5'd7),
        .b(_value_1__q)
    );
    wire [30:0] _node_300;
    MUX_UNSIGNED #(.width(31)) u_mux_325 (
        .y(_node_300),
        .sel(_node_299),
        .a(_T_383_7),
        .b(_node_298)
    );
    wire _node_301;
    EQ_UNSIGNED #(.width(5)) u_eq_326 (
        .y(_node_301),
        .a(5'd8),
        .b(_value_1__q)
    );
    wire [30:0] _node_302;
    MUX_UNSIGNED #(.width(31)) u_mux_327 (
        .y(_node_302),
        .sel(_node_301),
        .a(_T_383_8),
        .b(_node_300)
    );
    wire _node_303;
    EQ_UNSIGNED #(.width(5)) u_eq_328 (
        .y(_node_303),
        .a(5'd9),
        .b(_value_1__q)
    );
    wire [30:0] _node_304;
    MUX_UNSIGNED #(.width(31)) u_mux_329 (
        .y(_node_304),
        .sel(_node_303),
        .a(_T_383_9),
        .b(_node_302)
    );
    wire _node_305;
    EQ_UNSIGNED #(.width(5)) u_eq_330 (
        .y(_node_305),
        .a(5'd10),
        .b(_value_1__q)
    );
    wire [30:0] _node_306;
    MUX_UNSIGNED #(.width(31)) u_mux_331 (
        .y(_node_306),
        .sel(_node_305),
        .a(_T_383_10),
        .b(_node_304)
    );
    wire _node_307;
    EQ_UNSIGNED #(.width(5)) u_eq_332 (
        .y(_node_307),
        .a(5'd11),
        .b(_value_1__q)
    );
    wire [30:0] _node_308;
    MUX_UNSIGNED #(.width(31)) u_mux_333 (
        .y(_node_308),
        .sel(_node_307),
        .a(_T_383_11),
        .b(_node_306)
    );
    wire _node_309;
    EQ_UNSIGNED #(.width(5)) u_eq_334 (
        .y(_node_309),
        .a(5'd12),
        .b(_value_1__q)
    );
    wire [30:0] _node_310;
    MUX_UNSIGNED #(.width(31)) u_mux_335 (
        .y(_node_310),
        .sel(_node_309),
        .a(_T_383_12),
        .b(_node_308)
    );
    wire _node_311;
    EQ_UNSIGNED #(.width(5)) u_eq_336 (
        .y(_node_311),
        .a(5'd13),
        .b(_value_1__q)
    );
    wire [30:0] _node_312;
    MUX_UNSIGNED #(.width(31)) u_mux_337 (
        .y(_node_312),
        .sel(_node_311),
        .a(_T_383_13),
        .b(_node_310)
    );
    wire _node_313;
    EQ_UNSIGNED #(.width(5)) u_eq_338 (
        .y(_node_313),
        .a(5'd14),
        .b(_value_1__q)
    );
    wire [30:0] _node_314;
    MUX_UNSIGNED #(.width(31)) u_mux_339 (
        .y(_node_314),
        .sel(_node_313),
        .a(_T_383_14),
        .b(_node_312)
    );
    wire _node_315;
    EQ_UNSIGNED #(.width(5)) u_eq_340 (
        .y(_node_315),
        .a(5'd15),
        .b(_value_1__q)
    );
    wire [30:0] _node_316;
    MUX_UNSIGNED #(.width(31)) u_mux_341 (
        .y(_node_316),
        .sel(_node_315),
        .a(_T_383_15),
        .b(_node_314)
    );
    wire _node_317;
    EQ_UNSIGNED #(.width(5)) u_eq_342 (
        .y(_node_317),
        .a(5'd16),
        .b(_value_1__q)
    );
    wire [30:0] _node_318;
    MUX_UNSIGNED #(.width(31)) u_mux_343 (
        .y(_node_318),
        .sel(_node_317),
        .a(_T_383_16),
        .b(_node_316)
    );
    wire _node_319;
    EQ_UNSIGNED #(.width(5)) u_eq_344 (
        .y(_node_319),
        .a(5'd17),
        .b(_value_1__q)
    );
    wire [30:0] _node_320;
    MUX_UNSIGNED #(.width(31)) u_mux_345 (
        .y(_node_320),
        .sel(_node_319),
        .a(_T_383_17),
        .b(_node_318)
    );
    wire _node_321;
    EQ_UNSIGNED #(.width(5)) u_eq_346 (
        .y(_node_321),
        .a(5'd18),
        .b(_value_1__q)
    );
    wire [30:0] _node_322;
    MUX_UNSIGNED #(.width(31)) u_mux_347 (
        .y(_node_322),
        .sel(_node_321),
        .a(_T_383_18),
        .b(_node_320)
    );
    wire _node_323;
    EQ_UNSIGNED #(.width(5)) u_eq_348 (
        .y(_node_323),
        .a(5'd19),
        .b(_value_1__q)
    );
    wire [30:0] _node_324;
    MUX_UNSIGNED #(.width(31)) u_mux_349 (
        .y(_node_324),
        .sel(_node_323),
        .a(_T_383_19),
        .b(_node_322)
    );
    wire _node_325;
    EQ_UNSIGNED #(.width(5)) u_eq_350 (
        .y(_node_325),
        .a(5'd20),
        .b(_value_1__q)
    );
    wire [30:0] _node_326;
    MUX_UNSIGNED #(.width(31)) u_mux_351 (
        .y(_node_326),
        .sel(_node_325),
        .a(_T_383_20),
        .b(_node_324)
    );
    wire _node_327;
    EQ_UNSIGNED #(.width(5)) u_eq_352 (
        .y(_node_327),
        .a(5'd21),
        .b(_value_1__q)
    );
    wire [30:0] _node_328;
    MUX_UNSIGNED #(.width(31)) u_mux_353 (
        .y(_node_328),
        .sel(_node_327),
        .a(_T_383_21),
        .b(_node_326)
    );
    wire _node_329;
    EQ_UNSIGNED #(.width(5)) u_eq_354 (
        .y(_node_329),
        .a(5'd22),
        .b(_value_1__q)
    );
    wire [30:0] _node_330;
    MUX_UNSIGNED #(.width(31)) u_mux_355 (
        .y(_node_330),
        .sel(_node_329),
        .a(_T_383_22),
        .b(_node_328)
    );
    wire _node_331;
    EQ_UNSIGNED #(.width(5)) u_eq_356 (
        .y(_node_331),
        .a(5'd23),
        .b(_value_1__q)
    );
    wire [30:0] _node_332;
    MUX_UNSIGNED #(.width(31)) u_mux_357 (
        .y(_node_332),
        .sel(_node_331),
        .a(_T_383_23),
        .b(_node_330)
    );
    wire _node_333;
    EQ_UNSIGNED #(.width(5)) u_eq_358 (
        .y(_node_333),
        .a(5'd24),
        .b(_value_1__q)
    );
    wire [30:0] _node_334;
    MUX_UNSIGNED #(.width(31)) u_mux_359 (
        .y(_node_334),
        .sel(_node_333),
        .a(_T_383_24),
        .b(_node_332)
    );
    wire [5:0] _T_414;
    BITS #(.width(8), .high(5), .low(0)) bits_360 (
        .y(_T_414),
        .in(__T_4__q)
    );
    wire _node_335;
    EQ_UNSIGNED #(.width(6)) u_eq_361 (
        .y(_node_335),
        .a(6'd0),
        .b(_T_414)
    );
    wire _node_336;
    assign _node_336 = _T_243_0;
    wire _node_337;
    EQ_UNSIGNED #(.width(6)) u_eq_362 (
        .y(_node_337),
        .a(6'd1),
        .b(_T_414)
    );
    wire _node_338;
    MUX_UNSIGNED #(.width(1)) u_mux_363 (
        .y(_node_338),
        .sel(_node_337),
        .a(_T_243_1),
        .b(_node_336)
    );
    wire _node_339;
    EQ_UNSIGNED #(.width(6)) u_eq_364 (
        .y(_node_339),
        .a(6'd2),
        .b(_T_414)
    );
    wire _node_340;
    MUX_UNSIGNED #(.width(1)) u_mux_365 (
        .y(_node_340),
        .sel(_node_339),
        .a(_T_243_2),
        .b(_node_338)
    );
    wire _node_341;
    EQ_UNSIGNED #(.width(6)) u_eq_366 (
        .y(_node_341),
        .a(6'd3),
        .b(_T_414)
    );
    wire _node_342;
    MUX_UNSIGNED #(.width(1)) u_mux_367 (
        .y(_node_342),
        .sel(_node_341),
        .a(_T_243_3),
        .b(_node_340)
    );
    wire _node_343;
    EQ_UNSIGNED #(.width(6)) u_eq_368 (
        .y(_node_343),
        .a(6'd4),
        .b(_T_414)
    );
    wire _node_344;
    MUX_UNSIGNED #(.width(1)) u_mux_369 (
        .y(_node_344),
        .sel(_node_343),
        .a(_T_243_4),
        .b(_node_342)
    );
    wire _node_345;
    EQ_UNSIGNED #(.width(6)) u_eq_370 (
        .y(_node_345),
        .a(6'd5),
        .b(_T_414)
    );
    wire _node_346;
    MUX_UNSIGNED #(.width(1)) u_mux_371 (
        .y(_node_346),
        .sel(_node_345),
        .a(_T_243_5),
        .b(_node_344)
    );
    wire _node_347;
    EQ_UNSIGNED #(.width(6)) u_eq_372 (
        .y(_node_347),
        .a(6'd6),
        .b(_T_414)
    );
    wire _node_348;
    MUX_UNSIGNED #(.width(1)) u_mux_373 (
        .y(_node_348),
        .sel(_node_347),
        .a(_T_243_6),
        .b(_node_346)
    );
    wire _node_349;
    EQ_UNSIGNED #(.width(6)) u_eq_374 (
        .y(_node_349),
        .a(6'd7),
        .b(_T_414)
    );
    wire _node_350;
    MUX_UNSIGNED #(.width(1)) u_mux_375 (
        .y(_node_350),
        .sel(_node_349),
        .a(_T_243_7),
        .b(_node_348)
    );
    wire _node_351;
    EQ_UNSIGNED #(.width(6)) u_eq_376 (
        .y(_node_351),
        .a(6'd8),
        .b(_T_414)
    );
    wire _node_352;
    MUX_UNSIGNED #(.width(1)) u_mux_377 (
        .y(_node_352),
        .sel(_node_351),
        .a(_T_243_8),
        .b(_node_350)
    );
    wire _node_353;
    EQ_UNSIGNED #(.width(6)) u_eq_378 (
        .y(_node_353),
        .a(6'd9),
        .b(_T_414)
    );
    wire _node_354;
    MUX_UNSIGNED #(.width(1)) u_mux_379 (
        .y(_node_354),
        .sel(_node_353),
        .a(_T_243_9),
        .b(_node_352)
    );
    wire _node_355;
    EQ_UNSIGNED #(.width(6)) u_eq_380 (
        .y(_node_355),
        .a(6'd10),
        .b(_T_414)
    );
    wire _node_356;
    MUX_UNSIGNED #(.width(1)) u_mux_381 (
        .y(_node_356),
        .sel(_node_355),
        .a(_T_243_10),
        .b(_node_354)
    );
    wire _node_357;
    EQ_UNSIGNED #(.width(6)) u_eq_382 (
        .y(_node_357),
        .a(6'd11),
        .b(_T_414)
    );
    wire _node_358;
    MUX_UNSIGNED #(.width(1)) u_mux_383 (
        .y(_node_358),
        .sel(_node_357),
        .a(_T_243_11),
        .b(_node_356)
    );
    wire _node_359;
    EQ_UNSIGNED #(.width(6)) u_eq_384 (
        .y(_node_359),
        .a(6'd12),
        .b(_T_414)
    );
    wire _node_360;
    MUX_UNSIGNED #(.width(1)) u_mux_385 (
        .y(_node_360),
        .sel(_node_359),
        .a(_T_243_12),
        .b(_node_358)
    );
    wire _node_361;
    EQ_UNSIGNED #(.width(6)) u_eq_386 (
        .y(_node_361),
        .a(6'd13),
        .b(_T_414)
    );
    wire _node_362;
    MUX_UNSIGNED #(.width(1)) u_mux_387 (
        .y(_node_362),
        .sel(_node_361),
        .a(_T_243_13),
        .b(_node_360)
    );
    wire _node_363;
    EQ_UNSIGNED #(.width(6)) u_eq_388 (
        .y(_node_363),
        .a(6'd14),
        .b(_T_414)
    );
    wire _node_364;
    MUX_UNSIGNED #(.width(1)) u_mux_389 (
        .y(_node_364),
        .sel(_node_363),
        .a(_T_243_14),
        .b(_node_362)
    );
    wire _node_365;
    EQ_UNSIGNED #(.width(6)) u_eq_390 (
        .y(_node_365),
        .a(6'd15),
        .b(_T_414)
    );
    wire _node_366;
    MUX_UNSIGNED #(.width(1)) u_mux_391 (
        .y(_node_366),
        .sel(_node_365),
        .a(_T_243_15),
        .b(_node_364)
    );
    wire _node_367;
    EQ_UNSIGNED #(.width(6)) u_eq_392 (
        .y(_node_367),
        .a(6'd16),
        .b(_T_414)
    );
    wire _node_368;
    MUX_UNSIGNED #(.width(1)) u_mux_393 (
        .y(_node_368),
        .sel(_node_367),
        .a(_T_243_16),
        .b(_node_366)
    );
    wire _node_369;
    EQ_UNSIGNED #(.width(6)) u_eq_394 (
        .y(_node_369),
        .a(6'd17),
        .b(_T_414)
    );
    wire _node_370;
    MUX_UNSIGNED #(.width(1)) u_mux_395 (
        .y(_node_370),
        .sel(_node_369),
        .a(_T_243_17),
        .b(_node_368)
    );
    wire _node_371;
    EQ_UNSIGNED #(.width(6)) u_eq_396 (
        .y(_node_371),
        .a(6'd18),
        .b(_T_414)
    );
    wire _node_372;
    MUX_UNSIGNED #(.width(1)) u_mux_397 (
        .y(_node_372),
        .sel(_node_371),
        .a(_T_243_18),
        .b(_node_370)
    );
    wire _node_373;
    EQ_UNSIGNED #(.width(6)) u_eq_398 (
        .y(_node_373),
        .a(6'd19),
        .b(_T_414)
    );
    wire _node_374;
    MUX_UNSIGNED #(.width(1)) u_mux_399 (
        .y(_node_374),
        .sel(_node_373),
        .a(_T_243_19),
        .b(_node_372)
    );
    wire _node_375;
    EQ_UNSIGNED #(.width(6)) u_eq_400 (
        .y(_node_375),
        .a(6'd20),
        .b(_T_414)
    );
    wire _node_376;
    MUX_UNSIGNED #(.width(1)) u_mux_401 (
        .y(_node_376),
        .sel(_node_375),
        .a(_T_243_20),
        .b(_node_374)
    );
    wire _node_377;
    EQ_UNSIGNED #(.width(6)) u_eq_402 (
        .y(_node_377),
        .a(6'd21),
        .b(_T_414)
    );
    wire _node_378;
    MUX_UNSIGNED #(.width(1)) u_mux_403 (
        .y(_node_378),
        .sel(_node_377),
        .a(_T_243_21),
        .b(_node_376)
    );
    wire _node_379;
    EQ_UNSIGNED #(.width(6)) u_eq_404 (
        .y(_node_379),
        .a(6'd22),
        .b(_T_414)
    );
    wire _node_380;
    MUX_UNSIGNED #(.width(1)) u_mux_405 (
        .y(_node_380),
        .sel(_node_379),
        .a(_T_243_22),
        .b(_node_378)
    );
    wire _node_381;
    EQ_UNSIGNED #(.width(6)) u_eq_406 (
        .y(_node_381),
        .a(6'd23),
        .b(_T_414)
    );
    wire _node_382;
    MUX_UNSIGNED #(.width(1)) u_mux_407 (
        .y(_node_382),
        .sel(_node_381),
        .a(_T_243_23),
        .b(_node_380)
    );
    wire _node_383;
    EQ_UNSIGNED #(.width(6)) u_eq_408 (
        .y(_node_383),
        .a(6'd24),
        .b(_T_414)
    );
    wire _node_384;
    MUX_UNSIGNED #(.width(1)) u_mux_409 (
        .y(_node_384),
        .sel(_node_383),
        .a(_T_243_24),
        .b(_node_382)
    );
    wire _node_385;
    EQ_UNSIGNED #(.width(6)) u_eq_410 (
        .y(_node_385),
        .a(6'd25),
        .b(_T_414)
    );
    wire _node_386;
    MUX_UNSIGNED #(.width(1)) u_mux_411 (
        .y(_node_386),
        .sel(_node_385),
        .a(_T_243_25),
        .b(_node_384)
    );
    wire _node_387;
    EQ_UNSIGNED #(.width(6)) u_eq_412 (
        .y(_node_387),
        .a(6'd26),
        .b(_T_414)
    );
    wire _node_388;
    MUX_UNSIGNED #(.width(1)) u_mux_413 (
        .y(_node_388),
        .sel(_node_387),
        .a(_T_243_26),
        .b(_node_386)
    );
    wire _node_389;
    EQ_UNSIGNED #(.width(6)) u_eq_414 (
        .y(_node_389),
        .a(6'd27),
        .b(_T_414)
    );
    wire _node_390;
    MUX_UNSIGNED #(.width(1)) u_mux_415 (
        .y(_node_390),
        .sel(_node_389),
        .a(_T_243_27),
        .b(_node_388)
    );
    wire _node_391;
    EQ_UNSIGNED #(.width(6)) u_eq_416 (
        .y(_node_391),
        .a(6'd28),
        .b(_T_414)
    );
    wire _node_392;
    MUX_UNSIGNED #(.width(1)) u_mux_417 (
        .y(_node_392),
        .sel(_node_391),
        .a(_T_243_28),
        .b(_node_390)
    );
    wire _node_393;
    EQ_UNSIGNED #(.width(6)) u_eq_418 (
        .y(_node_393),
        .a(6'd29),
        .b(_T_414)
    );
    wire _node_394;
    MUX_UNSIGNED #(.width(1)) u_mux_419 (
        .y(_node_394),
        .sel(_node_393),
        .a(_T_243_29),
        .b(_node_392)
    );
    wire _node_395;
    EQ_UNSIGNED #(.width(6)) u_eq_420 (
        .y(_node_395),
        .a(6'd30),
        .b(_T_414)
    );
    wire _node_396;
    MUX_UNSIGNED #(.width(1)) u_mux_421 (
        .y(_node_396),
        .sel(_node_395),
        .a(_T_243_30),
        .b(_node_394)
    );
    wire _node_397;
    EQ_UNSIGNED #(.width(6)) u_eq_422 (
        .y(_node_397),
        .a(6'd31),
        .b(_T_414)
    );
    wire _node_398;
    MUX_UNSIGNED #(.width(1)) u_mux_423 (
        .y(_node_398),
        .sel(_node_397),
        .a(_T_243_31),
        .b(_node_396)
    );
    wire _node_399;
    EQ_UNSIGNED #(.width(6)) u_eq_424 (
        .y(_node_399),
        .a(6'd32),
        .b(_T_414)
    );
    wire _node_400;
    MUX_UNSIGNED #(.width(1)) u_mux_425 (
        .y(_node_400),
        .sel(_node_399),
        .a(_T_243_32),
        .b(_node_398)
    );
    wire _node_401;
    EQ_UNSIGNED #(.width(6)) u_eq_426 (
        .y(_node_401),
        .a(6'd33),
        .b(_T_414)
    );
    wire _node_402;
    MUX_UNSIGNED #(.width(1)) u_mux_427 (
        .y(_node_402),
        .sel(_node_401),
        .a(_T_243_33),
        .b(_node_400)
    );
    wire _node_403;
    EQ_UNSIGNED #(.width(6)) u_eq_428 (
        .y(_node_403),
        .a(6'd34),
        .b(_T_414)
    );
    wire _node_404;
    MUX_UNSIGNED #(.width(1)) u_mux_429 (
        .y(_node_404),
        .sel(_node_403),
        .a(_T_243_34),
        .b(_node_402)
    );
    wire _node_405;
    EQ_UNSIGNED #(.width(6)) u_eq_430 (
        .y(_node_405),
        .a(6'd35),
        .b(_T_414)
    );
    wire _node_406;
    MUX_UNSIGNED #(.width(1)) u_mux_431 (
        .y(_node_406),
        .sel(_node_405),
        .a(_T_243_35),
        .b(_node_404)
    );
    wire _node_407;
    EQ_UNSIGNED #(.width(6)) u_eq_432 (
        .y(_node_407),
        .a(6'd36),
        .b(_T_414)
    );
    wire _node_408;
    MUX_UNSIGNED #(.width(1)) u_mux_433 (
        .y(_node_408),
        .sel(_node_407),
        .a(_T_243_36),
        .b(_node_406)
    );
    wire _node_409;
    EQ_UNSIGNED #(.width(6)) u_eq_434 (
        .y(_node_409),
        .a(6'd37),
        .b(_T_414)
    );
    wire _node_410;
    MUX_UNSIGNED #(.width(1)) u_mux_435 (
        .y(_node_410),
        .sel(_node_409),
        .a(_T_243_37),
        .b(_node_408)
    );
    wire _node_411;
    EQ_UNSIGNED #(.width(6)) u_eq_436 (
        .y(_node_411),
        .a(6'd38),
        .b(_T_414)
    );
    wire _node_412;
    MUX_UNSIGNED #(.width(1)) u_mux_437 (
        .y(_node_412),
        .sel(_node_411),
        .a(_T_243_38),
        .b(_node_410)
    );
    wire _node_413;
    EQ_UNSIGNED #(.width(6)) u_eq_438 (
        .y(_node_413),
        .a(6'd39),
        .b(_T_414)
    );
    wire _node_414;
    MUX_UNSIGNED #(.width(1)) u_mux_439 (
        .y(_node_414),
        .sel(_node_413),
        .a(_T_243_39),
        .b(_node_412)
    );
    wire _node_415;
    EQ_UNSIGNED #(.width(6)) u_eq_440 (
        .y(_node_415),
        .a(6'd40),
        .b(_T_414)
    );
    wire _node_416;
    MUX_UNSIGNED #(.width(1)) u_mux_441 (
        .y(_node_416),
        .sel(_node_415),
        .a(_T_243_40),
        .b(_node_414)
    );
    wire _node_417;
    EQ_UNSIGNED #(.width(6)) u_eq_442 (
        .y(_node_417),
        .a(6'd41),
        .b(_T_414)
    );
    wire _node_418;
    MUX_UNSIGNED #(.width(1)) u_mux_443 (
        .y(_node_418),
        .sel(_node_417),
        .a(_T_243_41),
        .b(_node_416)
    );
    wire _node_419;
    EQ_UNSIGNED #(.width(6)) u_eq_444 (
        .y(_node_419),
        .a(6'd42),
        .b(_T_414)
    );
    wire _node_420;
    MUX_UNSIGNED #(.width(1)) u_mux_445 (
        .y(_node_420),
        .sel(_node_419),
        .a(_T_243_42),
        .b(_node_418)
    );
    wire _node_421;
    EQ_UNSIGNED #(.width(6)) u_eq_446 (
        .y(_node_421),
        .a(6'd43),
        .b(_T_414)
    );
    wire _node_422;
    MUX_UNSIGNED #(.width(1)) u_mux_447 (
        .y(_node_422),
        .sel(_node_421),
        .a(_T_243_43),
        .b(_node_420)
    );
    wire _node_423;
    EQ_UNSIGNED #(.width(6)) u_eq_448 (
        .y(_node_423),
        .a(6'd44),
        .b(_T_414)
    );
    wire _node_424;
    MUX_UNSIGNED #(.width(1)) u_mux_449 (
        .y(_node_424),
        .sel(_node_423),
        .a(_T_243_44),
        .b(_node_422)
    );
    wire _node_425;
    EQ_UNSIGNED #(.width(6)) u_eq_450 (
        .y(_node_425),
        .a(6'd45),
        .b(_T_414)
    );
    wire _node_426;
    MUX_UNSIGNED #(.width(1)) u_mux_451 (
        .y(_node_426),
        .sel(_node_425),
        .a(_T_243_45),
        .b(_node_424)
    );
    wire _node_427;
    EQ_UNSIGNED #(.width(6)) u_eq_452 (
        .y(_node_427),
        .a(6'd46),
        .b(_T_414)
    );
    wire _node_428;
    MUX_UNSIGNED #(.width(1)) u_mux_453 (
        .y(_node_428),
        .sel(_node_427),
        .a(_T_243_46),
        .b(_node_426)
    );
    wire _node_429;
    EQ_UNSIGNED #(.width(6)) u_eq_454 (
        .y(_node_429),
        .a(6'd47),
        .b(_T_414)
    );
    wire _node_430;
    MUX_UNSIGNED #(.width(1)) u_mux_455 (
        .y(_node_430),
        .sel(_node_429),
        .a(_T_243_47),
        .b(_node_428)
    );
    wire _node_431;
    EQ_UNSIGNED #(.width(6)) u_eq_456 (
        .y(_node_431),
        .a(6'd48),
        .b(_T_414)
    );
    wire _node_432;
    MUX_UNSIGNED #(.width(1)) u_mux_457 (
        .y(_node_432),
        .sel(_node_431),
        .a(_T_243_48),
        .b(_node_430)
    );
    wire _node_433;
    EQ_UNSIGNED #(.width(6)) u_eq_458 (
        .y(_node_433),
        .a(6'd49),
        .b(_T_414)
    );
    wire _node_434;
    MUX_UNSIGNED #(.width(1)) u_mux_459 (
        .y(_node_434),
        .sel(_node_433),
        .a(_T_243_49),
        .b(_node_432)
    );
    wire _node_435;
    EQ_UNSIGNED #(.width(6)) u_eq_460 (
        .y(_node_435),
        .a(6'd50),
        .b(_T_414)
    );
    wire _node_436;
    MUX_UNSIGNED #(.width(1)) u_mux_461 (
        .y(_node_436),
        .sel(_node_435),
        .a(_T_243_50),
        .b(_node_434)
    );
    wire _node_437;
    EQ_UNSIGNED #(.width(6)) u_eq_462 (
        .y(_node_437),
        .a(6'd51),
        .b(_T_414)
    );
    wire _node_438;
    MUX_UNSIGNED #(.width(1)) u_mux_463 (
        .y(_node_438),
        .sel(_node_437),
        .a(_T_243_51),
        .b(_node_436)
    );
    wire _node_439;
    EQ_UNSIGNED #(.width(6)) u_eq_464 (
        .y(_node_439),
        .a(6'd52),
        .b(_T_414)
    );
    wire _node_440;
    MUX_UNSIGNED #(.width(1)) u_mux_465 (
        .y(_node_440),
        .sel(_node_439),
        .a(_T_243_52),
        .b(_node_438)
    );
    wire _T_415;
    BITWISEAND #(.width(1)) bitwiseand_466 (
        .y(_T_415),
        .a(_c__io_in_valid),
        .b(_c__io_in_ready)
    );
    wire _T_417;
    EQ_UNSIGNED #(.width(5)) u_eq_467 (
        .y(_T_417),
        .a(_value_1__q),
        .b(5'h17)
    );
    wire [5:0] _T_419;
    wire [4:0] _WTEMP_16;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_468 (
        .y(_WTEMP_16),
        .in(1'h1)
    );
    ADD_UNSIGNED #(.width(5)) u_add_469 (
        .y(_T_419),
        .a(_value_1__q),
        .b(_WTEMP_16)
    );
    wire [4:0] _T_420;
    TAIL #(.width(6), .n(1)) tail_470 (
        .y(_T_420),
        .in(_T_419)
    );
    wire _T_423;
    EQ_UNSIGNED #(.width(1)) u_eq_471 (
        .y(_T_423),
        .a(__T_7__q),
        .b(1'h0)
    );
    wire _T_425;
    wire [7:0] _WTEMP_17;
    PAD_UNSIGNED #(.width(6), .n(8)) u_pad_472 (
        .y(_WTEMP_17),
        .in(6'h33)
    );
    EQ_UNSIGNED #(.width(8)) u_eq_473 (
        .y(_T_425),
        .a(__T_4__q),
        .b(_WTEMP_17)
    );
    wire _node_441;
    MUX_UNSIGNED #(.width(1)) u_mux_474 (
        .y(_node_441),
        .sel(_T_173),
        .a(_node_233),
        .b(__T_7__q)
    );
    wire [8:0] _T_428;
    wire [7:0] _WTEMP_18;
    PAD_UNSIGNED #(.width(1), .n(8)) u_pad_475 (
        .y(_WTEMP_18),
        .in(1'h1)
    );
    ADD_UNSIGNED #(.width(8)) u_add_476 (
        .y(_T_428),
        .a(__T_4__q),
        .b(_WTEMP_18)
    );
    wire [7:0] _T_429;
    TAIL #(.width(9), .n(1)) tail_477 (
        .y(_T_429),
        .in(_T_428)
    );
    wire [7:0] _node_442;
    MUX_UNSIGNED #(.width(8)) u_mux_478 (
        .y(_node_442),
        .sel(_T_173),
        .a(_node_232),
        .b(__T_4__q)
    );
    wire _node_443;
    MUX_UNSIGNED #(.width(1)) u_mux_479 (
        .y(_node_443),
        .sel(_T_425),
        .a(1'h1),
        .b(_node_441)
    );
    wire _node_444;
    MUX_UNSIGNED #(.width(1)) u_mux_480 (
        .y(_node_444),
        .sel(_T_173),
        .a(_node_233),
        .b(__T_7__q)
    );
    wire [7:0] _node_445;
    MUX_UNSIGNED #(.width(8)) u_mux_481 (
        .y(_node_445),
        .sel(_T_423),
        .a(_T_429),
        .b(_node_442)
    );
    wire [7:0] _node_446;
    MUX_UNSIGNED #(.width(8)) u_mux_482 (
        .y(_node_446),
        .sel(_T_173),
        .a(_node_232),
        .b(__T_4__q)
    );
    wire _node_447;
    MUX_UNSIGNED #(.width(1)) u_mux_483 (
        .y(_node_447),
        .sel(_T_423),
        .a(_node_443),
        .b(_node_444)
    );
    wire _node_448;
    MUX_UNSIGNED #(.width(1)) u_mux_484 (
        .y(_node_448),
        .sel(_T_173),
        .a(_node_233),
        .b(__T_7__q)
    );
    wire [4:0] _node_449;
    wire [4:0] _WTEMP_19;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_485 (
        .y(_WTEMP_19),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(5)) u_mux_486 (
        .y(_node_449),
        .sel(_T_417),
        .a(_WTEMP_19),
        .b(_T_420)
    );
    wire _T_485_0;
    wire _T_485_1;
    wire _T_485_2;
    wire _T_485_3;
    wire _T_485_4;
    wire _T_485_5;
    wire _T_485_6;
    wire _T_485_7;
    wire _T_485_8;
    wire _T_485_9;
    wire _T_485_10;
    wire _T_485_11;
    wire _T_485_12;
    wire _T_485_13;
    wire _T_485_14;
    wire _T_485_15;
    wire _T_485_16;
    wire _T_485_17;
    wire _T_485_18;
    wire _T_485_19;
    wire _T_485_20;
    wire _T_485_21;
    wire _T_485_22;
    wire _T_485_23;
    wire _T_485_24;
    wire _T_485_25;
    wire _T_485_26;
    wire _T_485_27;
    wire _T_485_28;
    wire _T_485_29;
    wire _T_485_30;
    wire _T_485_31;
    wire _T_485_32;
    wire _T_485_33;
    wire _T_485_34;
    wire _T_485_35;
    wire _T_485_36;
    wire _T_485_37;
    wire _T_485_38;
    wire _T_485_39;
    wire _T_485_40;
    wire _T_485_41;
    wire _T_485_42;
    wire _T_485_43;
    wire _T_485_44;
    wire _T_485_45;
    wire _T_485_46;
    wire _T_485_47;
    wire _T_485_48;
    wire _T_485_49;
    wire _T_485_50;
    wire _T_485_51;
    wire _T_485_52;
    wire [4:0] _value_2__q;
    wire [4:0] _value_2__d;
    DFF_POSCLK #(.width(5)) value_2 (
        .q(_value_2__q),
        .d(_value_2__d),
        .clk(clock)
    );
    wire [4:0] _WTEMP_20;
    MUX_UNSIGNED #(.width(5)) u_mux_487 (
        .y(_value_2__d),
        .sel(reset),
        .a(5'h0),
        .b(_WTEMP_20)
    );
    wire [3:0] _T_565_0;
    wire [3:0] _T_565_1;
    wire [3:0] _T_565_2;
    wire [3:0] _T_565_3;
    wire [3:0] _T_565_4;
    wire [3:0] _T_565_5;
    wire [3:0] _T_565_6;
    wire [3:0] _T_565_7;
    wire [3:0] _T_565_8;
    wire [3:0] _T_565_9;
    wire [3:0] _T_565_10;
    wire [3:0] _T_565_11;
    wire [3:0] _T_565_12;
    wire [3:0] _T_565_13;
    wire [3:0] _T_565_14;
    wire [3:0] _T_565_15;
    wire [3:0] _T_565_16;
    wire [3:0] _T_565_17;
    wire [3:0] _T_565_18;
    wire [3:0] _T_565_19;
    wire [1:0] _T_610_0;
    wire [1:0] _T_610_1;
    wire [1:0] _T_610_2;
    wire [1:0] _T_610_3;
    wire [1:0] _T_610_4;
    wire [1:0] _T_610_5;
    wire [1:0] _T_610_6;
    wire [1:0] _T_610_7;
    wire [1:0] _T_610_8;
    wire [1:0] _T_610_9;
    wire [1:0] _T_610_10;
    wire [1:0] _T_610_11;
    wire [1:0] _T_610_12;
    wire [1:0] _T_610_13;
    wire [1:0] _T_610_14;
    wire [1:0] _T_610_15;
    wire [1:0] _T_610_16;
    wire [1:0] _T_610_17;
    wire [1:0] _T_610_18;
    wire [1:0] _T_610_19;
    wire _node_450;
    EQ_UNSIGNED #(.width(5)) u_eq_488 (
        .y(_node_450),
        .a(5'd0),
        .b(_value_2__q)
    );
    wire [3:0] _node_451;
    assign _node_451 = _T_565_0;
    wire _node_452;
    EQ_UNSIGNED #(.width(5)) u_eq_489 (
        .y(_node_452),
        .a(5'd1),
        .b(_value_2__q)
    );
    wire [3:0] _node_453;
    MUX_UNSIGNED #(.width(4)) u_mux_490 (
        .y(_node_453),
        .sel(_node_452),
        .a(_T_565_1),
        .b(_node_451)
    );
    wire _node_454;
    EQ_UNSIGNED #(.width(5)) u_eq_491 (
        .y(_node_454),
        .a(5'd2),
        .b(_value_2__q)
    );
    wire [3:0] _node_455;
    MUX_UNSIGNED #(.width(4)) u_mux_492 (
        .y(_node_455),
        .sel(_node_454),
        .a(_T_565_2),
        .b(_node_453)
    );
    wire _node_456;
    EQ_UNSIGNED #(.width(5)) u_eq_493 (
        .y(_node_456),
        .a(5'd3),
        .b(_value_2__q)
    );
    wire [3:0] _node_457;
    MUX_UNSIGNED #(.width(4)) u_mux_494 (
        .y(_node_457),
        .sel(_node_456),
        .a(_T_565_3),
        .b(_node_455)
    );
    wire _node_458;
    EQ_UNSIGNED #(.width(5)) u_eq_495 (
        .y(_node_458),
        .a(5'd4),
        .b(_value_2__q)
    );
    wire [3:0] _node_459;
    MUX_UNSIGNED #(.width(4)) u_mux_496 (
        .y(_node_459),
        .sel(_node_458),
        .a(_T_565_4),
        .b(_node_457)
    );
    wire _node_460;
    EQ_UNSIGNED #(.width(5)) u_eq_497 (
        .y(_node_460),
        .a(5'd5),
        .b(_value_2__q)
    );
    wire [3:0] _node_461;
    MUX_UNSIGNED #(.width(4)) u_mux_498 (
        .y(_node_461),
        .sel(_node_460),
        .a(_T_565_5),
        .b(_node_459)
    );
    wire _node_462;
    EQ_UNSIGNED #(.width(5)) u_eq_499 (
        .y(_node_462),
        .a(5'd6),
        .b(_value_2__q)
    );
    wire [3:0] _node_463;
    MUX_UNSIGNED #(.width(4)) u_mux_500 (
        .y(_node_463),
        .sel(_node_462),
        .a(_T_565_6),
        .b(_node_461)
    );
    wire _node_464;
    EQ_UNSIGNED #(.width(5)) u_eq_501 (
        .y(_node_464),
        .a(5'd7),
        .b(_value_2__q)
    );
    wire [3:0] _node_465;
    MUX_UNSIGNED #(.width(4)) u_mux_502 (
        .y(_node_465),
        .sel(_node_464),
        .a(_T_565_7),
        .b(_node_463)
    );
    wire _node_466;
    EQ_UNSIGNED #(.width(5)) u_eq_503 (
        .y(_node_466),
        .a(5'd8),
        .b(_value_2__q)
    );
    wire [3:0] _node_467;
    MUX_UNSIGNED #(.width(4)) u_mux_504 (
        .y(_node_467),
        .sel(_node_466),
        .a(_T_565_8),
        .b(_node_465)
    );
    wire _node_468;
    EQ_UNSIGNED #(.width(5)) u_eq_505 (
        .y(_node_468),
        .a(5'd9),
        .b(_value_2__q)
    );
    wire [3:0] _node_469;
    MUX_UNSIGNED #(.width(4)) u_mux_506 (
        .y(_node_469),
        .sel(_node_468),
        .a(_T_565_9),
        .b(_node_467)
    );
    wire _node_470;
    EQ_UNSIGNED #(.width(5)) u_eq_507 (
        .y(_node_470),
        .a(5'd10),
        .b(_value_2__q)
    );
    wire [3:0] _node_471;
    MUX_UNSIGNED #(.width(4)) u_mux_508 (
        .y(_node_471),
        .sel(_node_470),
        .a(_T_565_10),
        .b(_node_469)
    );
    wire _node_472;
    EQ_UNSIGNED #(.width(5)) u_eq_509 (
        .y(_node_472),
        .a(5'd11),
        .b(_value_2__q)
    );
    wire [3:0] _node_473;
    MUX_UNSIGNED #(.width(4)) u_mux_510 (
        .y(_node_473),
        .sel(_node_472),
        .a(_T_565_11),
        .b(_node_471)
    );
    wire _node_474;
    EQ_UNSIGNED #(.width(5)) u_eq_511 (
        .y(_node_474),
        .a(5'd12),
        .b(_value_2__q)
    );
    wire [3:0] _node_475;
    MUX_UNSIGNED #(.width(4)) u_mux_512 (
        .y(_node_475),
        .sel(_node_474),
        .a(_T_565_12),
        .b(_node_473)
    );
    wire _node_476;
    EQ_UNSIGNED #(.width(5)) u_eq_513 (
        .y(_node_476),
        .a(5'd13),
        .b(_value_2__q)
    );
    wire [3:0] _node_477;
    MUX_UNSIGNED #(.width(4)) u_mux_514 (
        .y(_node_477),
        .sel(_node_476),
        .a(_T_565_13),
        .b(_node_475)
    );
    wire _node_478;
    EQ_UNSIGNED #(.width(5)) u_eq_515 (
        .y(_node_478),
        .a(5'd14),
        .b(_value_2__q)
    );
    wire [3:0] _node_479;
    MUX_UNSIGNED #(.width(4)) u_mux_516 (
        .y(_node_479),
        .sel(_node_478),
        .a(_T_565_14),
        .b(_node_477)
    );
    wire _node_480;
    EQ_UNSIGNED #(.width(5)) u_eq_517 (
        .y(_node_480),
        .a(5'd15),
        .b(_value_2__q)
    );
    wire [3:0] _node_481;
    MUX_UNSIGNED #(.width(4)) u_mux_518 (
        .y(_node_481),
        .sel(_node_480),
        .a(_T_565_15),
        .b(_node_479)
    );
    wire _node_482;
    EQ_UNSIGNED #(.width(5)) u_eq_519 (
        .y(_node_482),
        .a(5'd16),
        .b(_value_2__q)
    );
    wire [3:0] _node_483;
    MUX_UNSIGNED #(.width(4)) u_mux_520 (
        .y(_node_483),
        .sel(_node_482),
        .a(_T_565_16),
        .b(_node_481)
    );
    wire _node_484;
    EQ_UNSIGNED #(.width(5)) u_eq_521 (
        .y(_node_484),
        .a(5'd17),
        .b(_value_2__q)
    );
    wire [3:0] _node_485;
    MUX_UNSIGNED #(.width(4)) u_mux_522 (
        .y(_node_485),
        .sel(_node_484),
        .a(_T_565_17),
        .b(_node_483)
    );
    wire _node_486;
    EQ_UNSIGNED #(.width(5)) u_eq_523 (
        .y(_node_486),
        .a(5'd18),
        .b(_value_2__q)
    );
    wire [3:0] _node_487;
    MUX_UNSIGNED #(.width(4)) u_mux_524 (
        .y(_node_487),
        .sel(_node_486),
        .a(_T_565_18),
        .b(_node_485)
    );
    wire _node_488;
    EQ_UNSIGNED #(.width(5)) u_eq_525 (
        .y(_node_488),
        .a(5'd19),
        .b(_value_2__q)
    );
    wire [3:0] _node_489;
    MUX_UNSIGNED #(.width(4)) u_mux_526 (
        .y(_node_489),
        .sel(_node_488),
        .a(_T_565_19),
        .b(_node_487)
    );
    wire _node_490;
    EQ_UNSIGNED #(.width(5)) u_eq_527 (
        .y(_node_490),
        .a(5'd0),
        .b(_value_2__q)
    );
    wire [1:0] _node_491;
    assign _node_491 = _T_610_0;
    wire _node_492;
    EQ_UNSIGNED #(.width(5)) u_eq_528 (
        .y(_node_492),
        .a(5'd1),
        .b(_value_2__q)
    );
    wire [1:0] _node_493;
    MUX_UNSIGNED #(.width(2)) u_mux_529 (
        .y(_node_493),
        .sel(_node_492),
        .a(_T_610_1),
        .b(_node_491)
    );
    wire _node_494;
    EQ_UNSIGNED #(.width(5)) u_eq_530 (
        .y(_node_494),
        .a(5'd2),
        .b(_value_2__q)
    );
    wire [1:0] _node_495;
    MUX_UNSIGNED #(.width(2)) u_mux_531 (
        .y(_node_495),
        .sel(_node_494),
        .a(_T_610_2),
        .b(_node_493)
    );
    wire _node_496;
    EQ_UNSIGNED #(.width(5)) u_eq_532 (
        .y(_node_496),
        .a(5'd3),
        .b(_value_2__q)
    );
    wire [1:0] _node_497;
    MUX_UNSIGNED #(.width(2)) u_mux_533 (
        .y(_node_497),
        .sel(_node_496),
        .a(_T_610_3),
        .b(_node_495)
    );
    wire _node_498;
    EQ_UNSIGNED #(.width(5)) u_eq_534 (
        .y(_node_498),
        .a(5'd4),
        .b(_value_2__q)
    );
    wire [1:0] _node_499;
    MUX_UNSIGNED #(.width(2)) u_mux_535 (
        .y(_node_499),
        .sel(_node_498),
        .a(_T_610_4),
        .b(_node_497)
    );
    wire _node_500;
    EQ_UNSIGNED #(.width(5)) u_eq_536 (
        .y(_node_500),
        .a(5'd5),
        .b(_value_2__q)
    );
    wire [1:0] _node_501;
    MUX_UNSIGNED #(.width(2)) u_mux_537 (
        .y(_node_501),
        .sel(_node_500),
        .a(_T_610_5),
        .b(_node_499)
    );
    wire _node_502;
    EQ_UNSIGNED #(.width(5)) u_eq_538 (
        .y(_node_502),
        .a(5'd6),
        .b(_value_2__q)
    );
    wire [1:0] _node_503;
    MUX_UNSIGNED #(.width(2)) u_mux_539 (
        .y(_node_503),
        .sel(_node_502),
        .a(_T_610_6),
        .b(_node_501)
    );
    wire _node_504;
    EQ_UNSIGNED #(.width(5)) u_eq_540 (
        .y(_node_504),
        .a(5'd7),
        .b(_value_2__q)
    );
    wire [1:0] _node_505;
    MUX_UNSIGNED #(.width(2)) u_mux_541 (
        .y(_node_505),
        .sel(_node_504),
        .a(_T_610_7),
        .b(_node_503)
    );
    wire _node_506;
    EQ_UNSIGNED #(.width(5)) u_eq_542 (
        .y(_node_506),
        .a(5'd8),
        .b(_value_2__q)
    );
    wire [1:0] _node_507;
    MUX_UNSIGNED #(.width(2)) u_mux_543 (
        .y(_node_507),
        .sel(_node_506),
        .a(_T_610_8),
        .b(_node_505)
    );
    wire _node_508;
    EQ_UNSIGNED #(.width(5)) u_eq_544 (
        .y(_node_508),
        .a(5'd9),
        .b(_value_2__q)
    );
    wire [1:0] _node_509;
    MUX_UNSIGNED #(.width(2)) u_mux_545 (
        .y(_node_509),
        .sel(_node_508),
        .a(_T_610_9),
        .b(_node_507)
    );
    wire _node_510;
    EQ_UNSIGNED #(.width(5)) u_eq_546 (
        .y(_node_510),
        .a(5'd10),
        .b(_value_2__q)
    );
    wire [1:0] _node_511;
    MUX_UNSIGNED #(.width(2)) u_mux_547 (
        .y(_node_511),
        .sel(_node_510),
        .a(_T_610_10),
        .b(_node_509)
    );
    wire _node_512;
    EQ_UNSIGNED #(.width(5)) u_eq_548 (
        .y(_node_512),
        .a(5'd11),
        .b(_value_2__q)
    );
    wire [1:0] _node_513;
    MUX_UNSIGNED #(.width(2)) u_mux_549 (
        .y(_node_513),
        .sel(_node_512),
        .a(_T_610_11),
        .b(_node_511)
    );
    wire _node_514;
    EQ_UNSIGNED #(.width(5)) u_eq_550 (
        .y(_node_514),
        .a(5'd12),
        .b(_value_2__q)
    );
    wire [1:0] _node_515;
    MUX_UNSIGNED #(.width(2)) u_mux_551 (
        .y(_node_515),
        .sel(_node_514),
        .a(_T_610_12),
        .b(_node_513)
    );
    wire _node_516;
    EQ_UNSIGNED #(.width(5)) u_eq_552 (
        .y(_node_516),
        .a(5'd13),
        .b(_value_2__q)
    );
    wire [1:0] _node_517;
    MUX_UNSIGNED #(.width(2)) u_mux_553 (
        .y(_node_517),
        .sel(_node_516),
        .a(_T_610_13),
        .b(_node_515)
    );
    wire _node_518;
    EQ_UNSIGNED #(.width(5)) u_eq_554 (
        .y(_node_518),
        .a(5'd14),
        .b(_value_2__q)
    );
    wire [1:0] _node_519;
    MUX_UNSIGNED #(.width(2)) u_mux_555 (
        .y(_node_519),
        .sel(_node_518),
        .a(_T_610_14),
        .b(_node_517)
    );
    wire _node_520;
    EQ_UNSIGNED #(.width(5)) u_eq_556 (
        .y(_node_520),
        .a(5'd15),
        .b(_value_2__q)
    );
    wire [1:0] _node_521;
    MUX_UNSIGNED #(.width(2)) u_mux_557 (
        .y(_node_521),
        .sel(_node_520),
        .a(_T_610_15),
        .b(_node_519)
    );
    wire _node_522;
    EQ_UNSIGNED #(.width(5)) u_eq_558 (
        .y(_node_522),
        .a(5'd16),
        .b(_value_2__q)
    );
    wire [1:0] _node_523;
    MUX_UNSIGNED #(.width(2)) u_mux_559 (
        .y(_node_523),
        .sel(_node_522),
        .a(_T_610_16),
        .b(_node_521)
    );
    wire _node_524;
    EQ_UNSIGNED #(.width(5)) u_eq_560 (
        .y(_node_524),
        .a(5'd17),
        .b(_value_2__q)
    );
    wire [1:0] _node_525;
    MUX_UNSIGNED #(.width(2)) u_mux_561 (
        .y(_node_525),
        .sel(_node_524),
        .a(_T_610_17),
        .b(_node_523)
    );
    wire _node_526;
    EQ_UNSIGNED #(.width(5)) u_eq_562 (
        .y(_node_526),
        .a(5'd18),
        .b(_value_2__q)
    );
    wire [1:0] _node_527;
    MUX_UNSIGNED #(.width(2)) u_mux_563 (
        .y(_node_527),
        .sel(_node_526),
        .a(_T_610_18),
        .b(_node_525)
    );
    wire _node_528;
    EQ_UNSIGNED #(.width(5)) u_eq_564 (
        .y(_node_528),
        .a(5'd19),
        .b(_value_2__q)
    );
    wire [1:0] _node_529;
    MUX_UNSIGNED #(.width(2)) u_mux_565 (
        .y(_node_529),
        .sel(_node_528),
        .a(_T_610_19),
        .b(_node_527)
    );
    wire [5:0] _T_636;
    BITS #(.width(8), .high(5), .low(0)) bits_566 (
        .y(_T_636),
        .in(__T_4__q)
    );
    wire _node_530;
    EQ_UNSIGNED #(.width(6)) u_eq_567 (
        .y(_node_530),
        .a(6'd0),
        .b(_T_636)
    );
    wire _node_531;
    assign _node_531 = _T_485_0;
    wire _node_532;
    EQ_UNSIGNED #(.width(6)) u_eq_568 (
        .y(_node_532),
        .a(6'd1),
        .b(_T_636)
    );
    wire _node_533;
    MUX_UNSIGNED #(.width(1)) u_mux_569 (
        .y(_node_533),
        .sel(_node_532),
        .a(_T_485_1),
        .b(_node_531)
    );
    wire _node_534;
    EQ_UNSIGNED #(.width(6)) u_eq_570 (
        .y(_node_534),
        .a(6'd2),
        .b(_T_636)
    );
    wire _node_535;
    MUX_UNSIGNED #(.width(1)) u_mux_571 (
        .y(_node_535),
        .sel(_node_534),
        .a(_T_485_2),
        .b(_node_533)
    );
    wire _node_536;
    EQ_UNSIGNED #(.width(6)) u_eq_572 (
        .y(_node_536),
        .a(6'd3),
        .b(_T_636)
    );
    wire _node_537;
    MUX_UNSIGNED #(.width(1)) u_mux_573 (
        .y(_node_537),
        .sel(_node_536),
        .a(_T_485_3),
        .b(_node_535)
    );
    wire _node_538;
    EQ_UNSIGNED #(.width(6)) u_eq_574 (
        .y(_node_538),
        .a(6'd4),
        .b(_T_636)
    );
    wire _node_539;
    MUX_UNSIGNED #(.width(1)) u_mux_575 (
        .y(_node_539),
        .sel(_node_538),
        .a(_T_485_4),
        .b(_node_537)
    );
    wire _node_540;
    EQ_UNSIGNED #(.width(6)) u_eq_576 (
        .y(_node_540),
        .a(6'd5),
        .b(_T_636)
    );
    wire _node_541;
    MUX_UNSIGNED #(.width(1)) u_mux_577 (
        .y(_node_541),
        .sel(_node_540),
        .a(_T_485_5),
        .b(_node_539)
    );
    wire _node_542;
    EQ_UNSIGNED #(.width(6)) u_eq_578 (
        .y(_node_542),
        .a(6'd6),
        .b(_T_636)
    );
    wire _node_543;
    MUX_UNSIGNED #(.width(1)) u_mux_579 (
        .y(_node_543),
        .sel(_node_542),
        .a(_T_485_6),
        .b(_node_541)
    );
    wire _node_544;
    EQ_UNSIGNED #(.width(6)) u_eq_580 (
        .y(_node_544),
        .a(6'd7),
        .b(_T_636)
    );
    wire _node_545;
    MUX_UNSIGNED #(.width(1)) u_mux_581 (
        .y(_node_545),
        .sel(_node_544),
        .a(_T_485_7),
        .b(_node_543)
    );
    wire _node_546;
    EQ_UNSIGNED #(.width(6)) u_eq_582 (
        .y(_node_546),
        .a(6'd8),
        .b(_T_636)
    );
    wire _node_547;
    MUX_UNSIGNED #(.width(1)) u_mux_583 (
        .y(_node_547),
        .sel(_node_546),
        .a(_T_485_8),
        .b(_node_545)
    );
    wire _node_548;
    EQ_UNSIGNED #(.width(6)) u_eq_584 (
        .y(_node_548),
        .a(6'd9),
        .b(_T_636)
    );
    wire _node_549;
    MUX_UNSIGNED #(.width(1)) u_mux_585 (
        .y(_node_549),
        .sel(_node_548),
        .a(_T_485_9),
        .b(_node_547)
    );
    wire _node_550;
    EQ_UNSIGNED #(.width(6)) u_eq_586 (
        .y(_node_550),
        .a(6'd10),
        .b(_T_636)
    );
    wire _node_551;
    MUX_UNSIGNED #(.width(1)) u_mux_587 (
        .y(_node_551),
        .sel(_node_550),
        .a(_T_485_10),
        .b(_node_549)
    );
    wire _node_552;
    EQ_UNSIGNED #(.width(6)) u_eq_588 (
        .y(_node_552),
        .a(6'd11),
        .b(_T_636)
    );
    wire _node_553;
    MUX_UNSIGNED #(.width(1)) u_mux_589 (
        .y(_node_553),
        .sel(_node_552),
        .a(_T_485_11),
        .b(_node_551)
    );
    wire _node_554;
    EQ_UNSIGNED #(.width(6)) u_eq_590 (
        .y(_node_554),
        .a(6'd12),
        .b(_T_636)
    );
    wire _node_555;
    MUX_UNSIGNED #(.width(1)) u_mux_591 (
        .y(_node_555),
        .sel(_node_554),
        .a(_T_485_12),
        .b(_node_553)
    );
    wire _node_556;
    EQ_UNSIGNED #(.width(6)) u_eq_592 (
        .y(_node_556),
        .a(6'd13),
        .b(_T_636)
    );
    wire _node_557;
    MUX_UNSIGNED #(.width(1)) u_mux_593 (
        .y(_node_557),
        .sel(_node_556),
        .a(_T_485_13),
        .b(_node_555)
    );
    wire _node_558;
    EQ_UNSIGNED #(.width(6)) u_eq_594 (
        .y(_node_558),
        .a(6'd14),
        .b(_T_636)
    );
    wire _node_559;
    MUX_UNSIGNED #(.width(1)) u_mux_595 (
        .y(_node_559),
        .sel(_node_558),
        .a(_T_485_14),
        .b(_node_557)
    );
    wire _node_560;
    EQ_UNSIGNED #(.width(6)) u_eq_596 (
        .y(_node_560),
        .a(6'd15),
        .b(_T_636)
    );
    wire _node_561;
    MUX_UNSIGNED #(.width(1)) u_mux_597 (
        .y(_node_561),
        .sel(_node_560),
        .a(_T_485_15),
        .b(_node_559)
    );
    wire _node_562;
    EQ_UNSIGNED #(.width(6)) u_eq_598 (
        .y(_node_562),
        .a(6'd16),
        .b(_T_636)
    );
    wire _node_563;
    MUX_UNSIGNED #(.width(1)) u_mux_599 (
        .y(_node_563),
        .sel(_node_562),
        .a(_T_485_16),
        .b(_node_561)
    );
    wire _node_564;
    EQ_UNSIGNED #(.width(6)) u_eq_600 (
        .y(_node_564),
        .a(6'd17),
        .b(_T_636)
    );
    wire _node_565;
    MUX_UNSIGNED #(.width(1)) u_mux_601 (
        .y(_node_565),
        .sel(_node_564),
        .a(_T_485_17),
        .b(_node_563)
    );
    wire _node_566;
    EQ_UNSIGNED #(.width(6)) u_eq_602 (
        .y(_node_566),
        .a(6'd18),
        .b(_T_636)
    );
    wire _node_567;
    MUX_UNSIGNED #(.width(1)) u_mux_603 (
        .y(_node_567),
        .sel(_node_566),
        .a(_T_485_18),
        .b(_node_565)
    );
    wire _node_568;
    EQ_UNSIGNED #(.width(6)) u_eq_604 (
        .y(_node_568),
        .a(6'd19),
        .b(_T_636)
    );
    wire _node_569;
    MUX_UNSIGNED #(.width(1)) u_mux_605 (
        .y(_node_569),
        .sel(_node_568),
        .a(_T_485_19),
        .b(_node_567)
    );
    wire _node_570;
    EQ_UNSIGNED #(.width(6)) u_eq_606 (
        .y(_node_570),
        .a(6'd20),
        .b(_T_636)
    );
    wire _node_571;
    MUX_UNSIGNED #(.width(1)) u_mux_607 (
        .y(_node_571),
        .sel(_node_570),
        .a(_T_485_20),
        .b(_node_569)
    );
    wire _node_572;
    EQ_UNSIGNED #(.width(6)) u_eq_608 (
        .y(_node_572),
        .a(6'd21),
        .b(_T_636)
    );
    wire _node_573;
    MUX_UNSIGNED #(.width(1)) u_mux_609 (
        .y(_node_573),
        .sel(_node_572),
        .a(_T_485_21),
        .b(_node_571)
    );
    wire _node_574;
    EQ_UNSIGNED #(.width(6)) u_eq_610 (
        .y(_node_574),
        .a(6'd22),
        .b(_T_636)
    );
    wire _node_575;
    MUX_UNSIGNED #(.width(1)) u_mux_611 (
        .y(_node_575),
        .sel(_node_574),
        .a(_T_485_22),
        .b(_node_573)
    );
    wire _node_576;
    EQ_UNSIGNED #(.width(6)) u_eq_612 (
        .y(_node_576),
        .a(6'd23),
        .b(_T_636)
    );
    wire _node_577;
    MUX_UNSIGNED #(.width(1)) u_mux_613 (
        .y(_node_577),
        .sel(_node_576),
        .a(_T_485_23),
        .b(_node_575)
    );
    wire _node_578;
    EQ_UNSIGNED #(.width(6)) u_eq_614 (
        .y(_node_578),
        .a(6'd24),
        .b(_T_636)
    );
    wire _node_579;
    MUX_UNSIGNED #(.width(1)) u_mux_615 (
        .y(_node_579),
        .sel(_node_578),
        .a(_T_485_24),
        .b(_node_577)
    );
    wire _node_580;
    EQ_UNSIGNED #(.width(6)) u_eq_616 (
        .y(_node_580),
        .a(6'd25),
        .b(_T_636)
    );
    wire _node_581;
    MUX_UNSIGNED #(.width(1)) u_mux_617 (
        .y(_node_581),
        .sel(_node_580),
        .a(_T_485_25),
        .b(_node_579)
    );
    wire _node_582;
    EQ_UNSIGNED #(.width(6)) u_eq_618 (
        .y(_node_582),
        .a(6'd26),
        .b(_T_636)
    );
    wire _node_583;
    MUX_UNSIGNED #(.width(1)) u_mux_619 (
        .y(_node_583),
        .sel(_node_582),
        .a(_T_485_26),
        .b(_node_581)
    );
    wire _node_584;
    EQ_UNSIGNED #(.width(6)) u_eq_620 (
        .y(_node_584),
        .a(6'd27),
        .b(_T_636)
    );
    wire _node_585;
    MUX_UNSIGNED #(.width(1)) u_mux_621 (
        .y(_node_585),
        .sel(_node_584),
        .a(_T_485_27),
        .b(_node_583)
    );
    wire _node_586;
    EQ_UNSIGNED #(.width(6)) u_eq_622 (
        .y(_node_586),
        .a(6'd28),
        .b(_T_636)
    );
    wire _node_587;
    MUX_UNSIGNED #(.width(1)) u_mux_623 (
        .y(_node_587),
        .sel(_node_586),
        .a(_T_485_28),
        .b(_node_585)
    );
    wire _node_588;
    EQ_UNSIGNED #(.width(6)) u_eq_624 (
        .y(_node_588),
        .a(6'd29),
        .b(_T_636)
    );
    wire _node_589;
    MUX_UNSIGNED #(.width(1)) u_mux_625 (
        .y(_node_589),
        .sel(_node_588),
        .a(_T_485_29),
        .b(_node_587)
    );
    wire _node_590;
    EQ_UNSIGNED #(.width(6)) u_eq_626 (
        .y(_node_590),
        .a(6'd30),
        .b(_T_636)
    );
    wire _node_591;
    MUX_UNSIGNED #(.width(1)) u_mux_627 (
        .y(_node_591),
        .sel(_node_590),
        .a(_T_485_30),
        .b(_node_589)
    );
    wire _node_592;
    EQ_UNSIGNED #(.width(6)) u_eq_628 (
        .y(_node_592),
        .a(6'd31),
        .b(_T_636)
    );
    wire _node_593;
    MUX_UNSIGNED #(.width(1)) u_mux_629 (
        .y(_node_593),
        .sel(_node_592),
        .a(_T_485_31),
        .b(_node_591)
    );
    wire _node_594;
    EQ_UNSIGNED #(.width(6)) u_eq_630 (
        .y(_node_594),
        .a(6'd32),
        .b(_T_636)
    );
    wire _node_595;
    MUX_UNSIGNED #(.width(1)) u_mux_631 (
        .y(_node_595),
        .sel(_node_594),
        .a(_T_485_32),
        .b(_node_593)
    );
    wire _node_596;
    EQ_UNSIGNED #(.width(6)) u_eq_632 (
        .y(_node_596),
        .a(6'd33),
        .b(_T_636)
    );
    wire _node_597;
    MUX_UNSIGNED #(.width(1)) u_mux_633 (
        .y(_node_597),
        .sel(_node_596),
        .a(_T_485_33),
        .b(_node_595)
    );
    wire _node_598;
    EQ_UNSIGNED #(.width(6)) u_eq_634 (
        .y(_node_598),
        .a(6'd34),
        .b(_T_636)
    );
    wire _node_599;
    MUX_UNSIGNED #(.width(1)) u_mux_635 (
        .y(_node_599),
        .sel(_node_598),
        .a(_T_485_34),
        .b(_node_597)
    );
    wire _node_600;
    EQ_UNSIGNED #(.width(6)) u_eq_636 (
        .y(_node_600),
        .a(6'd35),
        .b(_T_636)
    );
    wire _node_601;
    MUX_UNSIGNED #(.width(1)) u_mux_637 (
        .y(_node_601),
        .sel(_node_600),
        .a(_T_485_35),
        .b(_node_599)
    );
    wire _node_602;
    EQ_UNSIGNED #(.width(6)) u_eq_638 (
        .y(_node_602),
        .a(6'd36),
        .b(_T_636)
    );
    wire _node_603;
    MUX_UNSIGNED #(.width(1)) u_mux_639 (
        .y(_node_603),
        .sel(_node_602),
        .a(_T_485_36),
        .b(_node_601)
    );
    wire _node_604;
    EQ_UNSIGNED #(.width(6)) u_eq_640 (
        .y(_node_604),
        .a(6'd37),
        .b(_T_636)
    );
    wire _node_605;
    MUX_UNSIGNED #(.width(1)) u_mux_641 (
        .y(_node_605),
        .sel(_node_604),
        .a(_T_485_37),
        .b(_node_603)
    );
    wire _node_606;
    EQ_UNSIGNED #(.width(6)) u_eq_642 (
        .y(_node_606),
        .a(6'd38),
        .b(_T_636)
    );
    wire _node_607;
    MUX_UNSIGNED #(.width(1)) u_mux_643 (
        .y(_node_607),
        .sel(_node_606),
        .a(_T_485_38),
        .b(_node_605)
    );
    wire _node_608;
    EQ_UNSIGNED #(.width(6)) u_eq_644 (
        .y(_node_608),
        .a(6'd39),
        .b(_T_636)
    );
    wire _node_609;
    MUX_UNSIGNED #(.width(1)) u_mux_645 (
        .y(_node_609),
        .sel(_node_608),
        .a(_T_485_39),
        .b(_node_607)
    );
    wire _node_610;
    EQ_UNSIGNED #(.width(6)) u_eq_646 (
        .y(_node_610),
        .a(6'd40),
        .b(_T_636)
    );
    wire _node_611;
    MUX_UNSIGNED #(.width(1)) u_mux_647 (
        .y(_node_611),
        .sel(_node_610),
        .a(_T_485_40),
        .b(_node_609)
    );
    wire _node_612;
    EQ_UNSIGNED #(.width(6)) u_eq_648 (
        .y(_node_612),
        .a(6'd41),
        .b(_T_636)
    );
    wire _node_613;
    MUX_UNSIGNED #(.width(1)) u_mux_649 (
        .y(_node_613),
        .sel(_node_612),
        .a(_T_485_41),
        .b(_node_611)
    );
    wire _node_614;
    EQ_UNSIGNED #(.width(6)) u_eq_650 (
        .y(_node_614),
        .a(6'd42),
        .b(_T_636)
    );
    wire _node_615;
    MUX_UNSIGNED #(.width(1)) u_mux_651 (
        .y(_node_615),
        .sel(_node_614),
        .a(_T_485_42),
        .b(_node_613)
    );
    wire _node_616;
    EQ_UNSIGNED #(.width(6)) u_eq_652 (
        .y(_node_616),
        .a(6'd43),
        .b(_T_636)
    );
    wire _node_617;
    MUX_UNSIGNED #(.width(1)) u_mux_653 (
        .y(_node_617),
        .sel(_node_616),
        .a(_T_485_43),
        .b(_node_615)
    );
    wire _node_618;
    EQ_UNSIGNED #(.width(6)) u_eq_654 (
        .y(_node_618),
        .a(6'd44),
        .b(_T_636)
    );
    wire _node_619;
    MUX_UNSIGNED #(.width(1)) u_mux_655 (
        .y(_node_619),
        .sel(_node_618),
        .a(_T_485_44),
        .b(_node_617)
    );
    wire _node_620;
    EQ_UNSIGNED #(.width(6)) u_eq_656 (
        .y(_node_620),
        .a(6'd45),
        .b(_T_636)
    );
    wire _node_621;
    MUX_UNSIGNED #(.width(1)) u_mux_657 (
        .y(_node_621),
        .sel(_node_620),
        .a(_T_485_45),
        .b(_node_619)
    );
    wire _node_622;
    EQ_UNSIGNED #(.width(6)) u_eq_658 (
        .y(_node_622),
        .a(6'd46),
        .b(_T_636)
    );
    wire _node_623;
    MUX_UNSIGNED #(.width(1)) u_mux_659 (
        .y(_node_623),
        .sel(_node_622),
        .a(_T_485_46),
        .b(_node_621)
    );
    wire _node_624;
    EQ_UNSIGNED #(.width(6)) u_eq_660 (
        .y(_node_624),
        .a(6'd47),
        .b(_T_636)
    );
    wire _node_625;
    MUX_UNSIGNED #(.width(1)) u_mux_661 (
        .y(_node_625),
        .sel(_node_624),
        .a(_T_485_47),
        .b(_node_623)
    );
    wire _node_626;
    EQ_UNSIGNED #(.width(6)) u_eq_662 (
        .y(_node_626),
        .a(6'd48),
        .b(_T_636)
    );
    wire _node_627;
    MUX_UNSIGNED #(.width(1)) u_mux_663 (
        .y(_node_627),
        .sel(_node_626),
        .a(_T_485_48),
        .b(_node_625)
    );
    wire _node_628;
    EQ_UNSIGNED #(.width(6)) u_eq_664 (
        .y(_node_628),
        .a(6'd49),
        .b(_T_636)
    );
    wire _node_629;
    MUX_UNSIGNED #(.width(1)) u_mux_665 (
        .y(_node_629),
        .sel(_node_628),
        .a(_T_485_49),
        .b(_node_627)
    );
    wire _node_630;
    EQ_UNSIGNED #(.width(6)) u_eq_666 (
        .y(_node_630),
        .a(6'd50),
        .b(_T_636)
    );
    wire _node_631;
    MUX_UNSIGNED #(.width(1)) u_mux_667 (
        .y(_node_631),
        .sel(_node_630),
        .a(_T_485_50),
        .b(_node_629)
    );
    wire _node_632;
    EQ_UNSIGNED #(.width(6)) u_eq_668 (
        .y(_node_632),
        .a(6'd51),
        .b(_T_636)
    );
    wire _node_633;
    MUX_UNSIGNED #(.width(1)) u_mux_669 (
        .y(_node_633),
        .sel(_node_632),
        .a(_T_485_51),
        .b(_node_631)
    );
    wire _node_634;
    EQ_UNSIGNED #(.width(6)) u_eq_670 (
        .y(_node_634),
        .a(6'd52),
        .b(_T_636)
    );
    wire _node_635;
    MUX_UNSIGNED #(.width(1)) u_mux_671 (
        .y(_node_635),
        .sel(_node_634),
        .a(_T_485_52),
        .b(_node_633)
    );
    wire _T_637;
    BITWISEAND #(.width(1)) bitwiseand_672 (
        .y(_T_637),
        .a(_c__io_load_routing_table_request_valid),
        .b(_c__io_load_routing_table_request_ready)
    );
    wire _T_639;
    EQ_UNSIGNED #(.width(5)) u_eq_673 (
        .y(_T_639),
        .a(_value_2__q),
        .b(5'h12)
    );
    wire [5:0] _T_641;
    wire [4:0] _WTEMP_21;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_674 (
        .y(_WTEMP_21),
        .in(1'h1)
    );
    ADD_UNSIGNED #(.width(5)) u_add_675 (
        .y(_T_641),
        .a(_value_2__q),
        .b(_WTEMP_21)
    );
    wire [4:0] _T_642;
    TAIL #(.width(6), .n(1)) tail_676 (
        .y(_T_642),
        .in(_T_641)
    );
    wire _T_645;
    EQ_UNSIGNED #(.width(1)) u_eq_677 (
        .y(_T_645),
        .a(__T_7__q),
        .b(1'h0)
    );
    wire _T_647;
    wire [7:0] _WTEMP_22;
    PAD_UNSIGNED #(.width(6), .n(8)) u_pad_678 (
        .y(_WTEMP_22),
        .in(6'h33)
    );
    EQ_UNSIGNED #(.width(8)) u_eq_679 (
        .y(_T_647),
        .a(__T_4__q),
        .b(_WTEMP_22)
    );
    wire _node_636;
    MUX_UNSIGNED #(.width(1)) u_mux_680 (
        .y(_node_636),
        .sel(_T_415),
        .a(_node_447),
        .b(_node_448)
    );
    wire [8:0] _T_650;
    wire [7:0] _WTEMP_23;
    PAD_UNSIGNED #(.width(1), .n(8)) u_pad_681 (
        .y(_WTEMP_23),
        .in(1'h1)
    );
    ADD_UNSIGNED #(.width(8)) u_add_682 (
        .y(_T_650),
        .a(__T_4__q),
        .b(_WTEMP_23)
    );
    wire [7:0] _T_651;
    TAIL #(.width(9), .n(1)) tail_683 (
        .y(_T_651),
        .in(_T_650)
    );
    wire [7:0] _node_637;
    MUX_UNSIGNED #(.width(8)) u_mux_684 (
        .y(_node_637),
        .sel(_T_415),
        .a(_node_445),
        .b(_node_446)
    );
    wire _node_638;
    MUX_UNSIGNED #(.width(1)) u_mux_685 (
        .y(_node_638),
        .sel(_T_647),
        .a(1'h1),
        .b(_node_636)
    );
    wire _node_639;
    MUX_UNSIGNED #(.width(1)) u_mux_686 (
        .y(_node_639),
        .sel(_T_415),
        .a(_node_447),
        .b(_node_448)
    );
    wire [7:0] _node_640;
    MUX_UNSIGNED #(.width(8)) u_mux_687 (
        .y(_node_640),
        .sel(_T_645),
        .a(_T_651),
        .b(_node_637)
    );
    wire [7:0] _node_641;
    MUX_UNSIGNED #(.width(8)) u_mux_688 (
        .y(_node_641),
        .sel(_T_415),
        .a(_node_445),
        .b(_node_446)
    );
    wire _node_642;
    MUX_UNSIGNED #(.width(1)) u_mux_689 (
        .y(_node_642),
        .sel(_T_645),
        .a(_node_638),
        .b(_node_639)
    );
    wire _node_643;
    MUX_UNSIGNED #(.width(1)) u_mux_690 (
        .y(_node_643),
        .sel(_T_415),
        .a(_node_447),
        .b(_node_448)
    );
    wire [4:0] _node_644;
    wire [4:0] _WTEMP_24;
    PAD_UNSIGNED #(.width(1), .n(5)) u_pad_691 (
        .y(_WTEMP_24),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(5)) u_mux_692 (
        .y(_node_644),
        .sel(_T_639),
        .a(_WTEMP_24),
        .b(_T_642)
    );
    wire _T_707_0;
    wire _T_707_1;
    wire _T_707_2;
    wire _T_707_3;
    wire _T_707_4;
    wire _T_707_5;
    wire _T_707_6;
    wire _T_707_7;
    wire _T_707_8;
    wire _T_707_9;
    wire _T_707_10;
    wire _T_707_11;
    wire _T_707_12;
    wire _T_707_13;
    wire _T_707_14;
    wire _T_707_15;
    wire _T_707_16;
    wire _T_707_17;
    wire _T_707_18;
    wire _T_707_19;
    wire _T_707_20;
    wire _T_707_21;
    wire _T_707_22;
    wire _T_707_23;
    wire _T_707_24;
    wire _T_707_25;
    wire _T_707_26;
    wire _T_707_27;
    wire _T_707_28;
    wire _T_707_29;
    wire _T_707_30;
    wire _T_707_31;
    wire _T_707_32;
    wire _T_707_33;
    wire _T_707_34;
    wire _T_707_35;
    wire _T_707_36;
    wire _T_707_37;
    wire _T_707_38;
    wire _T_707_39;
    wire _T_707_40;
    wire _T_707_41;
    wire _T_707_42;
    wire _T_707_43;
    wire _T_707_44;
    wire _T_707_45;
    wire _T_707_46;
    wire _T_707_47;
    wire _T_707_48;
    wire _T_707_49;
    wire _T_707_50;
    wire _T_707_51;
    wire _T_707_52;
    wire [5:0] _value_3__q;
    wire [5:0] _value_3__d;
    DFF_POSCLK #(.width(6)) value_3 (
        .q(_value_3__q),
        .d(_value_3__d),
        .clk(clock)
    );
    wire [5:0] _WTEMP_25;
    MUX_UNSIGNED #(.width(6)) u_mux_693 (
        .y(_value_3__d),
        .sel(reset),
        .a(6'h0),
        .b(_WTEMP_25)
    );
    wire [30:0] _T_773_0;
    wire [30:0] _T_773_1;
    wire [30:0] _T_773_2;
    wire [30:0] _T_773_3;
    wire [30:0] _T_773_4;
    wire [30:0] _T_773_5;
    wire [5:0] _T_783;
    BITS #(.width(8), .high(5), .low(0)) bits_694 (
        .y(_T_783),
        .in(__T_10__q)
    );
    wire _node_645;
    EQ_UNSIGNED #(.width(6)) u_eq_695 (
        .y(_node_645),
        .a(6'd0),
        .b(_T_783)
    );
    wire _node_646;
    assign _node_646 = _T_707_0;
    wire _node_647;
    EQ_UNSIGNED #(.width(6)) u_eq_696 (
        .y(_node_647),
        .a(6'd1),
        .b(_T_783)
    );
    wire _node_648;
    MUX_UNSIGNED #(.width(1)) u_mux_697 (
        .y(_node_648),
        .sel(_node_647),
        .a(_T_707_1),
        .b(_node_646)
    );
    wire _node_649;
    EQ_UNSIGNED #(.width(6)) u_eq_698 (
        .y(_node_649),
        .a(6'd2),
        .b(_T_783)
    );
    wire _node_650;
    MUX_UNSIGNED #(.width(1)) u_mux_699 (
        .y(_node_650),
        .sel(_node_649),
        .a(_T_707_2),
        .b(_node_648)
    );
    wire _node_651;
    EQ_UNSIGNED #(.width(6)) u_eq_700 (
        .y(_node_651),
        .a(6'd3),
        .b(_T_783)
    );
    wire _node_652;
    MUX_UNSIGNED #(.width(1)) u_mux_701 (
        .y(_node_652),
        .sel(_node_651),
        .a(_T_707_3),
        .b(_node_650)
    );
    wire _node_653;
    EQ_UNSIGNED #(.width(6)) u_eq_702 (
        .y(_node_653),
        .a(6'd4),
        .b(_T_783)
    );
    wire _node_654;
    MUX_UNSIGNED #(.width(1)) u_mux_703 (
        .y(_node_654),
        .sel(_node_653),
        .a(_T_707_4),
        .b(_node_652)
    );
    wire _node_655;
    EQ_UNSIGNED #(.width(6)) u_eq_704 (
        .y(_node_655),
        .a(6'd5),
        .b(_T_783)
    );
    wire _node_656;
    MUX_UNSIGNED #(.width(1)) u_mux_705 (
        .y(_node_656),
        .sel(_node_655),
        .a(_T_707_5),
        .b(_node_654)
    );
    wire _node_657;
    EQ_UNSIGNED #(.width(6)) u_eq_706 (
        .y(_node_657),
        .a(6'd6),
        .b(_T_783)
    );
    wire _node_658;
    MUX_UNSIGNED #(.width(1)) u_mux_707 (
        .y(_node_658),
        .sel(_node_657),
        .a(_T_707_6),
        .b(_node_656)
    );
    wire _node_659;
    EQ_UNSIGNED #(.width(6)) u_eq_708 (
        .y(_node_659),
        .a(6'd7),
        .b(_T_783)
    );
    wire _node_660;
    MUX_UNSIGNED #(.width(1)) u_mux_709 (
        .y(_node_660),
        .sel(_node_659),
        .a(_T_707_7),
        .b(_node_658)
    );
    wire _node_661;
    EQ_UNSIGNED #(.width(6)) u_eq_710 (
        .y(_node_661),
        .a(6'd8),
        .b(_T_783)
    );
    wire _node_662;
    MUX_UNSIGNED #(.width(1)) u_mux_711 (
        .y(_node_662),
        .sel(_node_661),
        .a(_T_707_8),
        .b(_node_660)
    );
    wire _node_663;
    EQ_UNSIGNED #(.width(6)) u_eq_712 (
        .y(_node_663),
        .a(6'd9),
        .b(_T_783)
    );
    wire _node_664;
    MUX_UNSIGNED #(.width(1)) u_mux_713 (
        .y(_node_664),
        .sel(_node_663),
        .a(_T_707_9),
        .b(_node_662)
    );
    wire _node_665;
    EQ_UNSIGNED #(.width(6)) u_eq_714 (
        .y(_node_665),
        .a(6'd10),
        .b(_T_783)
    );
    wire _node_666;
    MUX_UNSIGNED #(.width(1)) u_mux_715 (
        .y(_node_666),
        .sel(_node_665),
        .a(_T_707_10),
        .b(_node_664)
    );
    wire _node_667;
    EQ_UNSIGNED #(.width(6)) u_eq_716 (
        .y(_node_667),
        .a(6'd11),
        .b(_T_783)
    );
    wire _node_668;
    MUX_UNSIGNED #(.width(1)) u_mux_717 (
        .y(_node_668),
        .sel(_node_667),
        .a(_T_707_11),
        .b(_node_666)
    );
    wire _node_669;
    EQ_UNSIGNED #(.width(6)) u_eq_718 (
        .y(_node_669),
        .a(6'd12),
        .b(_T_783)
    );
    wire _node_670;
    MUX_UNSIGNED #(.width(1)) u_mux_719 (
        .y(_node_670),
        .sel(_node_669),
        .a(_T_707_12),
        .b(_node_668)
    );
    wire _node_671;
    EQ_UNSIGNED #(.width(6)) u_eq_720 (
        .y(_node_671),
        .a(6'd13),
        .b(_T_783)
    );
    wire _node_672;
    MUX_UNSIGNED #(.width(1)) u_mux_721 (
        .y(_node_672),
        .sel(_node_671),
        .a(_T_707_13),
        .b(_node_670)
    );
    wire _node_673;
    EQ_UNSIGNED #(.width(6)) u_eq_722 (
        .y(_node_673),
        .a(6'd14),
        .b(_T_783)
    );
    wire _node_674;
    MUX_UNSIGNED #(.width(1)) u_mux_723 (
        .y(_node_674),
        .sel(_node_673),
        .a(_T_707_14),
        .b(_node_672)
    );
    wire _node_675;
    EQ_UNSIGNED #(.width(6)) u_eq_724 (
        .y(_node_675),
        .a(6'd15),
        .b(_T_783)
    );
    wire _node_676;
    MUX_UNSIGNED #(.width(1)) u_mux_725 (
        .y(_node_676),
        .sel(_node_675),
        .a(_T_707_15),
        .b(_node_674)
    );
    wire _node_677;
    EQ_UNSIGNED #(.width(6)) u_eq_726 (
        .y(_node_677),
        .a(6'd16),
        .b(_T_783)
    );
    wire _node_678;
    MUX_UNSIGNED #(.width(1)) u_mux_727 (
        .y(_node_678),
        .sel(_node_677),
        .a(_T_707_16),
        .b(_node_676)
    );
    wire _node_679;
    EQ_UNSIGNED #(.width(6)) u_eq_728 (
        .y(_node_679),
        .a(6'd17),
        .b(_T_783)
    );
    wire _node_680;
    MUX_UNSIGNED #(.width(1)) u_mux_729 (
        .y(_node_680),
        .sel(_node_679),
        .a(_T_707_17),
        .b(_node_678)
    );
    wire _node_681;
    EQ_UNSIGNED #(.width(6)) u_eq_730 (
        .y(_node_681),
        .a(6'd18),
        .b(_T_783)
    );
    wire _node_682;
    MUX_UNSIGNED #(.width(1)) u_mux_731 (
        .y(_node_682),
        .sel(_node_681),
        .a(_T_707_18),
        .b(_node_680)
    );
    wire _node_683;
    EQ_UNSIGNED #(.width(6)) u_eq_732 (
        .y(_node_683),
        .a(6'd19),
        .b(_T_783)
    );
    wire _node_684;
    MUX_UNSIGNED #(.width(1)) u_mux_733 (
        .y(_node_684),
        .sel(_node_683),
        .a(_T_707_19),
        .b(_node_682)
    );
    wire _node_685;
    EQ_UNSIGNED #(.width(6)) u_eq_734 (
        .y(_node_685),
        .a(6'd20),
        .b(_T_783)
    );
    wire _node_686;
    MUX_UNSIGNED #(.width(1)) u_mux_735 (
        .y(_node_686),
        .sel(_node_685),
        .a(_T_707_20),
        .b(_node_684)
    );
    wire _node_687;
    EQ_UNSIGNED #(.width(6)) u_eq_736 (
        .y(_node_687),
        .a(6'd21),
        .b(_T_783)
    );
    wire _node_688;
    MUX_UNSIGNED #(.width(1)) u_mux_737 (
        .y(_node_688),
        .sel(_node_687),
        .a(_T_707_21),
        .b(_node_686)
    );
    wire _node_689;
    EQ_UNSIGNED #(.width(6)) u_eq_738 (
        .y(_node_689),
        .a(6'd22),
        .b(_T_783)
    );
    wire _node_690;
    MUX_UNSIGNED #(.width(1)) u_mux_739 (
        .y(_node_690),
        .sel(_node_689),
        .a(_T_707_22),
        .b(_node_688)
    );
    wire _node_691;
    EQ_UNSIGNED #(.width(6)) u_eq_740 (
        .y(_node_691),
        .a(6'd23),
        .b(_T_783)
    );
    wire _node_692;
    MUX_UNSIGNED #(.width(1)) u_mux_741 (
        .y(_node_692),
        .sel(_node_691),
        .a(_T_707_23),
        .b(_node_690)
    );
    wire _node_693;
    EQ_UNSIGNED #(.width(6)) u_eq_742 (
        .y(_node_693),
        .a(6'd24),
        .b(_T_783)
    );
    wire _node_694;
    MUX_UNSIGNED #(.width(1)) u_mux_743 (
        .y(_node_694),
        .sel(_node_693),
        .a(_T_707_24),
        .b(_node_692)
    );
    wire _node_695;
    EQ_UNSIGNED #(.width(6)) u_eq_744 (
        .y(_node_695),
        .a(6'd25),
        .b(_T_783)
    );
    wire _node_696;
    MUX_UNSIGNED #(.width(1)) u_mux_745 (
        .y(_node_696),
        .sel(_node_695),
        .a(_T_707_25),
        .b(_node_694)
    );
    wire _node_697;
    EQ_UNSIGNED #(.width(6)) u_eq_746 (
        .y(_node_697),
        .a(6'd26),
        .b(_T_783)
    );
    wire _node_698;
    MUX_UNSIGNED #(.width(1)) u_mux_747 (
        .y(_node_698),
        .sel(_node_697),
        .a(_T_707_26),
        .b(_node_696)
    );
    wire _node_699;
    EQ_UNSIGNED #(.width(6)) u_eq_748 (
        .y(_node_699),
        .a(6'd27),
        .b(_T_783)
    );
    wire _node_700;
    MUX_UNSIGNED #(.width(1)) u_mux_749 (
        .y(_node_700),
        .sel(_node_699),
        .a(_T_707_27),
        .b(_node_698)
    );
    wire _node_701;
    EQ_UNSIGNED #(.width(6)) u_eq_750 (
        .y(_node_701),
        .a(6'd28),
        .b(_T_783)
    );
    wire _node_702;
    MUX_UNSIGNED #(.width(1)) u_mux_751 (
        .y(_node_702),
        .sel(_node_701),
        .a(_T_707_28),
        .b(_node_700)
    );
    wire _node_703;
    EQ_UNSIGNED #(.width(6)) u_eq_752 (
        .y(_node_703),
        .a(6'd29),
        .b(_T_783)
    );
    wire _node_704;
    MUX_UNSIGNED #(.width(1)) u_mux_753 (
        .y(_node_704),
        .sel(_node_703),
        .a(_T_707_29),
        .b(_node_702)
    );
    wire _node_705;
    EQ_UNSIGNED #(.width(6)) u_eq_754 (
        .y(_node_705),
        .a(6'd30),
        .b(_T_783)
    );
    wire _node_706;
    MUX_UNSIGNED #(.width(1)) u_mux_755 (
        .y(_node_706),
        .sel(_node_705),
        .a(_T_707_30),
        .b(_node_704)
    );
    wire _node_707;
    EQ_UNSIGNED #(.width(6)) u_eq_756 (
        .y(_node_707),
        .a(6'd31),
        .b(_T_783)
    );
    wire _node_708;
    MUX_UNSIGNED #(.width(1)) u_mux_757 (
        .y(_node_708),
        .sel(_node_707),
        .a(_T_707_31),
        .b(_node_706)
    );
    wire _node_709;
    EQ_UNSIGNED #(.width(6)) u_eq_758 (
        .y(_node_709),
        .a(6'd32),
        .b(_T_783)
    );
    wire _node_710;
    MUX_UNSIGNED #(.width(1)) u_mux_759 (
        .y(_node_710),
        .sel(_node_709),
        .a(_T_707_32),
        .b(_node_708)
    );
    wire _node_711;
    EQ_UNSIGNED #(.width(6)) u_eq_760 (
        .y(_node_711),
        .a(6'd33),
        .b(_T_783)
    );
    wire _node_712;
    MUX_UNSIGNED #(.width(1)) u_mux_761 (
        .y(_node_712),
        .sel(_node_711),
        .a(_T_707_33),
        .b(_node_710)
    );
    wire _node_713;
    EQ_UNSIGNED #(.width(6)) u_eq_762 (
        .y(_node_713),
        .a(6'd34),
        .b(_T_783)
    );
    wire _node_714;
    MUX_UNSIGNED #(.width(1)) u_mux_763 (
        .y(_node_714),
        .sel(_node_713),
        .a(_T_707_34),
        .b(_node_712)
    );
    wire _node_715;
    EQ_UNSIGNED #(.width(6)) u_eq_764 (
        .y(_node_715),
        .a(6'd35),
        .b(_T_783)
    );
    wire _node_716;
    MUX_UNSIGNED #(.width(1)) u_mux_765 (
        .y(_node_716),
        .sel(_node_715),
        .a(_T_707_35),
        .b(_node_714)
    );
    wire _node_717;
    EQ_UNSIGNED #(.width(6)) u_eq_766 (
        .y(_node_717),
        .a(6'd36),
        .b(_T_783)
    );
    wire _node_718;
    MUX_UNSIGNED #(.width(1)) u_mux_767 (
        .y(_node_718),
        .sel(_node_717),
        .a(_T_707_36),
        .b(_node_716)
    );
    wire _node_719;
    EQ_UNSIGNED #(.width(6)) u_eq_768 (
        .y(_node_719),
        .a(6'd37),
        .b(_T_783)
    );
    wire _node_720;
    MUX_UNSIGNED #(.width(1)) u_mux_769 (
        .y(_node_720),
        .sel(_node_719),
        .a(_T_707_37),
        .b(_node_718)
    );
    wire _node_721;
    EQ_UNSIGNED #(.width(6)) u_eq_770 (
        .y(_node_721),
        .a(6'd38),
        .b(_T_783)
    );
    wire _node_722;
    MUX_UNSIGNED #(.width(1)) u_mux_771 (
        .y(_node_722),
        .sel(_node_721),
        .a(_T_707_38),
        .b(_node_720)
    );
    wire _node_723;
    EQ_UNSIGNED #(.width(6)) u_eq_772 (
        .y(_node_723),
        .a(6'd39),
        .b(_T_783)
    );
    wire _node_724;
    MUX_UNSIGNED #(.width(1)) u_mux_773 (
        .y(_node_724),
        .sel(_node_723),
        .a(_T_707_39),
        .b(_node_722)
    );
    wire _node_725;
    EQ_UNSIGNED #(.width(6)) u_eq_774 (
        .y(_node_725),
        .a(6'd40),
        .b(_T_783)
    );
    wire _node_726;
    MUX_UNSIGNED #(.width(1)) u_mux_775 (
        .y(_node_726),
        .sel(_node_725),
        .a(_T_707_40),
        .b(_node_724)
    );
    wire _node_727;
    EQ_UNSIGNED #(.width(6)) u_eq_776 (
        .y(_node_727),
        .a(6'd41),
        .b(_T_783)
    );
    wire _node_728;
    MUX_UNSIGNED #(.width(1)) u_mux_777 (
        .y(_node_728),
        .sel(_node_727),
        .a(_T_707_41),
        .b(_node_726)
    );
    wire _node_729;
    EQ_UNSIGNED #(.width(6)) u_eq_778 (
        .y(_node_729),
        .a(6'd42),
        .b(_T_783)
    );
    wire _node_730;
    MUX_UNSIGNED #(.width(1)) u_mux_779 (
        .y(_node_730),
        .sel(_node_729),
        .a(_T_707_42),
        .b(_node_728)
    );
    wire _node_731;
    EQ_UNSIGNED #(.width(6)) u_eq_780 (
        .y(_node_731),
        .a(6'd43),
        .b(_T_783)
    );
    wire _node_732;
    MUX_UNSIGNED #(.width(1)) u_mux_781 (
        .y(_node_732),
        .sel(_node_731),
        .a(_T_707_43),
        .b(_node_730)
    );
    wire _node_733;
    EQ_UNSIGNED #(.width(6)) u_eq_782 (
        .y(_node_733),
        .a(6'd44),
        .b(_T_783)
    );
    wire _node_734;
    MUX_UNSIGNED #(.width(1)) u_mux_783 (
        .y(_node_734),
        .sel(_node_733),
        .a(_T_707_44),
        .b(_node_732)
    );
    wire _node_735;
    EQ_UNSIGNED #(.width(6)) u_eq_784 (
        .y(_node_735),
        .a(6'd45),
        .b(_T_783)
    );
    wire _node_736;
    MUX_UNSIGNED #(.width(1)) u_mux_785 (
        .y(_node_736),
        .sel(_node_735),
        .a(_T_707_45),
        .b(_node_734)
    );
    wire _node_737;
    EQ_UNSIGNED #(.width(6)) u_eq_786 (
        .y(_node_737),
        .a(6'd46),
        .b(_T_783)
    );
    wire _node_738;
    MUX_UNSIGNED #(.width(1)) u_mux_787 (
        .y(_node_738),
        .sel(_node_737),
        .a(_T_707_46),
        .b(_node_736)
    );
    wire _node_739;
    EQ_UNSIGNED #(.width(6)) u_eq_788 (
        .y(_node_739),
        .a(6'd47),
        .b(_T_783)
    );
    wire _node_740;
    MUX_UNSIGNED #(.width(1)) u_mux_789 (
        .y(_node_740),
        .sel(_node_739),
        .a(_T_707_47),
        .b(_node_738)
    );
    wire _node_741;
    EQ_UNSIGNED #(.width(6)) u_eq_790 (
        .y(_node_741),
        .a(6'd48),
        .b(_T_783)
    );
    wire _node_742;
    MUX_UNSIGNED #(.width(1)) u_mux_791 (
        .y(_node_742),
        .sel(_node_741),
        .a(_T_707_48),
        .b(_node_740)
    );
    wire _node_743;
    EQ_UNSIGNED #(.width(6)) u_eq_792 (
        .y(_node_743),
        .a(6'd49),
        .b(_T_783)
    );
    wire _node_744;
    MUX_UNSIGNED #(.width(1)) u_mux_793 (
        .y(_node_744),
        .sel(_node_743),
        .a(_T_707_49),
        .b(_node_742)
    );
    wire _node_745;
    EQ_UNSIGNED #(.width(6)) u_eq_794 (
        .y(_node_745),
        .a(6'd50),
        .b(_T_783)
    );
    wire _node_746;
    MUX_UNSIGNED #(.width(1)) u_mux_795 (
        .y(_node_746),
        .sel(_node_745),
        .a(_T_707_50),
        .b(_node_744)
    );
    wire _node_747;
    EQ_UNSIGNED #(.width(6)) u_eq_796 (
        .y(_node_747),
        .a(6'd51),
        .b(_T_783)
    );
    wire _node_748;
    MUX_UNSIGNED #(.width(1)) u_mux_797 (
        .y(_node_748),
        .sel(_node_747),
        .a(_T_707_51),
        .b(_node_746)
    );
    wire _node_749;
    EQ_UNSIGNED #(.width(6)) u_eq_798 (
        .y(_node_749),
        .a(6'd52),
        .b(_T_783)
    );
    wire _node_750;
    MUX_UNSIGNED #(.width(1)) u_mux_799 (
        .y(_node_750),
        .sel(_node_749),
        .a(_T_707_52),
        .b(_node_748)
    );
    wire _T_784;
    BITWISEAND #(.width(1)) bitwiseand_800 (
        .y(_T_784),
        .a(_c__io_outs_1_ready),
        .b(_c__io_outs_1_valid)
    );
    wire [2:0] _T_786;
    BITS #(.width(6), .high(2), .low(0)) bits_801 (
        .y(_T_786),
        .in(_value_3__q)
    );
    wire _T_788;
    EQ_UNSIGNED #(.width(1)) u_eq_802 (
        .y(_T_788),
        .a(reset),
        .b(1'h0)
    );
    wire [2:0] _T_790;
    BITS #(.width(6), .high(2), .low(0)) bits_803 (
        .y(_T_790),
        .in(_value_3__q)
    );
    wire _node_751;
    EQ_UNSIGNED #(.width(3)) u_eq_804 (
        .y(_node_751),
        .a(3'd0),
        .b(_T_790)
    );
    wire [30:0] _node_752;
    assign _node_752 = _T_773_0;
    wire _node_753;
    EQ_UNSIGNED #(.width(3)) u_eq_805 (
        .y(_node_753),
        .a(3'd1),
        .b(_T_790)
    );
    wire [30:0] _node_754;
    MUX_UNSIGNED #(.width(31)) u_mux_806 (
        .y(_node_754),
        .sel(_node_753),
        .a(_T_773_1),
        .b(_node_752)
    );
    wire _node_755;
    EQ_UNSIGNED #(.width(3)) u_eq_807 (
        .y(_node_755),
        .a(3'd2),
        .b(_T_790)
    );
    wire [30:0] _node_756;
    MUX_UNSIGNED #(.width(31)) u_mux_808 (
        .y(_node_756),
        .sel(_node_755),
        .a(_T_773_2),
        .b(_node_754)
    );
    wire _node_757;
    EQ_UNSIGNED #(.width(3)) u_eq_809 (
        .y(_node_757),
        .a(3'd3),
        .b(_T_790)
    );
    wire [30:0] _node_758;
    MUX_UNSIGNED #(.width(31)) u_mux_810 (
        .y(_node_758),
        .sel(_node_757),
        .a(_T_773_3),
        .b(_node_756)
    );
    wire _node_759;
    EQ_UNSIGNED #(.width(3)) u_eq_811 (
        .y(_node_759),
        .a(3'd4),
        .b(_T_790)
    );
    wire [30:0] _node_760;
    MUX_UNSIGNED #(.width(31)) u_mux_812 (
        .y(_node_760),
        .sel(_node_759),
        .a(_T_773_4),
        .b(_node_758)
    );
    wire _node_761;
    EQ_UNSIGNED #(.width(3)) u_eq_813 (
        .y(_node_761),
        .a(3'd5),
        .b(_T_790)
    );
    wire [30:0] _node_762;
    MUX_UNSIGNED #(.width(31)) u_mux_814 (
        .y(_node_762),
        .sel(_node_761),
        .a(_T_773_5),
        .b(_node_760)
    );
    wire _T_791;
    wire [63:0] _WTEMP_26;
    PAD_UNSIGNED #(.width(31), .n(64)) u_pad_815 (
        .y(_WTEMP_26),
        .in(_node_762)
    );
    NEQ_UNSIGNED #(.width(64)) u_neq_816 (
        .y(_T_791),
        .a(_c__io_outs_1_bits_body),
        .b(_WTEMP_26)
    );
    wire [2:0] _T_793;
    BITS #(.width(6), .high(2), .low(0)) bits_817 (
        .y(_T_793),
        .in(_value_3__q)
    );
    wire _T_795;
    EQ_UNSIGNED #(.width(1)) u_eq_818 (
        .y(_T_795),
        .a(reset),
        .b(1'h0)
    );
    wire _T_797;
    BITWISEOR #(.width(1)) bitwiseor_819 (
        .y(_T_797),
        .a(1'h0),
        .b(reset)
    );
    wire _T_799;
    EQ_UNSIGNED #(.width(1)) u_eq_820 (
        .y(_T_799),
        .a(_T_797),
        .b(1'h0)
    );
    wire _T_801;
    EQ_UNSIGNED #(.width(1)) u_eq_821 (
        .y(_T_801),
        .a(reset),
        .b(1'h0)
    );
    wire _T_803;
    EQ_UNSIGNED #(.width(6)) u_eq_822 (
        .y(_T_803),
        .a(_value_3__q),
        .b(6'h20)
    );
    wire [6:0] _T_805;
    wire [5:0] _WTEMP_27;
    PAD_UNSIGNED #(.width(1), .n(6)) u_pad_823 (
        .y(_WTEMP_27),
        .in(1'h1)
    );
    ADD_UNSIGNED #(.width(6)) u_add_824 (
        .y(_T_805),
        .a(_value_3__q),
        .b(_WTEMP_27)
    );
    wire [5:0] _T_806;
    TAIL #(.width(7), .n(1)) tail_825 (
        .y(_T_806),
        .in(_T_805)
    );
    wire _T_809;
    EQ_UNSIGNED #(.width(1)) u_eq_826 (
        .y(_T_809),
        .a(__T_13__q),
        .b(1'h0)
    );
    wire _T_811;
    wire [7:0] _WTEMP_28;
    PAD_UNSIGNED #(.width(6), .n(8)) u_pad_827 (
        .y(_WTEMP_28),
        .in(6'h20)
    );
    EQ_UNSIGNED #(.width(8)) u_eq_828 (
        .y(_T_811),
        .a(__T_10__q),
        .b(_WTEMP_28)
    );
    wire [8:0] _T_814;
    wire [7:0] _WTEMP_29;
    PAD_UNSIGNED #(.width(1), .n(8)) u_pad_829 (
        .y(_WTEMP_29),
        .in(1'h1)
    );
    ADD_UNSIGNED #(.width(8)) u_add_830 (
        .y(_T_814),
        .a(__T_10__q),
        .b(_WTEMP_29)
    );
    wire [7:0] _T_815;
    TAIL #(.width(9), .n(1)) tail_831 (
        .y(_T_815),
        .in(_T_814)
    );
    wire _node_763;
    MUX_UNSIGNED #(.width(1)) u_mux_832 (
        .y(_node_763),
        .sel(_T_811),
        .a(1'h1),
        .b(__T_13__q)
    );
    wire [7:0] _node_764;
    MUX_UNSIGNED #(.width(8)) u_mux_833 (
        .y(_node_764),
        .sel(_T_809),
        .a(_T_815),
        .b(__T_10__q)
    );
    wire _node_765;
    MUX_UNSIGNED #(.width(1)) u_mux_834 (
        .y(_node_765),
        .sel(_T_809),
        .a(_node_763),
        .b(__T_13__q)
    );
    wire [5:0] _node_766;
    wire [5:0] _WTEMP_30;
    PAD_UNSIGNED #(.width(1), .n(6)) u_pad_835 (
        .y(_WTEMP_30),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(6)) u_mux_836 (
        .y(_node_766),
        .sel(_T_803),
        .a(_WTEMP_30),
        .b(_T_806)
    );
    wire _T_871_0;
    wire _T_871_1;
    wire _T_871_2;
    wire _T_871_3;
    wire _T_871_4;
    wire _T_871_5;
    wire _T_871_6;
    wire _T_871_7;
    wire _T_871_8;
    wire _T_871_9;
    wire _T_871_10;
    wire _T_871_11;
    wire _T_871_12;
    wire _T_871_13;
    wire _T_871_14;
    wire _T_871_15;
    wire _T_871_16;
    wire _T_871_17;
    wire _T_871_18;
    wire _T_871_19;
    wire _T_871_20;
    wire _T_871_21;
    wire _T_871_22;
    wire _T_871_23;
    wire _T_871_24;
    wire _T_871_25;
    wire _T_871_26;
    wire _T_871_27;
    wire _T_871_28;
    wire _T_871_29;
    wire _T_871_30;
    wire _T_871_31;
    wire _T_871_32;
    wire _T_871_33;
    wire _T_871_34;
    wire _T_871_35;
    wire _T_871_36;
    wire _T_871_37;
    wire _T_871_38;
    wire _T_871_39;
    wire _T_871_40;
    wire _T_871_41;
    wire _T_871_42;
    wire _T_871_43;
    wire _T_871_44;
    wire _T_871_45;
    wire _T_871_46;
    wire _T_871_47;
    wire _T_871_48;
    wire _T_871_49;
    wire _T_871_50;
    wire _T_871_51;
    wire _T_871_52;
    wire [5:0] _value_4__q;
    wire [5:0] _value_4__d;
    DFF_POSCLK #(.width(6)) value_4 (
        .q(_value_4__q),
        .d(_value_4__d),
        .clk(clock)
    );
    wire [5:0] _WTEMP_31;
    MUX_UNSIGNED #(.width(6)) u_mux_837 (
        .y(_value_4__d),
        .sel(reset),
        .a(6'h0),
        .b(_WTEMP_31)
    );
    wire [30:0] _T_942_0;
    wire [30:0] _T_942_1;
    wire [30:0] _T_942_2;
    wire [30:0] _T_942_3;
    wire [30:0] _T_942_4;
    wire [30:0] _T_942_5;
    wire [30:0] _T_942_6;
    wire [30:0] _T_942_7;
    wire [30:0] _T_942_8;
    wire [30:0] _T_942_9;
    wire [30:0] _T_942_10;
    wire [5:0] _T_957;
    BITS #(.width(8), .high(5), .low(0)) bits_838 (
        .y(_T_957),
        .in(__T_10__q)
    );
    wire _node_767;
    EQ_UNSIGNED #(.width(6)) u_eq_839 (
        .y(_node_767),
        .a(6'd0),
        .b(_T_957)
    );
    wire _node_768;
    assign _node_768 = _T_871_0;
    wire _node_769;
    EQ_UNSIGNED #(.width(6)) u_eq_840 (
        .y(_node_769),
        .a(6'd1),
        .b(_T_957)
    );
    wire _node_770;
    MUX_UNSIGNED #(.width(1)) u_mux_841 (
        .y(_node_770),
        .sel(_node_769),
        .a(_T_871_1),
        .b(_node_768)
    );
    wire _node_771;
    EQ_UNSIGNED #(.width(6)) u_eq_842 (
        .y(_node_771),
        .a(6'd2),
        .b(_T_957)
    );
    wire _node_772;
    MUX_UNSIGNED #(.width(1)) u_mux_843 (
        .y(_node_772),
        .sel(_node_771),
        .a(_T_871_2),
        .b(_node_770)
    );
    wire _node_773;
    EQ_UNSIGNED #(.width(6)) u_eq_844 (
        .y(_node_773),
        .a(6'd3),
        .b(_T_957)
    );
    wire _node_774;
    MUX_UNSIGNED #(.width(1)) u_mux_845 (
        .y(_node_774),
        .sel(_node_773),
        .a(_T_871_3),
        .b(_node_772)
    );
    wire _node_775;
    EQ_UNSIGNED #(.width(6)) u_eq_846 (
        .y(_node_775),
        .a(6'd4),
        .b(_T_957)
    );
    wire _node_776;
    MUX_UNSIGNED #(.width(1)) u_mux_847 (
        .y(_node_776),
        .sel(_node_775),
        .a(_T_871_4),
        .b(_node_774)
    );
    wire _node_777;
    EQ_UNSIGNED #(.width(6)) u_eq_848 (
        .y(_node_777),
        .a(6'd5),
        .b(_T_957)
    );
    wire _node_778;
    MUX_UNSIGNED #(.width(1)) u_mux_849 (
        .y(_node_778),
        .sel(_node_777),
        .a(_T_871_5),
        .b(_node_776)
    );
    wire _node_779;
    EQ_UNSIGNED #(.width(6)) u_eq_850 (
        .y(_node_779),
        .a(6'd6),
        .b(_T_957)
    );
    wire _node_780;
    MUX_UNSIGNED #(.width(1)) u_mux_851 (
        .y(_node_780),
        .sel(_node_779),
        .a(_T_871_6),
        .b(_node_778)
    );
    wire _node_781;
    EQ_UNSIGNED #(.width(6)) u_eq_852 (
        .y(_node_781),
        .a(6'd7),
        .b(_T_957)
    );
    wire _node_782;
    MUX_UNSIGNED #(.width(1)) u_mux_853 (
        .y(_node_782),
        .sel(_node_781),
        .a(_T_871_7),
        .b(_node_780)
    );
    wire _node_783;
    EQ_UNSIGNED #(.width(6)) u_eq_854 (
        .y(_node_783),
        .a(6'd8),
        .b(_T_957)
    );
    wire _node_784;
    MUX_UNSIGNED #(.width(1)) u_mux_855 (
        .y(_node_784),
        .sel(_node_783),
        .a(_T_871_8),
        .b(_node_782)
    );
    wire _node_785;
    EQ_UNSIGNED #(.width(6)) u_eq_856 (
        .y(_node_785),
        .a(6'd9),
        .b(_T_957)
    );
    wire _node_786;
    MUX_UNSIGNED #(.width(1)) u_mux_857 (
        .y(_node_786),
        .sel(_node_785),
        .a(_T_871_9),
        .b(_node_784)
    );
    wire _node_787;
    EQ_UNSIGNED #(.width(6)) u_eq_858 (
        .y(_node_787),
        .a(6'd10),
        .b(_T_957)
    );
    wire _node_788;
    MUX_UNSIGNED #(.width(1)) u_mux_859 (
        .y(_node_788),
        .sel(_node_787),
        .a(_T_871_10),
        .b(_node_786)
    );
    wire _node_789;
    EQ_UNSIGNED #(.width(6)) u_eq_860 (
        .y(_node_789),
        .a(6'd11),
        .b(_T_957)
    );
    wire _node_790;
    MUX_UNSIGNED #(.width(1)) u_mux_861 (
        .y(_node_790),
        .sel(_node_789),
        .a(_T_871_11),
        .b(_node_788)
    );
    wire _node_791;
    EQ_UNSIGNED #(.width(6)) u_eq_862 (
        .y(_node_791),
        .a(6'd12),
        .b(_T_957)
    );
    wire _node_792;
    MUX_UNSIGNED #(.width(1)) u_mux_863 (
        .y(_node_792),
        .sel(_node_791),
        .a(_T_871_12),
        .b(_node_790)
    );
    wire _node_793;
    EQ_UNSIGNED #(.width(6)) u_eq_864 (
        .y(_node_793),
        .a(6'd13),
        .b(_T_957)
    );
    wire _node_794;
    MUX_UNSIGNED #(.width(1)) u_mux_865 (
        .y(_node_794),
        .sel(_node_793),
        .a(_T_871_13),
        .b(_node_792)
    );
    wire _node_795;
    EQ_UNSIGNED #(.width(6)) u_eq_866 (
        .y(_node_795),
        .a(6'd14),
        .b(_T_957)
    );
    wire _node_796;
    MUX_UNSIGNED #(.width(1)) u_mux_867 (
        .y(_node_796),
        .sel(_node_795),
        .a(_T_871_14),
        .b(_node_794)
    );
    wire _node_797;
    EQ_UNSIGNED #(.width(6)) u_eq_868 (
        .y(_node_797),
        .a(6'd15),
        .b(_T_957)
    );
    wire _node_798;
    MUX_UNSIGNED #(.width(1)) u_mux_869 (
        .y(_node_798),
        .sel(_node_797),
        .a(_T_871_15),
        .b(_node_796)
    );
    wire _node_799;
    EQ_UNSIGNED #(.width(6)) u_eq_870 (
        .y(_node_799),
        .a(6'd16),
        .b(_T_957)
    );
    wire _node_800;
    MUX_UNSIGNED #(.width(1)) u_mux_871 (
        .y(_node_800),
        .sel(_node_799),
        .a(_T_871_16),
        .b(_node_798)
    );
    wire _node_801;
    EQ_UNSIGNED #(.width(6)) u_eq_872 (
        .y(_node_801),
        .a(6'd17),
        .b(_T_957)
    );
    wire _node_802;
    MUX_UNSIGNED #(.width(1)) u_mux_873 (
        .y(_node_802),
        .sel(_node_801),
        .a(_T_871_17),
        .b(_node_800)
    );
    wire _node_803;
    EQ_UNSIGNED #(.width(6)) u_eq_874 (
        .y(_node_803),
        .a(6'd18),
        .b(_T_957)
    );
    wire _node_804;
    MUX_UNSIGNED #(.width(1)) u_mux_875 (
        .y(_node_804),
        .sel(_node_803),
        .a(_T_871_18),
        .b(_node_802)
    );
    wire _node_805;
    EQ_UNSIGNED #(.width(6)) u_eq_876 (
        .y(_node_805),
        .a(6'd19),
        .b(_T_957)
    );
    wire _node_806;
    MUX_UNSIGNED #(.width(1)) u_mux_877 (
        .y(_node_806),
        .sel(_node_805),
        .a(_T_871_19),
        .b(_node_804)
    );
    wire _node_807;
    EQ_UNSIGNED #(.width(6)) u_eq_878 (
        .y(_node_807),
        .a(6'd20),
        .b(_T_957)
    );
    wire _node_808;
    MUX_UNSIGNED #(.width(1)) u_mux_879 (
        .y(_node_808),
        .sel(_node_807),
        .a(_T_871_20),
        .b(_node_806)
    );
    wire _node_809;
    EQ_UNSIGNED #(.width(6)) u_eq_880 (
        .y(_node_809),
        .a(6'd21),
        .b(_T_957)
    );
    wire _node_810;
    MUX_UNSIGNED #(.width(1)) u_mux_881 (
        .y(_node_810),
        .sel(_node_809),
        .a(_T_871_21),
        .b(_node_808)
    );
    wire _node_811;
    EQ_UNSIGNED #(.width(6)) u_eq_882 (
        .y(_node_811),
        .a(6'd22),
        .b(_T_957)
    );
    wire _node_812;
    MUX_UNSIGNED #(.width(1)) u_mux_883 (
        .y(_node_812),
        .sel(_node_811),
        .a(_T_871_22),
        .b(_node_810)
    );
    wire _node_813;
    EQ_UNSIGNED #(.width(6)) u_eq_884 (
        .y(_node_813),
        .a(6'd23),
        .b(_T_957)
    );
    wire _node_814;
    MUX_UNSIGNED #(.width(1)) u_mux_885 (
        .y(_node_814),
        .sel(_node_813),
        .a(_T_871_23),
        .b(_node_812)
    );
    wire _node_815;
    EQ_UNSIGNED #(.width(6)) u_eq_886 (
        .y(_node_815),
        .a(6'd24),
        .b(_T_957)
    );
    wire _node_816;
    MUX_UNSIGNED #(.width(1)) u_mux_887 (
        .y(_node_816),
        .sel(_node_815),
        .a(_T_871_24),
        .b(_node_814)
    );
    wire _node_817;
    EQ_UNSIGNED #(.width(6)) u_eq_888 (
        .y(_node_817),
        .a(6'd25),
        .b(_T_957)
    );
    wire _node_818;
    MUX_UNSIGNED #(.width(1)) u_mux_889 (
        .y(_node_818),
        .sel(_node_817),
        .a(_T_871_25),
        .b(_node_816)
    );
    wire _node_819;
    EQ_UNSIGNED #(.width(6)) u_eq_890 (
        .y(_node_819),
        .a(6'd26),
        .b(_T_957)
    );
    wire _node_820;
    MUX_UNSIGNED #(.width(1)) u_mux_891 (
        .y(_node_820),
        .sel(_node_819),
        .a(_T_871_26),
        .b(_node_818)
    );
    wire _node_821;
    EQ_UNSIGNED #(.width(6)) u_eq_892 (
        .y(_node_821),
        .a(6'd27),
        .b(_T_957)
    );
    wire _node_822;
    MUX_UNSIGNED #(.width(1)) u_mux_893 (
        .y(_node_822),
        .sel(_node_821),
        .a(_T_871_27),
        .b(_node_820)
    );
    wire _node_823;
    EQ_UNSIGNED #(.width(6)) u_eq_894 (
        .y(_node_823),
        .a(6'd28),
        .b(_T_957)
    );
    wire _node_824;
    MUX_UNSIGNED #(.width(1)) u_mux_895 (
        .y(_node_824),
        .sel(_node_823),
        .a(_T_871_28),
        .b(_node_822)
    );
    wire _node_825;
    EQ_UNSIGNED #(.width(6)) u_eq_896 (
        .y(_node_825),
        .a(6'd29),
        .b(_T_957)
    );
    wire _node_826;
    MUX_UNSIGNED #(.width(1)) u_mux_897 (
        .y(_node_826),
        .sel(_node_825),
        .a(_T_871_29),
        .b(_node_824)
    );
    wire _node_827;
    EQ_UNSIGNED #(.width(6)) u_eq_898 (
        .y(_node_827),
        .a(6'd30),
        .b(_T_957)
    );
    wire _node_828;
    MUX_UNSIGNED #(.width(1)) u_mux_899 (
        .y(_node_828),
        .sel(_node_827),
        .a(_T_871_30),
        .b(_node_826)
    );
    wire _node_829;
    EQ_UNSIGNED #(.width(6)) u_eq_900 (
        .y(_node_829),
        .a(6'd31),
        .b(_T_957)
    );
    wire _node_830;
    MUX_UNSIGNED #(.width(1)) u_mux_901 (
        .y(_node_830),
        .sel(_node_829),
        .a(_T_871_31),
        .b(_node_828)
    );
    wire _node_831;
    EQ_UNSIGNED #(.width(6)) u_eq_902 (
        .y(_node_831),
        .a(6'd32),
        .b(_T_957)
    );
    wire _node_832;
    MUX_UNSIGNED #(.width(1)) u_mux_903 (
        .y(_node_832),
        .sel(_node_831),
        .a(_T_871_32),
        .b(_node_830)
    );
    wire _node_833;
    EQ_UNSIGNED #(.width(6)) u_eq_904 (
        .y(_node_833),
        .a(6'd33),
        .b(_T_957)
    );
    wire _node_834;
    MUX_UNSIGNED #(.width(1)) u_mux_905 (
        .y(_node_834),
        .sel(_node_833),
        .a(_T_871_33),
        .b(_node_832)
    );
    wire _node_835;
    EQ_UNSIGNED #(.width(6)) u_eq_906 (
        .y(_node_835),
        .a(6'd34),
        .b(_T_957)
    );
    wire _node_836;
    MUX_UNSIGNED #(.width(1)) u_mux_907 (
        .y(_node_836),
        .sel(_node_835),
        .a(_T_871_34),
        .b(_node_834)
    );
    wire _node_837;
    EQ_UNSIGNED #(.width(6)) u_eq_908 (
        .y(_node_837),
        .a(6'd35),
        .b(_T_957)
    );
    wire _node_838;
    MUX_UNSIGNED #(.width(1)) u_mux_909 (
        .y(_node_838),
        .sel(_node_837),
        .a(_T_871_35),
        .b(_node_836)
    );
    wire _node_839;
    EQ_UNSIGNED #(.width(6)) u_eq_910 (
        .y(_node_839),
        .a(6'd36),
        .b(_T_957)
    );
    wire _node_840;
    MUX_UNSIGNED #(.width(1)) u_mux_911 (
        .y(_node_840),
        .sel(_node_839),
        .a(_T_871_36),
        .b(_node_838)
    );
    wire _node_841;
    EQ_UNSIGNED #(.width(6)) u_eq_912 (
        .y(_node_841),
        .a(6'd37),
        .b(_T_957)
    );
    wire _node_842;
    MUX_UNSIGNED #(.width(1)) u_mux_913 (
        .y(_node_842),
        .sel(_node_841),
        .a(_T_871_37),
        .b(_node_840)
    );
    wire _node_843;
    EQ_UNSIGNED #(.width(6)) u_eq_914 (
        .y(_node_843),
        .a(6'd38),
        .b(_T_957)
    );
    wire _node_844;
    MUX_UNSIGNED #(.width(1)) u_mux_915 (
        .y(_node_844),
        .sel(_node_843),
        .a(_T_871_38),
        .b(_node_842)
    );
    wire _node_845;
    EQ_UNSIGNED #(.width(6)) u_eq_916 (
        .y(_node_845),
        .a(6'd39),
        .b(_T_957)
    );
    wire _node_846;
    MUX_UNSIGNED #(.width(1)) u_mux_917 (
        .y(_node_846),
        .sel(_node_845),
        .a(_T_871_39),
        .b(_node_844)
    );
    wire _node_847;
    EQ_UNSIGNED #(.width(6)) u_eq_918 (
        .y(_node_847),
        .a(6'd40),
        .b(_T_957)
    );
    wire _node_848;
    MUX_UNSIGNED #(.width(1)) u_mux_919 (
        .y(_node_848),
        .sel(_node_847),
        .a(_T_871_40),
        .b(_node_846)
    );
    wire _node_849;
    EQ_UNSIGNED #(.width(6)) u_eq_920 (
        .y(_node_849),
        .a(6'd41),
        .b(_T_957)
    );
    wire _node_850;
    MUX_UNSIGNED #(.width(1)) u_mux_921 (
        .y(_node_850),
        .sel(_node_849),
        .a(_T_871_41),
        .b(_node_848)
    );
    wire _node_851;
    EQ_UNSIGNED #(.width(6)) u_eq_922 (
        .y(_node_851),
        .a(6'd42),
        .b(_T_957)
    );
    wire _node_852;
    MUX_UNSIGNED #(.width(1)) u_mux_923 (
        .y(_node_852),
        .sel(_node_851),
        .a(_T_871_42),
        .b(_node_850)
    );
    wire _node_853;
    EQ_UNSIGNED #(.width(6)) u_eq_924 (
        .y(_node_853),
        .a(6'd43),
        .b(_T_957)
    );
    wire _node_854;
    MUX_UNSIGNED #(.width(1)) u_mux_925 (
        .y(_node_854),
        .sel(_node_853),
        .a(_T_871_43),
        .b(_node_852)
    );
    wire _node_855;
    EQ_UNSIGNED #(.width(6)) u_eq_926 (
        .y(_node_855),
        .a(6'd44),
        .b(_T_957)
    );
    wire _node_856;
    MUX_UNSIGNED #(.width(1)) u_mux_927 (
        .y(_node_856),
        .sel(_node_855),
        .a(_T_871_44),
        .b(_node_854)
    );
    wire _node_857;
    EQ_UNSIGNED #(.width(6)) u_eq_928 (
        .y(_node_857),
        .a(6'd45),
        .b(_T_957)
    );
    wire _node_858;
    MUX_UNSIGNED #(.width(1)) u_mux_929 (
        .y(_node_858),
        .sel(_node_857),
        .a(_T_871_45),
        .b(_node_856)
    );
    wire _node_859;
    EQ_UNSIGNED #(.width(6)) u_eq_930 (
        .y(_node_859),
        .a(6'd46),
        .b(_T_957)
    );
    wire _node_860;
    MUX_UNSIGNED #(.width(1)) u_mux_931 (
        .y(_node_860),
        .sel(_node_859),
        .a(_T_871_46),
        .b(_node_858)
    );
    wire _node_861;
    EQ_UNSIGNED #(.width(6)) u_eq_932 (
        .y(_node_861),
        .a(6'd47),
        .b(_T_957)
    );
    wire _node_862;
    MUX_UNSIGNED #(.width(1)) u_mux_933 (
        .y(_node_862),
        .sel(_node_861),
        .a(_T_871_47),
        .b(_node_860)
    );
    wire _node_863;
    EQ_UNSIGNED #(.width(6)) u_eq_934 (
        .y(_node_863),
        .a(6'd48),
        .b(_T_957)
    );
    wire _node_864;
    MUX_UNSIGNED #(.width(1)) u_mux_935 (
        .y(_node_864),
        .sel(_node_863),
        .a(_T_871_48),
        .b(_node_862)
    );
    wire _node_865;
    EQ_UNSIGNED #(.width(6)) u_eq_936 (
        .y(_node_865),
        .a(6'd49),
        .b(_T_957)
    );
    wire _node_866;
    MUX_UNSIGNED #(.width(1)) u_mux_937 (
        .y(_node_866),
        .sel(_node_865),
        .a(_T_871_49),
        .b(_node_864)
    );
    wire _node_867;
    EQ_UNSIGNED #(.width(6)) u_eq_938 (
        .y(_node_867),
        .a(6'd50),
        .b(_T_957)
    );
    wire _node_868;
    MUX_UNSIGNED #(.width(1)) u_mux_939 (
        .y(_node_868),
        .sel(_node_867),
        .a(_T_871_50),
        .b(_node_866)
    );
    wire _node_869;
    EQ_UNSIGNED #(.width(6)) u_eq_940 (
        .y(_node_869),
        .a(6'd51),
        .b(_T_957)
    );
    wire _node_870;
    MUX_UNSIGNED #(.width(1)) u_mux_941 (
        .y(_node_870),
        .sel(_node_869),
        .a(_T_871_51),
        .b(_node_868)
    );
    wire _node_871;
    EQ_UNSIGNED #(.width(6)) u_eq_942 (
        .y(_node_871),
        .a(6'd52),
        .b(_T_957)
    );
    wire _node_872;
    MUX_UNSIGNED #(.width(1)) u_mux_943 (
        .y(_node_872),
        .sel(_node_871),
        .a(_T_871_52),
        .b(_node_870)
    );
    wire _T_958;
    BITWISEAND #(.width(1)) bitwiseand_944 (
        .y(_T_958),
        .a(_c__io_outs_2_ready),
        .b(_c__io_outs_2_valid)
    );
    wire [3:0] _T_960;
    BITS #(.width(6), .high(3), .low(0)) bits_945 (
        .y(_T_960),
        .in(_value_4__q)
    );
    wire _T_962;
    EQ_UNSIGNED #(.width(1)) u_eq_946 (
        .y(_T_962),
        .a(reset),
        .b(1'h0)
    );
    wire [3:0] _T_964;
    BITS #(.width(6), .high(3), .low(0)) bits_947 (
        .y(_T_964),
        .in(_value_4__q)
    );
    wire _node_873;
    EQ_UNSIGNED #(.width(4)) u_eq_948 (
        .y(_node_873),
        .a(4'd0),
        .b(_T_964)
    );
    wire [30:0] _node_874;
    assign _node_874 = _T_942_0;
    wire _node_875;
    EQ_UNSIGNED #(.width(4)) u_eq_949 (
        .y(_node_875),
        .a(4'd1),
        .b(_T_964)
    );
    wire [30:0] _node_876;
    MUX_UNSIGNED #(.width(31)) u_mux_950 (
        .y(_node_876),
        .sel(_node_875),
        .a(_T_942_1),
        .b(_node_874)
    );
    wire _node_877;
    EQ_UNSIGNED #(.width(4)) u_eq_951 (
        .y(_node_877),
        .a(4'd2),
        .b(_T_964)
    );
    wire [30:0] _node_878;
    MUX_UNSIGNED #(.width(31)) u_mux_952 (
        .y(_node_878),
        .sel(_node_877),
        .a(_T_942_2),
        .b(_node_876)
    );
    wire _node_879;
    EQ_UNSIGNED #(.width(4)) u_eq_953 (
        .y(_node_879),
        .a(4'd3),
        .b(_T_964)
    );
    wire [30:0] _node_880;
    MUX_UNSIGNED #(.width(31)) u_mux_954 (
        .y(_node_880),
        .sel(_node_879),
        .a(_T_942_3),
        .b(_node_878)
    );
    wire _node_881;
    EQ_UNSIGNED #(.width(4)) u_eq_955 (
        .y(_node_881),
        .a(4'd4),
        .b(_T_964)
    );
    wire [30:0] _node_882;
    MUX_UNSIGNED #(.width(31)) u_mux_956 (
        .y(_node_882),
        .sel(_node_881),
        .a(_T_942_4),
        .b(_node_880)
    );
    wire _node_883;
    EQ_UNSIGNED #(.width(4)) u_eq_957 (
        .y(_node_883),
        .a(4'd5),
        .b(_T_964)
    );
    wire [30:0] _node_884;
    MUX_UNSIGNED #(.width(31)) u_mux_958 (
        .y(_node_884),
        .sel(_node_883),
        .a(_T_942_5),
        .b(_node_882)
    );
    wire _node_885;
    EQ_UNSIGNED #(.width(4)) u_eq_959 (
        .y(_node_885),
        .a(4'd6),
        .b(_T_964)
    );
    wire [30:0] _node_886;
    MUX_UNSIGNED #(.width(31)) u_mux_960 (
        .y(_node_886),
        .sel(_node_885),
        .a(_T_942_6),
        .b(_node_884)
    );
    wire _node_887;
    EQ_UNSIGNED #(.width(4)) u_eq_961 (
        .y(_node_887),
        .a(4'd7),
        .b(_T_964)
    );
    wire [30:0] _node_888;
    MUX_UNSIGNED #(.width(31)) u_mux_962 (
        .y(_node_888),
        .sel(_node_887),
        .a(_T_942_7),
        .b(_node_886)
    );
    wire _node_889;
    EQ_UNSIGNED #(.width(4)) u_eq_963 (
        .y(_node_889),
        .a(4'd8),
        .b(_T_964)
    );
    wire [30:0] _node_890;
    MUX_UNSIGNED #(.width(31)) u_mux_964 (
        .y(_node_890),
        .sel(_node_889),
        .a(_T_942_8),
        .b(_node_888)
    );
    wire _node_891;
    EQ_UNSIGNED #(.width(4)) u_eq_965 (
        .y(_node_891),
        .a(4'd9),
        .b(_T_964)
    );
    wire [30:0] _node_892;
    MUX_UNSIGNED #(.width(31)) u_mux_966 (
        .y(_node_892),
        .sel(_node_891),
        .a(_T_942_9),
        .b(_node_890)
    );
    wire _node_893;
    EQ_UNSIGNED #(.width(4)) u_eq_967 (
        .y(_node_893),
        .a(4'd10),
        .b(_T_964)
    );
    wire [30:0] _node_894;
    MUX_UNSIGNED #(.width(31)) u_mux_968 (
        .y(_node_894),
        .sel(_node_893),
        .a(_T_942_10),
        .b(_node_892)
    );
    wire _T_965;
    wire [63:0] _WTEMP_32;
    PAD_UNSIGNED #(.width(31), .n(64)) u_pad_969 (
        .y(_WTEMP_32),
        .in(_node_894)
    );
    NEQ_UNSIGNED #(.width(64)) u_neq_970 (
        .y(_T_965),
        .a(_c__io_outs_2_bits_body),
        .b(_WTEMP_32)
    );
    wire [3:0] _T_967;
    BITS #(.width(6), .high(3), .low(0)) bits_971 (
        .y(_T_967),
        .in(_value_4__q)
    );
    wire _T_969;
    EQ_UNSIGNED #(.width(1)) u_eq_972 (
        .y(_T_969),
        .a(reset),
        .b(1'h0)
    );
    wire _T_971;
    BITWISEOR #(.width(1)) bitwiseor_973 (
        .y(_T_971),
        .a(1'h0),
        .b(reset)
    );
    wire _T_973;
    EQ_UNSIGNED #(.width(1)) u_eq_974 (
        .y(_T_973),
        .a(_T_971),
        .b(1'h0)
    );
    wire _T_975;
    EQ_UNSIGNED #(.width(1)) u_eq_975 (
        .y(_T_975),
        .a(reset),
        .b(1'h0)
    );
    wire _T_977;
    EQ_UNSIGNED #(.width(6)) u_eq_976 (
        .y(_T_977),
        .a(_value_4__q),
        .b(6'h20)
    );
    wire [6:0] _T_979;
    wire [5:0] _WTEMP_33;
    PAD_UNSIGNED #(.width(1), .n(6)) u_pad_977 (
        .y(_WTEMP_33),
        .in(1'h1)
    );
    ADD_UNSIGNED #(.width(6)) u_add_978 (
        .y(_T_979),
        .a(_value_4__q),
        .b(_WTEMP_33)
    );
    wire [5:0] _T_980;
    TAIL #(.width(7), .n(1)) tail_979 (
        .y(_T_980),
        .in(_T_979)
    );
    wire _T_983;
    EQ_UNSIGNED #(.width(1)) u_eq_980 (
        .y(_T_983),
        .a(__T_13__q),
        .b(1'h0)
    );
    wire _T_985;
    wire [7:0] _WTEMP_34;
    PAD_UNSIGNED #(.width(6), .n(8)) u_pad_981 (
        .y(_WTEMP_34),
        .in(6'h20)
    );
    EQ_UNSIGNED #(.width(8)) u_eq_982 (
        .y(_T_985),
        .a(__T_10__q),
        .b(_WTEMP_34)
    );
    wire _node_895;
    MUX_UNSIGNED #(.width(1)) u_mux_983 (
        .y(_node_895),
        .sel(_T_784),
        .a(_node_765),
        .b(__T_13__q)
    );
    wire [8:0] _T_988;
    wire [7:0] _WTEMP_35;
    PAD_UNSIGNED #(.width(1), .n(8)) u_pad_984 (
        .y(_WTEMP_35),
        .in(1'h1)
    );
    ADD_UNSIGNED #(.width(8)) u_add_985 (
        .y(_T_988),
        .a(__T_10__q),
        .b(_WTEMP_35)
    );
    wire [7:0] _T_989;
    TAIL #(.width(9), .n(1)) tail_986 (
        .y(_T_989),
        .in(_T_988)
    );
    wire [7:0] _node_896;
    MUX_UNSIGNED #(.width(8)) u_mux_987 (
        .y(_node_896),
        .sel(_T_784),
        .a(_node_764),
        .b(__T_10__q)
    );
    wire _node_897;
    MUX_UNSIGNED #(.width(1)) u_mux_988 (
        .y(_node_897),
        .sel(_T_985),
        .a(1'h1),
        .b(_node_895)
    );
    wire _node_898;
    MUX_UNSIGNED #(.width(1)) u_mux_989 (
        .y(_node_898),
        .sel(_T_784),
        .a(_node_765),
        .b(__T_13__q)
    );
    wire [7:0] _node_899;
    MUX_UNSIGNED #(.width(8)) u_mux_990 (
        .y(_node_899),
        .sel(_T_983),
        .a(_T_989),
        .b(_node_896)
    );
    wire [7:0] _node_900;
    MUX_UNSIGNED #(.width(8)) u_mux_991 (
        .y(_node_900),
        .sel(_T_784),
        .a(_node_764),
        .b(__T_10__q)
    );
    wire _node_901;
    MUX_UNSIGNED #(.width(1)) u_mux_992 (
        .y(_node_901),
        .sel(_T_983),
        .a(_node_897),
        .b(_node_898)
    );
    wire _node_902;
    MUX_UNSIGNED #(.width(1)) u_mux_993 (
        .y(_node_902),
        .sel(_T_784),
        .a(_node_765),
        .b(__T_13__q)
    );
    wire [5:0] _node_903;
    wire [5:0] _WTEMP_36;
    PAD_UNSIGNED #(.width(1), .n(6)) u_pad_994 (
        .y(_WTEMP_36),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(6)) u_mux_995 (
        .y(_node_903),
        .sel(_T_977),
        .a(_WTEMP_36),
        .b(_T_980)
    );
    wire _T_1045_0;
    wire _T_1045_1;
    wire _T_1045_2;
    wire _T_1045_3;
    wire _T_1045_4;
    wire _T_1045_5;
    wire _T_1045_6;
    wire _T_1045_7;
    wire _T_1045_8;
    wire _T_1045_9;
    wire _T_1045_10;
    wire _T_1045_11;
    wire _T_1045_12;
    wire _T_1045_13;
    wire _T_1045_14;
    wire _T_1045_15;
    wire _T_1045_16;
    wire _T_1045_17;
    wire _T_1045_18;
    wire _T_1045_19;
    wire _T_1045_20;
    wire _T_1045_21;
    wire _T_1045_22;
    wire _T_1045_23;
    wire _T_1045_24;
    wire _T_1045_25;
    wire _T_1045_26;
    wire _T_1045_27;
    wire _T_1045_28;
    wire _T_1045_29;
    wire _T_1045_30;
    wire _T_1045_31;
    wire _T_1045_32;
    wire _T_1045_33;
    wire _T_1045_34;
    wire _T_1045_35;
    wire _T_1045_36;
    wire _T_1045_37;
    wire _T_1045_38;
    wire _T_1045_39;
    wire _T_1045_40;
    wire _T_1045_41;
    wire _T_1045_42;
    wire _T_1045_43;
    wire _T_1045_44;
    wire _T_1045_45;
    wire _T_1045_46;
    wire _T_1045_47;
    wire _T_1045_48;
    wire _T_1045_49;
    wire _T_1045_50;
    wire _T_1045_51;
    wire _T_1045_52;
    wire [5:0] _value_5__q;
    wire [5:0] _value_5__d;
    DFF_POSCLK #(.width(6)) value_5 (
        .q(_value_5__q),
        .d(_value_5__d),
        .clk(clock)
    );
    wire [5:0] _WTEMP_37;
    MUX_UNSIGNED #(.width(6)) u_mux_996 (
        .y(_value_5__d),
        .sel(reset),
        .a(6'h0),
        .b(_WTEMP_37)
    );
    wire [30:0] _T_1111_0;
    wire [30:0] _T_1111_1;
    wire [30:0] _T_1111_2;
    wire [30:0] _T_1111_3;
    wire [30:0] _T_1111_4;
    wire [30:0] _T_1111_5;
    wire [5:0] _T_1121;
    BITS #(.width(8), .high(5), .low(0)) bits_997 (
        .y(_T_1121),
        .in(__T_10__q)
    );
    wire _node_904;
    EQ_UNSIGNED #(.width(6)) u_eq_998 (
        .y(_node_904),
        .a(6'd0),
        .b(_T_1121)
    );
    wire _node_905;
    assign _node_905 = _T_1045_0;
    wire _node_906;
    EQ_UNSIGNED #(.width(6)) u_eq_999 (
        .y(_node_906),
        .a(6'd1),
        .b(_T_1121)
    );
    wire _node_907;
    MUX_UNSIGNED #(.width(1)) u_mux_1000 (
        .y(_node_907),
        .sel(_node_906),
        .a(_T_1045_1),
        .b(_node_905)
    );
    wire _node_908;
    EQ_UNSIGNED #(.width(6)) u_eq_1001 (
        .y(_node_908),
        .a(6'd2),
        .b(_T_1121)
    );
    wire _node_909;
    MUX_UNSIGNED #(.width(1)) u_mux_1002 (
        .y(_node_909),
        .sel(_node_908),
        .a(_T_1045_2),
        .b(_node_907)
    );
    wire _node_910;
    EQ_UNSIGNED #(.width(6)) u_eq_1003 (
        .y(_node_910),
        .a(6'd3),
        .b(_T_1121)
    );
    wire _node_911;
    MUX_UNSIGNED #(.width(1)) u_mux_1004 (
        .y(_node_911),
        .sel(_node_910),
        .a(_T_1045_3),
        .b(_node_909)
    );
    wire _node_912;
    EQ_UNSIGNED #(.width(6)) u_eq_1005 (
        .y(_node_912),
        .a(6'd4),
        .b(_T_1121)
    );
    wire _node_913;
    MUX_UNSIGNED #(.width(1)) u_mux_1006 (
        .y(_node_913),
        .sel(_node_912),
        .a(_T_1045_4),
        .b(_node_911)
    );
    wire _node_914;
    EQ_UNSIGNED #(.width(6)) u_eq_1007 (
        .y(_node_914),
        .a(6'd5),
        .b(_T_1121)
    );
    wire _node_915;
    MUX_UNSIGNED #(.width(1)) u_mux_1008 (
        .y(_node_915),
        .sel(_node_914),
        .a(_T_1045_5),
        .b(_node_913)
    );
    wire _node_916;
    EQ_UNSIGNED #(.width(6)) u_eq_1009 (
        .y(_node_916),
        .a(6'd6),
        .b(_T_1121)
    );
    wire _node_917;
    MUX_UNSIGNED #(.width(1)) u_mux_1010 (
        .y(_node_917),
        .sel(_node_916),
        .a(_T_1045_6),
        .b(_node_915)
    );
    wire _node_918;
    EQ_UNSIGNED #(.width(6)) u_eq_1011 (
        .y(_node_918),
        .a(6'd7),
        .b(_T_1121)
    );
    wire _node_919;
    MUX_UNSIGNED #(.width(1)) u_mux_1012 (
        .y(_node_919),
        .sel(_node_918),
        .a(_T_1045_7),
        .b(_node_917)
    );
    wire _node_920;
    EQ_UNSIGNED #(.width(6)) u_eq_1013 (
        .y(_node_920),
        .a(6'd8),
        .b(_T_1121)
    );
    wire _node_921;
    MUX_UNSIGNED #(.width(1)) u_mux_1014 (
        .y(_node_921),
        .sel(_node_920),
        .a(_T_1045_8),
        .b(_node_919)
    );
    wire _node_922;
    EQ_UNSIGNED #(.width(6)) u_eq_1015 (
        .y(_node_922),
        .a(6'd9),
        .b(_T_1121)
    );
    wire _node_923;
    MUX_UNSIGNED #(.width(1)) u_mux_1016 (
        .y(_node_923),
        .sel(_node_922),
        .a(_T_1045_9),
        .b(_node_921)
    );
    wire _node_924;
    EQ_UNSIGNED #(.width(6)) u_eq_1017 (
        .y(_node_924),
        .a(6'd10),
        .b(_T_1121)
    );
    wire _node_925;
    MUX_UNSIGNED #(.width(1)) u_mux_1018 (
        .y(_node_925),
        .sel(_node_924),
        .a(_T_1045_10),
        .b(_node_923)
    );
    wire _node_926;
    EQ_UNSIGNED #(.width(6)) u_eq_1019 (
        .y(_node_926),
        .a(6'd11),
        .b(_T_1121)
    );
    wire _node_927;
    MUX_UNSIGNED #(.width(1)) u_mux_1020 (
        .y(_node_927),
        .sel(_node_926),
        .a(_T_1045_11),
        .b(_node_925)
    );
    wire _node_928;
    EQ_UNSIGNED #(.width(6)) u_eq_1021 (
        .y(_node_928),
        .a(6'd12),
        .b(_T_1121)
    );
    wire _node_929;
    MUX_UNSIGNED #(.width(1)) u_mux_1022 (
        .y(_node_929),
        .sel(_node_928),
        .a(_T_1045_12),
        .b(_node_927)
    );
    wire _node_930;
    EQ_UNSIGNED #(.width(6)) u_eq_1023 (
        .y(_node_930),
        .a(6'd13),
        .b(_T_1121)
    );
    wire _node_931;
    MUX_UNSIGNED #(.width(1)) u_mux_1024 (
        .y(_node_931),
        .sel(_node_930),
        .a(_T_1045_13),
        .b(_node_929)
    );
    wire _node_932;
    EQ_UNSIGNED #(.width(6)) u_eq_1025 (
        .y(_node_932),
        .a(6'd14),
        .b(_T_1121)
    );
    wire _node_933;
    MUX_UNSIGNED #(.width(1)) u_mux_1026 (
        .y(_node_933),
        .sel(_node_932),
        .a(_T_1045_14),
        .b(_node_931)
    );
    wire _node_934;
    EQ_UNSIGNED #(.width(6)) u_eq_1027 (
        .y(_node_934),
        .a(6'd15),
        .b(_T_1121)
    );
    wire _node_935;
    MUX_UNSIGNED #(.width(1)) u_mux_1028 (
        .y(_node_935),
        .sel(_node_934),
        .a(_T_1045_15),
        .b(_node_933)
    );
    wire _node_936;
    EQ_UNSIGNED #(.width(6)) u_eq_1029 (
        .y(_node_936),
        .a(6'd16),
        .b(_T_1121)
    );
    wire _node_937;
    MUX_UNSIGNED #(.width(1)) u_mux_1030 (
        .y(_node_937),
        .sel(_node_936),
        .a(_T_1045_16),
        .b(_node_935)
    );
    wire _node_938;
    EQ_UNSIGNED #(.width(6)) u_eq_1031 (
        .y(_node_938),
        .a(6'd17),
        .b(_T_1121)
    );
    wire _node_939;
    MUX_UNSIGNED #(.width(1)) u_mux_1032 (
        .y(_node_939),
        .sel(_node_938),
        .a(_T_1045_17),
        .b(_node_937)
    );
    wire _node_940;
    EQ_UNSIGNED #(.width(6)) u_eq_1033 (
        .y(_node_940),
        .a(6'd18),
        .b(_T_1121)
    );
    wire _node_941;
    MUX_UNSIGNED #(.width(1)) u_mux_1034 (
        .y(_node_941),
        .sel(_node_940),
        .a(_T_1045_18),
        .b(_node_939)
    );
    wire _node_942;
    EQ_UNSIGNED #(.width(6)) u_eq_1035 (
        .y(_node_942),
        .a(6'd19),
        .b(_T_1121)
    );
    wire _node_943;
    MUX_UNSIGNED #(.width(1)) u_mux_1036 (
        .y(_node_943),
        .sel(_node_942),
        .a(_T_1045_19),
        .b(_node_941)
    );
    wire _node_944;
    EQ_UNSIGNED #(.width(6)) u_eq_1037 (
        .y(_node_944),
        .a(6'd20),
        .b(_T_1121)
    );
    wire _node_945;
    MUX_UNSIGNED #(.width(1)) u_mux_1038 (
        .y(_node_945),
        .sel(_node_944),
        .a(_T_1045_20),
        .b(_node_943)
    );
    wire _node_946;
    EQ_UNSIGNED #(.width(6)) u_eq_1039 (
        .y(_node_946),
        .a(6'd21),
        .b(_T_1121)
    );
    wire _node_947;
    MUX_UNSIGNED #(.width(1)) u_mux_1040 (
        .y(_node_947),
        .sel(_node_946),
        .a(_T_1045_21),
        .b(_node_945)
    );
    wire _node_948;
    EQ_UNSIGNED #(.width(6)) u_eq_1041 (
        .y(_node_948),
        .a(6'd22),
        .b(_T_1121)
    );
    wire _node_949;
    MUX_UNSIGNED #(.width(1)) u_mux_1042 (
        .y(_node_949),
        .sel(_node_948),
        .a(_T_1045_22),
        .b(_node_947)
    );
    wire _node_950;
    EQ_UNSIGNED #(.width(6)) u_eq_1043 (
        .y(_node_950),
        .a(6'd23),
        .b(_T_1121)
    );
    wire _node_951;
    MUX_UNSIGNED #(.width(1)) u_mux_1044 (
        .y(_node_951),
        .sel(_node_950),
        .a(_T_1045_23),
        .b(_node_949)
    );
    wire _node_952;
    EQ_UNSIGNED #(.width(6)) u_eq_1045 (
        .y(_node_952),
        .a(6'd24),
        .b(_T_1121)
    );
    wire _node_953;
    MUX_UNSIGNED #(.width(1)) u_mux_1046 (
        .y(_node_953),
        .sel(_node_952),
        .a(_T_1045_24),
        .b(_node_951)
    );
    wire _node_954;
    EQ_UNSIGNED #(.width(6)) u_eq_1047 (
        .y(_node_954),
        .a(6'd25),
        .b(_T_1121)
    );
    wire _node_955;
    MUX_UNSIGNED #(.width(1)) u_mux_1048 (
        .y(_node_955),
        .sel(_node_954),
        .a(_T_1045_25),
        .b(_node_953)
    );
    wire _node_956;
    EQ_UNSIGNED #(.width(6)) u_eq_1049 (
        .y(_node_956),
        .a(6'd26),
        .b(_T_1121)
    );
    wire _node_957;
    MUX_UNSIGNED #(.width(1)) u_mux_1050 (
        .y(_node_957),
        .sel(_node_956),
        .a(_T_1045_26),
        .b(_node_955)
    );
    wire _node_958;
    EQ_UNSIGNED #(.width(6)) u_eq_1051 (
        .y(_node_958),
        .a(6'd27),
        .b(_T_1121)
    );
    wire _node_959;
    MUX_UNSIGNED #(.width(1)) u_mux_1052 (
        .y(_node_959),
        .sel(_node_958),
        .a(_T_1045_27),
        .b(_node_957)
    );
    wire _node_960;
    EQ_UNSIGNED #(.width(6)) u_eq_1053 (
        .y(_node_960),
        .a(6'd28),
        .b(_T_1121)
    );
    wire _node_961;
    MUX_UNSIGNED #(.width(1)) u_mux_1054 (
        .y(_node_961),
        .sel(_node_960),
        .a(_T_1045_28),
        .b(_node_959)
    );
    wire _node_962;
    EQ_UNSIGNED #(.width(6)) u_eq_1055 (
        .y(_node_962),
        .a(6'd29),
        .b(_T_1121)
    );
    wire _node_963;
    MUX_UNSIGNED #(.width(1)) u_mux_1056 (
        .y(_node_963),
        .sel(_node_962),
        .a(_T_1045_29),
        .b(_node_961)
    );
    wire _node_964;
    EQ_UNSIGNED #(.width(6)) u_eq_1057 (
        .y(_node_964),
        .a(6'd30),
        .b(_T_1121)
    );
    wire _node_965;
    MUX_UNSIGNED #(.width(1)) u_mux_1058 (
        .y(_node_965),
        .sel(_node_964),
        .a(_T_1045_30),
        .b(_node_963)
    );
    wire _node_966;
    EQ_UNSIGNED #(.width(6)) u_eq_1059 (
        .y(_node_966),
        .a(6'd31),
        .b(_T_1121)
    );
    wire _node_967;
    MUX_UNSIGNED #(.width(1)) u_mux_1060 (
        .y(_node_967),
        .sel(_node_966),
        .a(_T_1045_31),
        .b(_node_965)
    );
    wire _node_968;
    EQ_UNSIGNED #(.width(6)) u_eq_1061 (
        .y(_node_968),
        .a(6'd32),
        .b(_T_1121)
    );
    wire _node_969;
    MUX_UNSIGNED #(.width(1)) u_mux_1062 (
        .y(_node_969),
        .sel(_node_968),
        .a(_T_1045_32),
        .b(_node_967)
    );
    wire _node_970;
    EQ_UNSIGNED #(.width(6)) u_eq_1063 (
        .y(_node_970),
        .a(6'd33),
        .b(_T_1121)
    );
    wire _node_971;
    MUX_UNSIGNED #(.width(1)) u_mux_1064 (
        .y(_node_971),
        .sel(_node_970),
        .a(_T_1045_33),
        .b(_node_969)
    );
    wire _node_972;
    EQ_UNSIGNED #(.width(6)) u_eq_1065 (
        .y(_node_972),
        .a(6'd34),
        .b(_T_1121)
    );
    wire _node_973;
    MUX_UNSIGNED #(.width(1)) u_mux_1066 (
        .y(_node_973),
        .sel(_node_972),
        .a(_T_1045_34),
        .b(_node_971)
    );
    wire _node_974;
    EQ_UNSIGNED #(.width(6)) u_eq_1067 (
        .y(_node_974),
        .a(6'd35),
        .b(_T_1121)
    );
    wire _node_975;
    MUX_UNSIGNED #(.width(1)) u_mux_1068 (
        .y(_node_975),
        .sel(_node_974),
        .a(_T_1045_35),
        .b(_node_973)
    );
    wire _node_976;
    EQ_UNSIGNED #(.width(6)) u_eq_1069 (
        .y(_node_976),
        .a(6'd36),
        .b(_T_1121)
    );
    wire _node_977;
    MUX_UNSIGNED #(.width(1)) u_mux_1070 (
        .y(_node_977),
        .sel(_node_976),
        .a(_T_1045_36),
        .b(_node_975)
    );
    wire _node_978;
    EQ_UNSIGNED #(.width(6)) u_eq_1071 (
        .y(_node_978),
        .a(6'd37),
        .b(_T_1121)
    );
    wire _node_979;
    MUX_UNSIGNED #(.width(1)) u_mux_1072 (
        .y(_node_979),
        .sel(_node_978),
        .a(_T_1045_37),
        .b(_node_977)
    );
    wire _node_980;
    EQ_UNSIGNED #(.width(6)) u_eq_1073 (
        .y(_node_980),
        .a(6'd38),
        .b(_T_1121)
    );
    wire _node_981;
    MUX_UNSIGNED #(.width(1)) u_mux_1074 (
        .y(_node_981),
        .sel(_node_980),
        .a(_T_1045_38),
        .b(_node_979)
    );
    wire _node_982;
    EQ_UNSIGNED #(.width(6)) u_eq_1075 (
        .y(_node_982),
        .a(6'd39),
        .b(_T_1121)
    );
    wire _node_983;
    MUX_UNSIGNED #(.width(1)) u_mux_1076 (
        .y(_node_983),
        .sel(_node_982),
        .a(_T_1045_39),
        .b(_node_981)
    );
    wire _node_984;
    EQ_UNSIGNED #(.width(6)) u_eq_1077 (
        .y(_node_984),
        .a(6'd40),
        .b(_T_1121)
    );
    wire _node_985;
    MUX_UNSIGNED #(.width(1)) u_mux_1078 (
        .y(_node_985),
        .sel(_node_984),
        .a(_T_1045_40),
        .b(_node_983)
    );
    wire _node_986;
    EQ_UNSIGNED #(.width(6)) u_eq_1079 (
        .y(_node_986),
        .a(6'd41),
        .b(_T_1121)
    );
    wire _node_987;
    MUX_UNSIGNED #(.width(1)) u_mux_1080 (
        .y(_node_987),
        .sel(_node_986),
        .a(_T_1045_41),
        .b(_node_985)
    );
    wire _node_988;
    EQ_UNSIGNED #(.width(6)) u_eq_1081 (
        .y(_node_988),
        .a(6'd42),
        .b(_T_1121)
    );
    wire _node_989;
    MUX_UNSIGNED #(.width(1)) u_mux_1082 (
        .y(_node_989),
        .sel(_node_988),
        .a(_T_1045_42),
        .b(_node_987)
    );
    wire _node_990;
    EQ_UNSIGNED #(.width(6)) u_eq_1083 (
        .y(_node_990),
        .a(6'd43),
        .b(_T_1121)
    );
    wire _node_991;
    MUX_UNSIGNED #(.width(1)) u_mux_1084 (
        .y(_node_991),
        .sel(_node_990),
        .a(_T_1045_43),
        .b(_node_989)
    );
    wire _node_992;
    EQ_UNSIGNED #(.width(6)) u_eq_1085 (
        .y(_node_992),
        .a(6'd44),
        .b(_T_1121)
    );
    wire _node_993;
    MUX_UNSIGNED #(.width(1)) u_mux_1086 (
        .y(_node_993),
        .sel(_node_992),
        .a(_T_1045_44),
        .b(_node_991)
    );
    wire _node_994;
    EQ_UNSIGNED #(.width(6)) u_eq_1087 (
        .y(_node_994),
        .a(6'd45),
        .b(_T_1121)
    );
    wire _node_995;
    MUX_UNSIGNED #(.width(1)) u_mux_1088 (
        .y(_node_995),
        .sel(_node_994),
        .a(_T_1045_45),
        .b(_node_993)
    );
    wire _node_996;
    EQ_UNSIGNED #(.width(6)) u_eq_1089 (
        .y(_node_996),
        .a(6'd46),
        .b(_T_1121)
    );
    wire _node_997;
    MUX_UNSIGNED #(.width(1)) u_mux_1090 (
        .y(_node_997),
        .sel(_node_996),
        .a(_T_1045_46),
        .b(_node_995)
    );
    wire _node_998;
    EQ_UNSIGNED #(.width(6)) u_eq_1091 (
        .y(_node_998),
        .a(6'd47),
        .b(_T_1121)
    );
    wire _node_999;
    MUX_UNSIGNED #(.width(1)) u_mux_1092 (
        .y(_node_999),
        .sel(_node_998),
        .a(_T_1045_47),
        .b(_node_997)
    );
    wire _node_1000;
    EQ_UNSIGNED #(.width(6)) u_eq_1093 (
        .y(_node_1000),
        .a(6'd48),
        .b(_T_1121)
    );
    wire _node_1001;
    MUX_UNSIGNED #(.width(1)) u_mux_1094 (
        .y(_node_1001),
        .sel(_node_1000),
        .a(_T_1045_48),
        .b(_node_999)
    );
    wire _node_1002;
    EQ_UNSIGNED #(.width(6)) u_eq_1095 (
        .y(_node_1002),
        .a(6'd49),
        .b(_T_1121)
    );
    wire _node_1003;
    MUX_UNSIGNED #(.width(1)) u_mux_1096 (
        .y(_node_1003),
        .sel(_node_1002),
        .a(_T_1045_49),
        .b(_node_1001)
    );
    wire _node_1004;
    EQ_UNSIGNED #(.width(6)) u_eq_1097 (
        .y(_node_1004),
        .a(6'd50),
        .b(_T_1121)
    );
    wire _node_1005;
    MUX_UNSIGNED #(.width(1)) u_mux_1098 (
        .y(_node_1005),
        .sel(_node_1004),
        .a(_T_1045_50),
        .b(_node_1003)
    );
    wire _node_1006;
    EQ_UNSIGNED #(.width(6)) u_eq_1099 (
        .y(_node_1006),
        .a(6'd51),
        .b(_T_1121)
    );
    wire _node_1007;
    MUX_UNSIGNED #(.width(1)) u_mux_1100 (
        .y(_node_1007),
        .sel(_node_1006),
        .a(_T_1045_51),
        .b(_node_1005)
    );
    wire _node_1008;
    EQ_UNSIGNED #(.width(6)) u_eq_1101 (
        .y(_node_1008),
        .a(6'd52),
        .b(_T_1121)
    );
    wire _node_1009;
    MUX_UNSIGNED #(.width(1)) u_mux_1102 (
        .y(_node_1009),
        .sel(_node_1008),
        .a(_T_1045_52),
        .b(_node_1007)
    );
    wire _T_1122;
    BITWISEAND #(.width(1)) bitwiseand_1103 (
        .y(_T_1122),
        .a(_c__io_outs_3_ready),
        .b(_c__io_outs_3_valid)
    );
    wire [2:0] _T_1124;
    BITS #(.width(6), .high(2), .low(0)) bits_1104 (
        .y(_T_1124),
        .in(_value_5__q)
    );
    wire _T_1126;
    EQ_UNSIGNED #(.width(1)) u_eq_1105 (
        .y(_T_1126),
        .a(reset),
        .b(1'h0)
    );
    wire [2:0] _T_1128;
    BITS #(.width(6), .high(2), .low(0)) bits_1106 (
        .y(_T_1128),
        .in(_value_5__q)
    );
    wire _node_1010;
    EQ_UNSIGNED #(.width(3)) u_eq_1107 (
        .y(_node_1010),
        .a(3'd0),
        .b(_T_1128)
    );
    wire [30:0] _node_1011;
    assign _node_1011 = _T_1111_0;
    wire _node_1012;
    EQ_UNSIGNED #(.width(3)) u_eq_1108 (
        .y(_node_1012),
        .a(3'd1),
        .b(_T_1128)
    );
    wire [30:0] _node_1013;
    MUX_UNSIGNED #(.width(31)) u_mux_1109 (
        .y(_node_1013),
        .sel(_node_1012),
        .a(_T_1111_1),
        .b(_node_1011)
    );
    wire _node_1014;
    EQ_UNSIGNED #(.width(3)) u_eq_1110 (
        .y(_node_1014),
        .a(3'd2),
        .b(_T_1128)
    );
    wire [30:0] _node_1015;
    MUX_UNSIGNED #(.width(31)) u_mux_1111 (
        .y(_node_1015),
        .sel(_node_1014),
        .a(_T_1111_2),
        .b(_node_1013)
    );
    wire _node_1016;
    EQ_UNSIGNED #(.width(3)) u_eq_1112 (
        .y(_node_1016),
        .a(3'd3),
        .b(_T_1128)
    );
    wire [30:0] _node_1017;
    MUX_UNSIGNED #(.width(31)) u_mux_1113 (
        .y(_node_1017),
        .sel(_node_1016),
        .a(_T_1111_3),
        .b(_node_1015)
    );
    wire _node_1018;
    EQ_UNSIGNED #(.width(3)) u_eq_1114 (
        .y(_node_1018),
        .a(3'd4),
        .b(_T_1128)
    );
    wire [30:0] _node_1019;
    MUX_UNSIGNED #(.width(31)) u_mux_1115 (
        .y(_node_1019),
        .sel(_node_1018),
        .a(_T_1111_4),
        .b(_node_1017)
    );
    wire _node_1020;
    EQ_UNSIGNED #(.width(3)) u_eq_1116 (
        .y(_node_1020),
        .a(3'd5),
        .b(_T_1128)
    );
    wire [30:0] _node_1021;
    MUX_UNSIGNED #(.width(31)) u_mux_1117 (
        .y(_node_1021),
        .sel(_node_1020),
        .a(_T_1111_5),
        .b(_node_1019)
    );
    wire _T_1129;
    wire [63:0] _WTEMP_38;
    PAD_UNSIGNED #(.width(31), .n(64)) u_pad_1118 (
        .y(_WTEMP_38),
        .in(_node_1021)
    );
    NEQ_UNSIGNED #(.width(64)) u_neq_1119 (
        .y(_T_1129),
        .a(_c__io_outs_3_bits_body),
        .b(_WTEMP_38)
    );
    wire [2:0] _T_1131;
    BITS #(.width(6), .high(2), .low(0)) bits_1120 (
        .y(_T_1131),
        .in(_value_5__q)
    );
    wire _T_1133;
    EQ_UNSIGNED #(.width(1)) u_eq_1121 (
        .y(_T_1133),
        .a(reset),
        .b(1'h0)
    );
    wire _T_1135;
    BITWISEOR #(.width(1)) bitwiseor_1122 (
        .y(_T_1135),
        .a(1'h0),
        .b(reset)
    );
    wire _T_1137;
    EQ_UNSIGNED #(.width(1)) u_eq_1123 (
        .y(_T_1137),
        .a(_T_1135),
        .b(1'h0)
    );
    wire _T_1139;
    EQ_UNSIGNED #(.width(1)) u_eq_1124 (
        .y(_T_1139),
        .a(reset),
        .b(1'h0)
    );
    wire _T_1141;
    EQ_UNSIGNED #(.width(6)) u_eq_1125 (
        .y(_T_1141),
        .a(_value_5__q),
        .b(6'h20)
    );
    wire [6:0] _T_1143;
    wire [5:0] _WTEMP_39;
    PAD_UNSIGNED #(.width(1), .n(6)) u_pad_1126 (
        .y(_WTEMP_39),
        .in(1'h1)
    );
    ADD_UNSIGNED #(.width(6)) u_add_1127 (
        .y(_T_1143),
        .a(_value_5__q),
        .b(_WTEMP_39)
    );
    wire [5:0] _T_1144;
    TAIL #(.width(7), .n(1)) tail_1128 (
        .y(_T_1144),
        .in(_T_1143)
    );
    wire _T_1147;
    EQ_UNSIGNED #(.width(1)) u_eq_1129 (
        .y(_T_1147),
        .a(__T_13__q),
        .b(1'h0)
    );
    wire _T_1149;
    wire [7:0] _WTEMP_40;
    PAD_UNSIGNED #(.width(6), .n(8)) u_pad_1130 (
        .y(_WTEMP_40),
        .in(6'h20)
    );
    EQ_UNSIGNED #(.width(8)) u_eq_1131 (
        .y(_T_1149),
        .a(__T_10__q),
        .b(_WTEMP_40)
    );
    wire _node_1022;
    MUX_UNSIGNED #(.width(1)) u_mux_1132 (
        .y(_node_1022),
        .sel(_T_958),
        .a(_node_901),
        .b(_node_902)
    );
    wire [8:0] _T_1152;
    wire [7:0] _WTEMP_41;
    PAD_UNSIGNED #(.width(1), .n(8)) u_pad_1133 (
        .y(_WTEMP_41),
        .in(1'h1)
    );
    ADD_UNSIGNED #(.width(8)) u_add_1134 (
        .y(_T_1152),
        .a(__T_10__q),
        .b(_WTEMP_41)
    );
    wire [7:0] _T_1153;
    TAIL #(.width(9), .n(1)) tail_1135 (
        .y(_T_1153),
        .in(_T_1152)
    );
    wire [7:0] _node_1023;
    MUX_UNSIGNED #(.width(8)) u_mux_1136 (
        .y(_node_1023),
        .sel(_T_958),
        .a(_node_899),
        .b(_node_900)
    );
    wire _node_1024;
    MUX_UNSIGNED #(.width(1)) u_mux_1137 (
        .y(_node_1024),
        .sel(_T_1149),
        .a(1'h1),
        .b(_node_1022)
    );
    wire _node_1025;
    MUX_UNSIGNED #(.width(1)) u_mux_1138 (
        .y(_node_1025),
        .sel(_T_958),
        .a(_node_901),
        .b(_node_902)
    );
    wire [7:0] _node_1026;
    MUX_UNSIGNED #(.width(8)) u_mux_1139 (
        .y(_node_1026),
        .sel(_T_1147),
        .a(_T_1153),
        .b(_node_1023)
    );
    wire [7:0] _node_1027;
    MUX_UNSIGNED #(.width(8)) u_mux_1140 (
        .y(_node_1027),
        .sel(_T_958),
        .a(_node_899),
        .b(_node_900)
    );
    wire _node_1028;
    MUX_UNSIGNED #(.width(1)) u_mux_1141 (
        .y(_node_1028),
        .sel(_T_1147),
        .a(_node_1024),
        .b(_node_1025)
    );
    wire _node_1029;
    MUX_UNSIGNED #(.width(1)) u_mux_1142 (
        .y(_node_1029),
        .sel(_T_958),
        .a(_node_901),
        .b(_node_902)
    );
    wire [5:0] _node_1030;
    wire [5:0] _WTEMP_42;
    PAD_UNSIGNED #(.width(1), .n(6)) u_pad_1143 (
        .y(_WTEMP_42),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(6)) u_mux_1144 (
        .y(_node_1030),
        .sel(_T_1141),
        .a(_WTEMP_42),
        .b(_T_1144)
    );
    wire _T_1209_0;
    wire _T_1209_1;
    wire _T_1209_2;
    wire _T_1209_3;
    wire _T_1209_4;
    wire _T_1209_5;
    wire _T_1209_6;
    wire _T_1209_7;
    wire _T_1209_8;
    wire _T_1209_9;
    wire _T_1209_10;
    wire _T_1209_11;
    wire _T_1209_12;
    wire _T_1209_13;
    wire _T_1209_14;
    wire _T_1209_15;
    wire _T_1209_16;
    wire _T_1209_17;
    wire _T_1209_18;
    wire _T_1209_19;
    wire _T_1209_20;
    wire _T_1209_21;
    wire _T_1209_22;
    wire _T_1209_23;
    wire _T_1209_24;
    wire _T_1209_25;
    wire _T_1209_26;
    wire _T_1209_27;
    wire _T_1209_28;
    wire _T_1209_29;
    wire _T_1209_30;
    wire _T_1209_31;
    wire _T_1209_32;
    wire _T_1209_33;
    wire _T_1209_34;
    wire _T_1209_35;
    wire _T_1209_36;
    wire _T_1209_37;
    wire _T_1209_38;
    wire _T_1209_39;
    wire _T_1209_40;
    wire _T_1209_41;
    wire _T_1209_42;
    wire _T_1209_43;
    wire _T_1209_44;
    wire _T_1209_45;
    wire _T_1209_46;
    wire _T_1209_47;
    wire _T_1209_48;
    wire _T_1209_49;
    wire _T_1209_50;
    wire _T_1209_51;
    wire _T_1209_52;
    wire [5:0] _value_6__q;
    wire [5:0] _value_6__d;
    DFF_POSCLK #(.width(6)) value_6 (
        .q(_value_6__q),
        .d(_value_6__d),
        .clk(clock)
    );
    wire [5:0] _WTEMP_43;
    MUX_UNSIGNED #(.width(6)) u_mux_1145 (
        .y(_value_6__d),
        .sel(reset),
        .a(6'h0),
        .b(_WTEMP_43)
    );
    wire [28:0] _T_1274_0;
    wire [28:0] _T_1274_1;
    wire [28:0] _T_1274_2;
    wire [28:0] _T_1274_3;
    wire [28:0] _T_1274_4;
    wire [5:0] _T_1283;
    BITS #(.width(8), .high(5), .low(0)) bits_1146 (
        .y(_T_1283),
        .in(__T_10__q)
    );
    wire _node_1031;
    EQ_UNSIGNED #(.width(6)) u_eq_1147 (
        .y(_node_1031),
        .a(6'd0),
        .b(_T_1283)
    );
    wire _node_1032;
    assign _node_1032 = _T_1209_0;
    wire _node_1033;
    EQ_UNSIGNED #(.width(6)) u_eq_1148 (
        .y(_node_1033),
        .a(6'd1),
        .b(_T_1283)
    );
    wire _node_1034;
    MUX_UNSIGNED #(.width(1)) u_mux_1149 (
        .y(_node_1034),
        .sel(_node_1033),
        .a(_T_1209_1),
        .b(_node_1032)
    );
    wire _node_1035;
    EQ_UNSIGNED #(.width(6)) u_eq_1150 (
        .y(_node_1035),
        .a(6'd2),
        .b(_T_1283)
    );
    wire _node_1036;
    MUX_UNSIGNED #(.width(1)) u_mux_1151 (
        .y(_node_1036),
        .sel(_node_1035),
        .a(_T_1209_2),
        .b(_node_1034)
    );
    wire _node_1037;
    EQ_UNSIGNED #(.width(6)) u_eq_1152 (
        .y(_node_1037),
        .a(6'd3),
        .b(_T_1283)
    );
    wire _node_1038;
    MUX_UNSIGNED #(.width(1)) u_mux_1153 (
        .y(_node_1038),
        .sel(_node_1037),
        .a(_T_1209_3),
        .b(_node_1036)
    );
    wire _node_1039;
    EQ_UNSIGNED #(.width(6)) u_eq_1154 (
        .y(_node_1039),
        .a(6'd4),
        .b(_T_1283)
    );
    wire _node_1040;
    MUX_UNSIGNED #(.width(1)) u_mux_1155 (
        .y(_node_1040),
        .sel(_node_1039),
        .a(_T_1209_4),
        .b(_node_1038)
    );
    wire _node_1041;
    EQ_UNSIGNED #(.width(6)) u_eq_1156 (
        .y(_node_1041),
        .a(6'd5),
        .b(_T_1283)
    );
    wire _node_1042;
    MUX_UNSIGNED #(.width(1)) u_mux_1157 (
        .y(_node_1042),
        .sel(_node_1041),
        .a(_T_1209_5),
        .b(_node_1040)
    );
    wire _node_1043;
    EQ_UNSIGNED #(.width(6)) u_eq_1158 (
        .y(_node_1043),
        .a(6'd6),
        .b(_T_1283)
    );
    wire _node_1044;
    MUX_UNSIGNED #(.width(1)) u_mux_1159 (
        .y(_node_1044),
        .sel(_node_1043),
        .a(_T_1209_6),
        .b(_node_1042)
    );
    wire _node_1045;
    EQ_UNSIGNED #(.width(6)) u_eq_1160 (
        .y(_node_1045),
        .a(6'd7),
        .b(_T_1283)
    );
    wire _node_1046;
    MUX_UNSIGNED #(.width(1)) u_mux_1161 (
        .y(_node_1046),
        .sel(_node_1045),
        .a(_T_1209_7),
        .b(_node_1044)
    );
    wire _node_1047;
    EQ_UNSIGNED #(.width(6)) u_eq_1162 (
        .y(_node_1047),
        .a(6'd8),
        .b(_T_1283)
    );
    wire _node_1048;
    MUX_UNSIGNED #(.width(1)) u_mux_1163 (
        .y(_node_1048),
        .sel(_node_1047),
        .a(_T_1209_8),
        .b(_node_1046)
    );
    wire _node_1049;
    EQ_UNSIGNED #(.width(6)) u_eq_1164 (
        .y(_node_1049),
        .a(6'd9),
        .b(_T_1283)
    );
    wire _node_1050;
    MUX_UNSIGNED #(.width(1)) u_mux_1165 (
        .y(_node_1050),
        .sel(_node_1049),
        .a(_T_1209_9),
        .b(_node_1048)
    );
    wire _node_1051;
    EQ_UNSIGNED #(.width(6)) u_eq_1166 (
        .y(_node_1051),
        .a(6'd10),
        .b(_T_1283)
    );
    wire _node_1052;
    MUX_UNSIGNED #(.width(1)) u_mux_1167 (
        .y(_node_1052),
        .sel(_node_1051),
        .a(_T_1209_10),
        .b(_node_1050)
    );
    wire _node_1053;
    EQ_UNSIGNED #(.width(6)) u_eq_1168 (
        .y(_node_1053),
        .a(6'd11),
        .b(_T_1283)
    );
    wire _node_1054;
    MUX_UNSIGNED #(.width(1)) u_mux_1169 (
        .y(_node_1054),
        .sel(_node_1053),
        .a(_T_1209_11),
        .b(_node_1052)
    );
    wire _node_1055;
    EQ_UNSIGNED #(.width(6)) u_eq_1170 (
        .y(_node_1055),
        .a(6'd12),
        .b(_T_1283)
    );
    wire _node_1056;
    MUX_UNSIGNED #(.width(1)) u_mux_1171 (
        .y(_node_1056),
        .sel(_node_1055),
        .a(_T_1209_12),
        .b(_node_1054)
    );
    wire _node_1057;
    EQ_UNSIGNED #(.width(6)) u_eq_1172 (
        .y(_node_1057),
        .a(6'd13),
        .b(_T_1283)
    );
    wire _node_1058;
    MUX_UNSIGNED #(.width(1)) u_mux_1173 (
        .y(_node_1058),
        .sel(_node_1057),
        .a(_T_1209_13),
        .b(_node_1056)
    );
    wire _node_1059;
    EQ_UNSIGNED #(.width(6)) u_eq_1174 (
        .y(_node_1059),
        .a(6'd14),
        .b(_T_1283)
    );
    wire _node_1060;
    MUX_UNSIGNED #(.width(1)) u_mux_1175 (
        .y(_node_1060),
        .sel(_node_1059),
        .a(_T_1209_14),
        .b(_node_1058)
    );
    wire _node_1061;
    EQ_UNSIGNED #(.width(6)) u_eq_1176 (
        .y(_node_1061),
        .a(6'd15),
        .b(_T_1283)
    );
    wire _node_1062;
    MUX_UNSIGNED #(.width(1)) u_mux_1177 (
        .y(_node_1062),
        .sel(_node_1061),
        .a(_T_1209_15),
        .b(_node_1060)
    );
    wire _node_1063;
    EQ_UNSIGNED #(.width(6)) u_eq_1178 (
        .y(_node_1063),
        .a(6'd16),
        .b(_T_1283)
    );
    wire _node_1064;
    MUX_UNSIGNED #(.width(1)) u_mux_1179 (
        .y(_node_1064),
        .sel(_node_1063),
        .a(_T_1209_16),
        .b(_node_1062)
    );
    wire _node_1065;
    EQ_UNSIGNED #(.width(6)) u_eq_1180 (
        .y(_node_1065),
        .a(6'd17),
        .b(_T_1283)
    );
    wire _node_1066;
    MUX_UNSIGNED #(.width(1)) u_mux_1181 (
        .y(_node_1066),
        .sel(_node_1065),
        .a(_T_1209_17),
        .b(_node_1064)
    );
    wire _node_1067;
    EQ_UNSIGNED #(.width(6)) u_eq_1182 (
        .y(_node_1067),
        .a(6'd18),
        .b(_T_1283)
    );
    wire _node_1068;
    MUX_UNSIGNED #(.width(1)) u_mux_1183 (
        .y(_node_1068),
        .sel(_node_1067),
        .a(_T_1209_18),
        .b(_node_1066)
    );
    wire _node_1069;
    EQ_UNSIGNED #(.width(6)) u_eq_1184 (
        .y(_node_1069),
        .a(6'd19),
        .b(_T_1283)
    );
    wire _node_1070;
    MUX_UNSIGNED #(.width(1)) u_mux_1185 (
        .y(_node_1070),
        .sel(_node_1069),
        .a(_T_1209_19),
        .b(_node_1068)
    );
    wire _node_1071;
    EQ_UNSIGNED #(.width(6)) u_eq_1186 (
        .y(_node_1071),
        .a(6'd20),
        .b(_T_1283)
    );
    wire _node_1072;
    MUX_UNSIGNED #(.width(1)) u_mux_1187 (
        .y(_node_1072),
        .sel(_node_1071),
        .a(_T_1209_20),
        .b(_node_1070)
    );
    wire _node_1073;
    EQ_UNSIGNED #(.width(6)) u_eq_1188 (
        .y(_node_1073),
        .a(6'd21),
        .b(_T_1283)
    );
    wire _node_1074;
    MUX_UNSIGNED #(.width(1)) u_mux_1189 (
        .y(_node_1074),
        .sel(_node_1073),
        .a(_T_1209_21),
        .b(_node_1072)
    );
    wire _node_1075;
    EQ_UNSIGNED #(.width(6)) u_eq_1190 (
        .y(_node_1075),
        .a(6'd22),
        .b(_T_1283)
    );
    wire _node_1076;
    MUX_UNSIGNED #(.width(1)) u_mux_1191 (
        .y(_node_1076),
        .sel(_node_1075),
        .a(_T_1209_22),
        .b(_node_1074)
    );
    wire _node_1077;
    EQ_UNSIGNED #(.width(6)) u_eq_1192 (
        .y(_node_1077),
        .a(6'd23),
        .b(_T_1283)
    );
    wire _node_1078;
    MUX_UNSIGNED #(.width(1)) u_mux_1193 (
        .y(_node_1078),
        .sel(_node_1077),
        .a(_T_1209_23),
        .b(_node_1076)
    );
    wire _node_1079;
    EQ_UNSIGNED #(.width(6)) u_eq_1194 (
        .y(_node_1079),
        .a(6'd24),
        .b(_T_1283)
    );
    wire _node_1080;
    MUX_UNSIGNED #(.width(1)) u_mux_1195 (
        .y(_node_1080),
        .sel(_node_1079),
        .a(_T_1209_24),
        .b(_node_1078)
    );
    wire _node_1081;
    EQ_UNSIGNED #(.width(6)) u_eq_1196 (
        .y(_node_1081),
        .a(6'd25),
        .b(_T_1283)
    );
    wire _node_1082;
    MUX_UNSIGNED #(.width(1)) u_mux_1197 (
        .y(_node_1082),
        .sel(_node_1081),
        .a(_T_1209_25),
        .b(_node_1080)
    );
    wire _node_1083;
    EQ_UNSIGNED #(.width(6)) u_eq_1198 (
        .y(_node_1083),
        .a(6'd26),
        .b(_T_1283)
    );
    wire _node_1084;
    MUX_UNSIGNED #(.width(1)) u_mux_1199 (
        .y(_node_1084),
        .sel(_node_1083),
        .a(_T_1209_26),
        .b(_node_1082)
    );
    wire _node_1085;
    EQ_UNSIGNED #(.width(6)) u_eq_1200 (
        .y(_node_1085),
        .a(6'd27),
        .b(_T_1283)
    );
    wire _node_1086;
    MUX_UNSIGNED #(.width(1)) u_mux_1201 (
        .y(_node_1086),
        .sel(_node_1085),
        .a(_T_1209_27),
        .b(_node_1084)
    );
    wire _node_1087;
    EQ_UNSIGNED #(.width(6)) u_eq_1202 (
        .y(_node_1087),
        .a(6'd28),
        .b(_T_1283)
    );
    wire _node_1088;
    MUX_UNSIGNED #(.width(1)) u_mux_1203 (
        .y(_node_1088),
        .sel(_node_1087),
        .a(_T_1209_28),
        .b(_node_1086)
    );
    wire _node_1089;
    EQ_UNSIGNED #(.width(6)) u_eq_1204 (
        .y(_node_1089),
        .a(6'd29),
        .b(_T_1283)
    );
    wire _node_1090;
    MUX_UNSIGNED #(.width(1)) u_mux_1205 (
        .y(_node_1090),
        .sel(_node_1089),
        .a(_T_1209_29),
        .b(_node_1088)
    );
    wire _node_1091;
    EQ_UNSIGNED #(.width(6)) u_eq_1206 (
        .y(_node_1091),
        .a(6'd30),
        .b(_T_1283)
    );
    wire _node_1092;
    MUX_UNSIGNED #(.width(1)) u_mux_1207 (
        .y(_node_1092),
        .sel(_node_1091),
        .a(_T_1209_30),
        .b(_node_1090)
    );
    wire _node_1093;
    EQ_UNSIGNED #(.width(6)) u_eq_1208 (
        .y(_node_1093),
        .a(6'd31),
        .b(_T_1283)
    );
    wire _node_1094;
    MUX_UNSIGNED #(.width(1)) u_mux_1209 (
        .y(_node_1094),
        .sel(_node_1093),
        .a(_T_1209_31),
        .b(_node_1092)
    );
    wire _node_1095;
    EQ_UNSIGNED #(.width(6)) u_eq_1210 (
        .y(_node_1095),
        .a(6'd32),
        .b(_T_1283)
    );
    wire _node_1096;
    MUX_UNSIGNED #(.width(1)) u_mux_1211 (
        .y(_node_1096),
        .sel(_node_1095),
        .a(_T_1209_32),
        .b(_node_1094)
    );
    wire _node_1097;
    EQ_UNSIGNED #(.width(6)) u_eq_1212 (
        .y(_node_1097),
        .a(6'd33),
        .b(_T_1283)
    );
    wire _node_1098;
    MUX_UNSIGNED #(.width(1)) u_mux_1213 (
        .y(_node_1098),
        .sel(_node_1097),
        .a(_T_1209_33),
        .b(_node_1096)
    );
    wire _node_1099;
    EQ_UNSIGNED #(.width(6)) u_eq_1214 (
        .y(_node_1099),
        .a(6'd34),
        .b(_T_1283)
    );
    wire _node_1100;
    MUX_UNSIGNED #(.width(1)) u_mux_1215 (
        .y(_node_1100),
        .sel(_node_1099),
        .a(_T_1209_34),
        .b(_node_1098)
    );
    wire _node_1101;
    EQ_UNSIGNED #(.width(6)) u_eq_1216 (
        .y(_node_1101),
        .a(6'd35),
        .b(_T_1283)
    );
    wire _node_1102;
    MUX_UNSIGNED #(.width(1)) u_mux_1217 (
        .y(_node_1102),
        .sel(_node_1101),
        .a(_T_1209_35),
        .b(_node_1100)
    );
    wire _node_1103;
    EQ_UNSIGNED #(.width(6)) u_eq_1218 (
        .y(_node_1103),
        .a(6'd36),
        .b(_T_1283)
    );
    wire _node_1104;
    MUX_UNSIGNED #(.width(1)) u_mux_1219 (
        .y(_node_1104),
        .sel(_node_1103),
        .a(_T_1209_36),
        .b(_node_1102)
    );
    wire _node_1105;
    EQ_UNSIGNED #(.width(6)) u_eq_1220 (
        .y(_node_1105),
        .a(6'd37),
        .b(_T_1283)
    );
    wire _node_1106;
    MUX_UNSIGNED #(.width(1)) u_mux_1221 (
        .y(_node_1106),
        .sel(_node_1105),
        .a(_T_1209_37),
        .b(_node_1104)
    );
    wire _node_1107;
    EQ_UNSIGNED #(.width(6)) u_eq_1222 (
        .y(_node_1107),
        .a(6'd38),
        .b(_T_1283)
    );
    wire _node_1108;
    MUX_UNSIGNED #(.width(1)) u_mux_1223 (
        .y(_node_1108),
        .sel(_node_1107),
        .a(_T_1209_38),
        .b(_node_1106)
    );
    wire _node_1109;
    EQ_UNSIGNED #(.width(6)) u_eq_1224 (
        .y(_node_1109),
        .a(6'd39),
        .b(_T_1283)
    );
    wire _node_1110;
    MUX_UNSIGNED #(.width(1)) u_mux_1225 (
        .y(_node_1110),
        .sel(_node_1109),
        .a(_T_1209_39),
        .b(_node_1108)
    );
    wire _node_1111;
    EQ_UNSIGNED #(.width(6)) u_eq_1226 (
        .y(_node_1111),
        .a(6'd40),
        .b(_T_1283)
    );
    wire _node_1112;
    MUX_UNSIGNED #(.width(1)) u_mux_1227 (
        .y(_node_1112),
        .sel(_node_1111),
        .a(_T_1209_40),
        .b(_node_1110)
    );
    wire _node_1113;
    EQ_UNSIGNED #(.width(6)) u_eq_1228 (
        .y(_node_1113),
        .a(6'd41),
        .b(_T_1283)
    );
    wire _node_1114;
    MUX_UNSIGNED #(.width(1)) u_mux_1229 (
        .y(_node_1114),
        .sel(_node_1113),
        .a(_T_1209_41),
        .b(_node_1112)
    );
    wire _node_1115;
    EQ_UNSIGNED #(.width(6)) u_eq_1230 (
        .y(_node_1115),
        .a(6'd42),
        .b(_T_1283)
    );
    wire _node_1116;
    MUX_UNSIGNED #(.width(1)) u_mux_1231 (
        .y(_node_1116),
        .sel(_node_1115),
        .a(_T_1209_42),
        .b(_node_1114)
    );
    wire _node_1117;
    EQ_UNSIGNED #(.width(6)) u_eq_1232 (
        .y(_node_1117),
        .a(6'd43),
        .b(_T_1283)
    );
    wire _node_1118;
    MUX_UNSIGNED #(.width(1)) u_mux_1233 (
        .y(_node_1118),
        .sel(_node_1117),
        .a(_T_1209_43),
        .b(_node_1116)
    );
    wire _node_1119;
    EQ_UNSIGNED #(.width(6)) u_eq_1234 (
        .y(_node_1119),
        .a(6'd44),
        .b(_T_1283)
    );
    wire _node_1120;
    MUX_UNSIGNED #(.width(1)) u_mux_1235 (
        .y(_node_1120),
        .sel(_node_1119),
        .a(_T_1209_44),
        .b(_node_1118)
    );
    wire _node_1121;
    EQ_UNSIGNED #(.width(6)) u_eq_1236 (
        .y(_node_1121),
        .a(6'd45),
        .b(_T_1283)
    );
    wire _node_1122;
    MUX_UNSIGNED #(.width(1)) u_mux_1237 (
        .y(_node_1122),
        .sel(_node_1121),
        .a(_T_1209_45),
        .b(_node_1120)
    );
    wire _node_1123;
    EQ_UNSIGNED #(.width(6)) u_eq_1238 (
        .y(_node_1123),
        .a(6'd46),
        .b(_T_1283)
    );
    wire _node_1124;
    MUX_UNSIGNED #(.width(1)) u_mux_1239 (
        .y(_node_1124),
        .sel(_node_1123),
        .a(_T_1209_46),
        .b(_node_1122)
    );
    wire _node_1125;
    EQ_UNSIGNED #(.width(6)) u_eq_1240 (
        .y(_node_1125),
        .a(6'd47),
        .b(_T_1283)
    );
    wire _node_1126;
    MUX_UNSIGNED #(.width(1)) u_mux_1241 (
        .y(_node_1126),
        .sel(_node_1125),
        .a(_T_1209_47),
        .b(_node_1124)
    );
    wire _node_1127;
    EQ_UNSIGNED #(.width(6)) u_eq_1242 (
        .y(_node_1127),
        .a(6'd48),
        .b(_T_1283)
    );
    wire _node_1128;
    MUX_UNSIGNED #(.width(1)) u_mux_1243 (
        .y(_node_1128),
        .sel(_node_1127),
        .a(_T_1209_48),
        .b(_node_1126)
    );
    wire _node_1129;
    EQ_UNSIGNED #(.width(6)) u_eq_1244 (
        .y(_node_1129),
        .a(6'd49),
        .b(_T_1283)
    );
    wire _node_1130;
    MUX_UNSIGNED #(.width(1)) u_mux_1245 (
        .y(_node_1130),
        .sel(_node_1129),
        .a(_T_1209_49),
        .b(_node_1128)
    );
    wire _node_1131;
    EQ_UNSIGNED #(.width(6)) u_eq_1246 (
        .y(_node_1131),
        .a(6'd50),
        .b(_T_1283)
    );
    wire _node_1132;
    MUX_UNSIGNED #(.width(1)) u_mux_1247 (
        .y(_node_1132),
        .sel(_node_1131),
        .a(_T_1209_50),
        .b(_node_1130)
    );
    wire _node_1133;
    EQ_UNSIGNED #(.width(6)) u_eq_1248 (
        .y(_node_1133),
        .a(6'd51),
        .b(_T_1283)
    );
    wire _node_1134;
    MUX_UNSIGNED #(.width(1)) u_mux_1249 (
        .y(_node_1134),
        .sel(_node_1133),
        .a(_T_1209_51),
        .b(_node_1132)
    );
    wire _node_1135;
    EQ_UNSIGNED #(.width(6)) u_eq_1250 (
        .y(_node_1135),
        .a(6'd52),
        .b(_T_1283)
    );
    wire _node_1136;
    MUX_UNSIGNED #(.width(1)) u_mux_1251 (
        .y(_node_1136),
        .sel(_node_1135),
        .a(_T_1209_52),
        .b(_node_1134)
    );
    wire _T_1284;
    BITWISEAND #(.width(1)) bitwiseand_1252 (
        .y(_T_1284),
        .a(_c__io_outs_0_ready),
        .b(_c__io_outs_0_valid)
    );
    wire [2:0] _T_1286;
    BITS #(.width(6), .high(2), .low(0)) bits_1253 (
        .y(_T_1286),
        .in(_value_6__q)
    );
    wire _T_1288;
    EQ_UNSIGNED #(.width(1)) u_eq_1254 (
        .y(_T_1288),
        .a(reset),
        .b(1'h0)
    );
    wire [2:0] _T_1290;
    BITS #(.width(6), .high(2), .low(0)) bits_1255 (
        .y(_T_1290),
        .in(_value_6__q)
    );
    wire _node_1137;
    EQ_UNSIGNED #(.width(3)) u_eq_1256 (
        .y(_node_1137),
        .a(3'd0),
        .b(_T_1290)
    );
    wire [28:0] _node_1138;
    assign _node_1138 = _T_1274_0;
    wire _node_1139;
    EQ_UNSIGNED #(.width(3)) u_eq_1257 (
        .y(_node_1139),
        .a(3'd1),
        .b(_T_1290)
    );
    wire [28:0] _node_1140;
    MUX_UNSIGNED #(.width(29)) u_mux_1258 (
        .y(_node_1140),
        .sel(_node_1139),
        .a(_T_1274_1),
        .b(_node_1138)
    );
    wire _node_1141;
    EQ_UNSIGNED #(.width(3)) u_eq_1259 (
        .y(_node_1141),
        .a(3'd2),
        .b(_T_1290)
    );
    wire [28:0] _node_1142;
    MUX_UNSIGNED #(.width(29)) u_mux_1260 (
        .y(_node_1142),
        .sel(_node_1141),
        .a(_T_1274_2),
        .b(_node_1140)
    );
    wire _node_1143;
    EQ_UNSIGNED #(.width(3)) u_eq_1261 (
        .y(_node_1143),
        .a(3'd3),
        .b(_T_1290)
    );
    wire [28:0] _node_1144;
    MUX_UNSIGNED #(.width(29)) u_mux_1262 (
        .y(_node_1144),
        .sel(_node_1143),
        .a(_T_1274_3),
        .b(_node_1142)
    );
    wire _node_1145;
    EQ_UNSIGNED #(.width(3)) u_eq_1263 (
        .y(_node_1145),
        .a(3'd4),
        .b(_T_1290)
    );
    wire [28:0] _node_1146;
    MUX_UNSIGNED #(.width(29)) u_mux_1264 (
        .y(_node_1146),
        .sel(_node_1145),
        .a(_T_1274_4),
        .b(_node_1144)
    );
    wire _T_1291;
    wire [63:0] _WTEMP_44;
    PAD_UNSIGNED #(.width(29), .n(64)) u_pad_1265 (
        .y(_WTEMP_44),
        .in(_node_1146)
    );
    NEQ_UNSIGNED #(.width(64)) u_neq_1266 (
        .y(_T_1291),
        .a(_c__io_outs_0_bits_body),
        .b(_WTEMP_44)
    );
    wire [2:0] _T_1293;
    BITS #(.width(6), .high(2), .low(0)) bits_1267 (
        .y(_T_1293),
        .in(_value_6__q)
    );
    wire _T_1295;
    EQ_UNSIGNED #(.width(1)) u_eq_1268 (
        .y(_T_1295),
        .a(reset),
        .b(1'h0)
    );
    wire _T_1297;
    BITWISEOR #(.width(1)) bitwiseor_1269 (
        .y(_T_1297),
        .a(1'h0),
        .b(reset)
    );
    wire _T_1299;
    EQ_UNSIGNED #(.width(1)) u_eq_1270 (
        .y(_T_1299),
        .a(_T_1297),
        .b(1'h0)
    );
    wire _T_1301;
    EQ_UNSIGNED #(.width(1)) u_eq_1271 (
        .y(_T_1301),
        .a(reset),
        .b(1'h0)
    );
    wire _T_1303;
    EQ_UNSIGNED #(.width(6)) u_eq_1272 (
        .y(_T_1303),
        .a(_value_6__q),
        .b(6'h20)
    );
    wire [6:0] _T_1305;
    wire [5:0] _WTEMP_45;
    PAD_UNSIGNED #(.width(1), .n(6)) u_pad_1273 (
        .y(_WTEMP_45),
        .in(1'h1)
    );
    ADD_UNSIGNED #(.width(6)) u_add_1274 (
        .y(_T_1305),
        .a(_value_6__q),
        .b(_WTEMP_45)
    );
    wire [5:0] _T_1306;
    TAIL #(.width(7), .n(1)) tail_1275 (
        .y(_T_1306),
        .in(_T_1305)
    );
    wire _T_1309;
    EQ_UNSIGNED #(.width(1)) u_eq_1276 (
        .y(_T_1309),
        .a(__T_13__q),
        .b(1'h0)
    );
    wire _T_1311;
    wire [7:0] _WTEMP_46;
    PAD_UNSIGNED #(.width(6), .n(8)) u_pad_1277 (
        .y(_WTEMP_46),
        .in(6'h20)
    );
    EQ_UNSIGNED #(.width(8)) u_eq_1278 (
        .y(_T_1311),
        .a(__T_10__q),
        .b(_WTEMP_46)
    );
    wire _node_1147;
    MUX_UNSIGNED #(.width(1)) u_mux_1279 (
        .y(_node_1147),
        .sel(_T_1122),
        .a(_node_1028),
        .b(_node_1029)
    );
    wire [8:0] _T_1314;
    wire [7:0] _WTEMP_47;
    PAD_UNSIGNED #(.width(1), .n(8)) u_pad_1280 (
        .y(_WTEMP_47),
        .in(1'h1)
    );
    ADD_UNSIGNED #(.width(8)) u_add_1281 (
        .y(_T_1314),
        .a(__T_10__q),
        .b(_WTEMP_47)
    );
    wire [7:0] _T_1315;
    TAIL #(.width(9), .n(1)) tail_1282 (
        .y(_T_1315),
        .in(_T_1314)
    );
    wire [7:0] _node_1148;
    MUX_UNSIGNED #(.width(8)) u_mux_1283 (
        .y(_node_1148),
        .sel(_T_1122),
        .a(_node_1026),
        .b(_node_1027)
    );
    wire _node_1149;
    MUX_UNSIGNED #(.width(1)) u_mux_1284 (
        .y(_node_1149),
        .sel(_T_1311),
        .a(1'h1),
        .b(_node_1147)
    );
    wire _node_1150;
    MUX_UNSIGNED #(.width(1)) u_mux_1285 (
        .y(_node_1150),
        .sel(_T_1122),
        .a(_node_1028),
        .b(_node_1029)
    );
    wire [7:0] _node_1151;
    MUX_UNSIGNED #(.width(8)) u_mux_1286 (
        .y(_node_1151),
        .sel(_T_1309),
        .a(_T_1315),
        .b(_node_1148)
    );
    wire [7:0] _node_1152;
    MUX_UNSIGNED #(.width(8)) u_mux_1287 (
        .y(_node_1152),
        .sel(_T_1122),
        .a(_node_1026),
        .b(_node_1027)
    );
    wire _node_1153;
    MUX_UNSIGNED #(.width(1)) u_mux_1288 (
        .y(_node_1153),
        .sel(_T_1309),
        .a(_node_1149),
        .b(_node_1150)
    );
    wire _node_1154;
    MUX_UNSIGNED #(.width(1)) u_mux_1289 (
        .y(_node_1154),
        .sel(_T_1122),
        .a(_node_1028),
        .b(_node_1029)
    );
    wire [5:0] _node_1155;
    wire [5:0] _WTEMP_48;
    PAD_UNSIGNED #(.width(1), .n(6)) u_pad_1290 (
        .y(_WTEMP_48),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(6)) u_mux_1291 (
        .y(_node_1155),
        .sel(_T_1303),
        .a(_WTEMP_48),
        .b(_T_1306)
    );
    wire _T_1371_0;
    wire _T_1371_1;
    wire _T_1371_2;
    wire _T_1371_3;
    wire _T_1371_4;
    wire _T_1371_5;
    wire _T_1371_6;
    wire _T_1371_7;
    wire _T_1371_8;
    wire _T_1371_9;
    wire _T_1371_10;
    wire _T_1371_11;
    wire _T_1371_12;
    wire _T_1371_13;
    wire _T_1371_14;
    wire _T_1371_15;
    wire _T_1371_16;
    wire _T_1371_17;
    wire _T_1371_18;
    wire _T_1371_19;
    wire _T_1371_20;
    wire _T_1371_21;
    wire _T_1371_22;
    wire _T_1371_23;
    wire _T_1371_24;
    wire _T_1371_25;
    wire _T_1371_26;
    wire _T_1371_27;
    wire _T_1371_28;
    wire _T_1371_29;
    wire _T_1371_30;
    wire _T_1371_31;
    wire _T_1371_32;
    wire _T_1371_33;
    wire _T_1371_34;
    wire _T_1371_35;
    wire _T_1371_36;
    wire _T_1371_37;
    wire _T_1371_38;
    wire _T_1371_39;
    wire _T_1371_40;
    wire _T_1371_41;
    wire _T_1371_42;
    wire _T_1371_43;
    wire _T_1371_44;
    wire _T_1371_45;
    wire _T_1371_46;
    wire _T_1371_47;
    wire _T_1371_48;
    wire _T_1371_49;
    wire _T_1371_50;
    wire _T_1371_51;
    wire _T_1371_52;
    wire [5:0] _value_7__q;
    wire [5:0] _value_7__d;
    DFF_POSCLK #(.width(6)) value_7 (
        .q(_value_7__q),
        .d(_value_7__d),
        .clk(clock)
    );
    wire [5:0] _WTEMP_49;
    MUX_UNSIGNED #(.width(6)) u_mux_1292 (
        .y(_value_7__d),
        .sel(reset),
        .a(6'h0),
        .b(_WTEMP_49)
    );
    wire [1:0] _T_1441_0;
    wire [1:0] _T_1441_1;
    wire [1:0] _T_1441_2;
    wire [1:0] _T_1441_3;
    wire [1:0] _T_1441_4;
    wire [1:0] _T_1441_5;
    wire [1:0] _T_1441_6;
    wire [1:0] _T_1441_7;
    wire [1:0] _T_1441_8;
    wire [1:0] _T_1441_9;
    wire [5:0] _T_1455;
    BITS #(.width(8), .high(5), .low(0)) bits_1293 (
        .y(_T_1455),
        .in(__T_10__q)
    );
    wire _node_1156;
    EQ_UNSIGNED #(.width(6)) u_eq_1294 (
        .y(_node_1156),
        .a(6'd0),
        .b(_T_1455)
    );
    wire _node_1157;
    assign _node_1157 = _T_1371_0;
    wire _node_1158;
    EQ_UNSIGNED #(.width(6)) u_eq_1295 (
        .y(_node_1158),
        .a(6'd1),
        .b(_T_1455)
    );
    wire _node_1159;
    MUX_UNSIGNED #(.width(1)) u_mux_1296 (
        .y(_node_1159),
        .sel(_node_1158),
        .a(_T_1371_1),
        .b(_node_1157)
    );
    wire _node_1160;
    EQ_UNSIGNED #(.width(6)) u_eq_1297 (
        .y(_node_1160),
        .a(6'd2),
        .b(_T_1455)
    );
    wire _node_1161;
    MUX_UNSIGNED #(.width(1)) u_mux_1298 (
        .y(_node_1161),
        .sel(_node_1160),
        .a(_T_1371_2),
        .b(_node_1159)
    );
    wire _node_1162;
    EQ_UNSIGNED #(.width(6)) u_eq_1299 (
        .y(_node_1162),
        .a(6'd3),
        .b(_T_1455)
    );
    wire _node_1163;
    MUX_UNSIGNED #(.width(1)) u_mux_1300 (
        .y(_node_1163),
        .sel(_node_1162),
        .a(_T_1371_3),
        .b(_node_1161)
    );
    wire _node_1164;
    EQ_UNSIGNED #(.width(6)) u_eq_1301 (
        .y(_node_1164),
        .a(6'd4),
        .b(_T_1455)
    );
    wire _node_1165;
    MUX_UNSIGNED #(.width(1)) u_mux_1302 (
        .y(_node_1165),
        .sel(_node_1164),
        .a(_T_1371_4),
        .b(_node_1163)
    );
    wire _node_1166;
    EQ_UNSIGNED #(.width(6)) u_eq_1303 (
        .y(_node_1166),
        .a(6'd5),
        .b(_T_1455)
    );
    wire _node_1167;
    MUX_UNSIGNED #(.width(1)) u_mux_1304 (
        .y(_node_1167),
        .sel(_node_1166),
        .a(_T_1371_5),
        .b(_node_1165)
    );
    wire _node_1168;
    EQ_UNSIGNED #(.width(6)) u_eq_1305 (
        .y(_node_1168),
        .a(6'd6),
        .b(_T_1455)
    );
    wire _node_1169;
    MUX_UNSIGNED #(.width(1)) u_mux_1306 (
        .y(_node_1169),
        .sel(_node_1168),
        .a(_T_1371_6),
        .b(_node_1167)
    );
    wire _node_1170;
    EQ_UNSIGNED #(.width(6)) u_eq_1307 (
        .y(_node_1170),
        .a(6'd7),
        .b(_T_1455)
    );
    wire _node_1171;
    MUX_UNSIGNED #(.width(1)) u_mux_1308 (
        .y(_node_1171),
        .sel(_node_1170),
        .a(_T_1371_7),
        .b(_node_1169)
    );
    wire _node_1172;
    EQ_UNSIGNED #(.width(6)) u_eq_1309 (
        .y(_node_1172),
        .a(6'd8),
        .b(_T_1455)
    );
    wire _node_1173;
    MUX_UNSIGNED #(.width(1)) u_mux_1310 (
        .y(_node_1173),
        .sel(_node_1172),
        .a(_T_1371_8),
        .b(_node_1171)
    );
    wire _node_1174;
    EQ_UNSIGNED #(.width(6)) u_eq_1311 (
        .y(_node_1174),
        .a(6'd9),
        .b(_T_1455)
    );
    wire _node_1175;
    MUX_UNSIGNED #(.width(1)) u_mux_1312 (
        .y(_node_1175),
        .sel(_node_1174),
        .a(_T_1371_9),
        .b(_node_1173)
    );
    wire _node_1176;
    EQ_UNSIGNED #(.width(6)) u_eq_1313 (
        .y(_node_1176),
        .a(6'd10),
        .b(_T_1455)
    );
    wire _node_1177;
    MUX_UNSIGNED #(.width(1)) u_mux_1314 (
        .y(_node_1177),
        .sel(_node_1176),
        .a(_T_1371_10),
        .b(_node_1175)
    );
    wire _node_1178;
    EQ_UNSIGNED #(.width(6)) u_eq_1315 (
        .y(_node_1178),
        .a(6'd11),
        .b(_T_1455)
    );
    wire _node_1179;
    MUX_UNSIGNED #(.width(1)) u_mux_1316 (
        .y(_node_1179),
        .sel(_node_1178),
        .a(_T_1371_11),
        .b(_node_1177)
    );
    wire _node_1180;
    EQ_UNSIGNED #(.width(6)) u_eq_1317 (
        .y(_node_1180),
        .a(6'd12),
        .b(_T_1455)
    );
    wire _node_1181;
    MUX_UNSIGNED #(.width(1)) u_mux_1318 (
        .y(_node_1181),
        .sel(_node_1180),
        .a(_T_1371_12),
        .b(_node_1179)
    );
    wire _node_1182;
    EQ_UNSIGNED #(.width(6)) u_eq_1319 (
        .y(_node_1182),
        .a(6'd13),
        .b(_T_1455)
    );
    wire _node_1183;
    MUX_UNSIGNED #(.width(1)) u_mux_1320 (
        .y(_node_1183),
        .sel(_node_1182),
        .a(_T_1371_13),
        .b(_node_1181)
    );
    wire _node_1184;
    EQ_UNSIGNED #(.width(6)) u_eq_1321 (
        .y(_node_1184),
        .a(6'd14),
        .b(_T_1455)
    );
    wire _node_1185;
    MUX_UNSIGNED #(.width(1)) u_mux_1322 (
        .y(_node_1185),
        .sel(_node_1184),
        .a(_T_1371_14),
        .b(_node_1183)
    );
    wire _node_1186;
    EQ_UNSIGNED #(.width(6)) u_eq_1323 (
        .y(_node_1186),
        .a(6'd15),
        .b(_T_1455)
    );
    wire _node_1187;
    MUX_UNSIGNED #(.width(1)) u_mux_1324 (
        .y(_node_1187),
        .sel(_node_1186),
        .a(_T_1371_15),
        .b(_node_1185)
    );
    wire _node_1188;
    EQ_UNSIGNED #(.width(6)) u_eq_1325 (
        .y(_node_1188),
        .a(6'd16),
        .b(_T_1455)
    );
    wire _node_1189;
    MUX_UNSIGNED #(.width(1)) u_mux_1326 (
        .y(_node_1189),
        .sel(_node_1188),
        .a(_T_1371_16),
        .b(_node_1187)
    );
    wire _node_1190;
    EQ_UNSIGNED #(.width(6)) u_eq_1327 (
        .y(_node_1190),
        .a(6'd17),
        .b(_T_1455)
    );
    wire _node_1191;
    MUX_UNSIGNED #(.width(1)) u_mux_1328 (
        .y(_node_1191),
        .sel(_node_1190),
        .a(_T_1371_17),
        .b(_node_1189)
    );
    wire _node_1192;
    EQ_UNSIGNED #(.width(6)) u_eq_1329 (
        .y(_node_1192),
        .a(6'd18),
        .b(_T_1455)
    );
    wire _node_1193;
    MUX_UNSIGNED #(.width(1)) u_mux_1330 (
        .y(_node_1193),
        .sel(_node_1192),
        .a(_T_1371_18),
        .b(_node_1191)
    );
    wire _node_1194;
    EQ_UNSIGNED #(.width(6)) u_eq_1331 (
        .y(_node_1194),
        .a(6'd19),
        .b(_T_1455)
    );
    wire _node_1195;
    MUX_UNSIGNED #(.width(1)) u_mux_1332 (
        .y(_node_1195),
        .sel(_node_1194),
        .a(_T_1371_19),
        .b(_node_1193)
    );
    wire _node_1196;
    EQ_UNSIGNED #(.width(6)) u_eq_1333 (
        .y(_node_1196),
        .a(6'd20),
        .b(_T_1455)
    );
    wire _node_1197;
    MUX_UNSIGNED #(.width(1)) u_mux_1334 (
        .y(_node_1197),
        .sel(_node_1196),
        .a(_T_1371_20),
        .b(_node_1195)
    );
    wire _node_1198;
    EQ_UNSIGNED #(.width(6)) u_eq_1335 (
        .y(_node_1198),
        .a(6'd21),
        .b(_T_1455)
    );
    wire _node_1199;
    MUX_UNSIGNED #(.width(1)) u_mux_1336 (
        .y(_node_1199),
        .sel(_node_1198),
        .a(_T_1371_21),
        .b(_node_1197)
    );
    wire _node_1200;
    EQ_UNSIGNED #(.width(6)) u_eq_1337 (
        .y(_node_1200),
        .a(6'd22),
        .b(_T_1455)
    );
    wire _node_1201;
    MUX_UNSIGNED #(.width(1)) u_mux_1338 (
        .y(_node_1201),
        .sel(_node_1200),
        .a(_T_1371_22),
        .b(_node_1199)
    );
    wire _node_1202;
    EQ_UNSIGNED #(.width(6)) u_eq_1339 (
        .y(_node_1202),
        .a(6'd23),
        .b(_T_1455)
    );
    wire _node_1203;
    MUX_UNSIGNED #(.width(1)) u_mux_1340 (
        .y(_node_1203),
        .sel(_node_1202),
        .a(_T_1371_23),
        .b(_node_1201)
    );
    wire _node_1204;
    EQ_UNSIGNED #(.width(6)) u_eq_1341 (
        .y(_node_1204),
        .a(6'd24),
        .b(_T_1455)
    );
    wire _node_1205;
    MUX_UNSIGNED #(.width(1)) u_mux_1342 (
        .y(_node_1205),
        .sel(_node_1204),
        .a(_T_1371_24),
        .b(_node_1203)
    );
    wire _node_1206;
    EQ_UNSIGNED #(.width(6)) u_eq_1343 (
        .y(_node_1206),
        .a(6'd25),
        .b(_T_1455)
    );
    wire _node_1207;
    MUX_UNSIGNED #(.width(1)) u_mux_1344 (
        .y(_node_1207),
        .sel(_node_1206),
        .a(_T_1371_25),
        .b(_node_1205)
    );
    wire _node_1208;
    EQ_UNSIGNED #(.width(6)) u_eq_1345 (
        .y(_node_1208),
        .a(6'd26),
        .b(_T_1455)
    );
    wire _node_1209;
    MUX_UNSIGNED #(.width(1)) u_mux_1346 (
        .y(_node_1209),
        .sel(_node_1208),
        .a(_T_1371_26),
        .b(_node_1207)
    );
    wire _node_1210;
    EQ_UNSIGNED #(.width(6)) u_eq_1347 (
        .y(_node_1210),
        .a(6'd27),
        .b(_T_1455)
    );
    wire _node_1211;
    MUX_UNSIGNED #(.width(1)) u_mux_1348 (
        .y(_node_1211),
        .sel(_node_1210),
        .a(_T_1371_27),
        .b(_node_1209)
    );
    wire _node_1212;
    EQ_UNSIGNED #(.width(6)) u_eq_1349 (
        .y(_node_1212),
        .a(6'd28),
        .b(_T_1455)
    );
    wire _node_1213;
    MUX_UNSIGNED #(.width(1)) u_mux_1350 (
        .y(_node_1213),
        .sel(_node_1212),
        .a(_T_1371_28),
        .b(_node_1211)
    );
    wire _node_1214;
    EQ_UNSIGNED #(.width(6)) u_eq_1351 (
        .y(_node_1214),
        .a(6'd29),
        .b(_T_1455)
    );
    wire _node_1215;
    MUX_UNSIGNED #(.width(1)) u_mux_1352 (
        .y(_node_1215),
        .sel(_node_1214),
        .a(_T_1371_29),
        .b(_node_1213)
    );
    wire _node_1216;
    EQ_UNSIGNED #(.width(6)) u_eq_1353 (
        .y(_node_1216),
        .a(6'd30),
        .b(_T_1455)
    );
    wire _node_1217;
    MUX_UNSIGNED #(.width(1)) u_mux_1354 (
        .y(_node_1217),
        .sel(_node_1216),
        .a(_T_1371_30),
        .b(_node_1215)
    );
    wire _node_1218;
    EQ_UNSIGNED #(.width(6)) u_eq_1355 (
        .y(_node_1218),
        .a(6'd31),
        .b(_T_1455)
    );
    wire _node_1219;
    MUX_UNSIGNED #(.width(1)) u_mux_1356 (
        .y(_node_1219),
        .sel(_node_1218),
        .a(_T_1371_31),
        .b(_node_1217)
    );
    wire _node_1220;
    EQ_UNSIGNED #(.width(6)) u_eq_1357 (
        .y(_node_1220),
        .a(6'd32),
        .b(_T_1455)
    );
    wire _node_1221;
    MUX_UNSIGNED #(.width(1)) u_mux_1358 (
        .y(_node_1221),
        .sel(_node_1220),
        .a(_T_1371_32),
        .b(_node_1219)
    );
    wire _node_1222;
    EQ_UNSIGNED #(.width(6)) u_eq_1359 (
        .y(_node_1222),
        .a(6'd33),
        .b(_T_1455)
    );
    wire _node_1223;
    MUX_UNSIGNED #(.width(1)) u_mux_1360 (
        .y(_node_1223),
        .sel(_node_1222),
        .a(_T_1371_33),
        .b(_node_1221)
    );
    wire _node_1224;
    EQ_UNSIGNED #(.width(6)) u_eq_1361 (
        .y(_node_1224),
        .a(6'd34),
        .b(_T_1455)
    );
    wire _node_1225;
    MUX_UNSIGNED #(.width(1)) u_mux_1362 (
        .y(_node_1225),
        .sel(_node_1224),
        .a(_T_1371_34),
        .b(_node_1223)
    );
    wire _node_1226;
    EQ_UNSIGNED #(.width(6)) u_eq_1363 (
        .y(_node_1226),
        .a(6'd35),
        .b(_T_1455)
    );
    wire _node_1227;
    MUX_UNSIGNED #(.width(1)) u_mux_1364 (
        .y(_node_1227),
        .sel(_node_1226),
        .a(_T_1371_35),
        .b(_node_1225)
    );
    wire _node_1228;
    EQ_UNSIGNED #(.width(6)) u_eq_1365 (
        .y(_node_1228),
        .a(6'd36),
        .b(_T_1455)
    );
    wire _node_1229;
    MUX_UNSIGNED #(.width(1)) u_mux_1366 (
        .y(_node_1229),
        .sel(_node_1228),
        .a(_T_1371_36),
        .b(_node_1227)
    );
    wire _node_1230;
    EQ_UNSIGNED #(.width(6)) u_eq_1367 (
        .y(_node_1230),
        .a(6'd37),
        .b(_T_1455)
    );
    wire _node_1231;
    MUX_UNSIGNED #(.width(1)) u_mux_1368 (
        .y(_node_1231),
        .sel(_node_1230),
        .a(_T_1371_37),
        .b(_node_1229)
    );
    wire _node_1232;
    EQ_UNSIGNED #(.width(6)) u_eq_1369 (
        .y(_node_1232),
        .a(6'd38),
        .b(_T_1455)
    );
    wire _node_1233;
    MUX_UNSIGNED #(.width(1)) u_mux_1370 (
        .y(_node_1233),
        .sel(_node_1232),
        .a(_T_1371_38),
        .b(_node_1231)
    );
    wire _node_1234;
    EQ_UNSIGNED #(.width(6)) u_eq_1371 (
        .y(_node_1234),
        .a(6'd39),
        .b(_T_1455)
    );
    wire _node_1235;
    MUX_UNSIGNED #(.width(1)) u_mux_1372 (
        .y(_node_1235),
        .sel(_node_1234),
        .a(_T_1371_39),
        .b(_node_1233)
    );
    wire _node_1236;
    EQ_UNSIGNED #(.width(6)) u_eq_1373 (
        .y(_node_1236),
        .a(6'd40),
        .b(_T_1455)
    );
    wire _node_1237;
    MUX_UNSIGNED #(.width(1)) u_mux_1374 (
        .y(_node_1237),
        .sel(_node_1236),
        .a(_T_1371_40),
        .b(_node_1235)
    );
    wire _node_1238;
    EQ_UNSIGNED #(.width(6)) u_eq_1375 (
        .y(_node_1238),
        .a(6'd41),
        .b(_T_1455)
    );
    wire _node_1239;
    MUX_UNSIGNED #(.width(1)) u_mux_1376 (
        .y(_node_1239),
        .sel(_node_1238),
        .a(_T_1371_41),
        .b(_node_1237)
    );
    wire _node_1240;
    EQ_UNSIGNED #(.width(6)) u_eq_1377 (
        .y(_node_1240),
        .a(6'd42),
        .b(_T_1455)
    );
    wire _node_1241;
    MUX_UNSIGNED #(.width(1)) u_mux_1378 (
        .y(_node_1241),
        .sel(_node_1240),
        .a(_T_1371_42),
        .b(_node_1239)
    );
    wire _node_1242;
    EQ_UNSIGNED #(.width(6)) u_eq_1379 (
        .y(_node_1242),
        .a(6'd43),
        .b(_T_1455)
    );
    wire _node_1243;
    MUX_UNSIGNED #(.width(1)) u_mux_1380 (
        .y(_node_1243),
        .sel(_node_1242),
        .a(_T_1371_43),
        .b(_node_1241)
    );
    wire _node_1244;
    EQ_UNSIGNED #(.width(6)) u_eq_1381 (
        .y(_node_1244),
        .a(6'd44),
        .b(_T_1455)
    );
    wire _node_1245;
    MUX_UNSIGNED #(.width(1)) u_mux_1382 (
        .y(_node_1245),
        .sel(_node_1244),
        .a(_T_1371_44),
        .b(_node_1243)
    );
    wire _node_1246;
    EQ_UNSIGNED #(.width(6)) u_eq_1383 (
        .y(_node_1246),
        .a(6'd45),
        .b(_T_1455)
    );
    wire _node_1247;
    MUX_UNSIGNED #(.width(1)) u_mux_1384 (
        .y(_node_1247),
        .sel(_node_1246),
        .a(_T_1371_45),
        .b(_node_1245)
    );
    wire _node_1248;
    EQ_UNSIGNED #(.width(6)) u_eq_1385 (
        .y(_node_1248),
        .a(6'd46),
        .b(_T_1455)
    );
    wire _node_1249;
    MUX_UNSIGNED #(.width(1)) u_mux_1386 (
        .y(_node_1249),
        .sel(_node_1248),
        .a(_T_1371_46),
        .b(_node_1247)
    );
    wire _node_1250;
    EQ_UNSIGNED #(.width(6)) u_eq_1387 (
        .y(_node_1250),
        .a(6'd47),
        .b(_T_1455)
    );
    wire _node_1251;
    MUX_UNSIGNED #(.width(1)) u_mux_1388 (
        .y(_node_1251),
        .sel(_node_1250),
        .a(_T_1371_47),
        .b(_node_1249)
    );
    wire _node_1252;
    EQ_UNSIGNED #(.width(6)) u_eq_1389 (
        .y(_node_1252),
        .a(6'd48),
        .b(_T_1455)
    );
    wire _node_1253;
    MUX_UNSIGNED #(.width(1)) u_mux_1390 (
        .y(_node_1253),
        .sel(_node_1252),
        .a(_T_1371_48),
        .b(_node_1251)
    );
    wire _node_1254;
    EQ_UNSIGNED #(.width(6)) u_eq_1391 (
        .y(_node_1254),
        .a(6'd49),
        .b(_T_1455)
    );
    wire _node_1255;
    MUX_UNSIGNED #(.width(1)) u_mux_1392 (
        .y(_node_1255),
        .sel(_node_1254),
        .a(_T_1371_49),
        .b(_node_1253)
    );
    wire _node_1256;
    EQ_UNSIGNED #(.width(6)) u_eq_1393 (
        .y(_node_1256),
        .a(6'd50),
        .b(_T_1455)
    );
    wire _node_1257;
    MUX_UNSIGNED #(.width(1)) u_mux_1394 (
        .y(_node_1257),
        .sel(_node_1256),
        .a(_T_1371_50),
        .b(_node_1255)
    );
    wire _node_1258;
    EQ_UNSIGNED #(.width(6)) u_eq_1395 (
        .y(_node_1258),
        .a(6'd51),
        .b(_T_1455)
    );
    wire _node_1259;
    MUX_UNSIGNED #(.width(1)) u_mux_1396 (
        .y(_node_1259),
        .sel(_node_1258),
        .a(_T_1371_51),
        .b(_node_1257)
    );
    wire _node_1260;
    EQ_UNSIGNED #(.width(6)) u_eq_1397 (
        .y(_node_1260),
        .a(6'd52),
        .b(_T_1455)
    );
    wire _node_1261;
    MUX_UNSIGNED #(.width(1)) u_mux_1398 (
        .y(_node_1261),
        .sel(_node_1260),
        .a(_T_1371_52),
        .b(_node_1259)
    );
    wire _T_1456;
    BITWISEAND #(.width(1)) bitwiseand_1399 (
        .y(_T_1456),
        .a(_c__io_read_routing_table_response_ready),
        .b(_c__io_read_routing_table_response_valid)
    );
    wire [3:0] _T_1458;
    BITS #(.width(6), .high(3), .low(0)) bits_1400 (
        .y(_T_1458),
        .in(_value_7__q)
    );
    wire _T_1460;
    EQ_UNSIGNED #(.width(1)) u_eq_1401 (
        .y(_T_1460),
        .a(reset),
        .b(1'h0)
    );
    wire [3:0] _T_1462;
    BITS #(.width(6), .high(3), .low(0)) bits_1402 (
        .y(_T_1462),
        .in(_value_7__q)
    );
    wire _node_1262;
    EQ_UNSIGNED #(.width(4)) u_eq_1403 (
        .y(_node_1262),
        .a(4'd0),
        .b(_T_1462)
    );
    wire [1:0] _node_1263;
    assign _node_1263 = _T_1441_0;
    wire _node_1264;
    EQ_UNSIGNED #(.width(4)) u_eq_1404 (
        .y(_node_1264),
        .a(4'd1),
        .b(_T_1462)
    );
    wire [1:0] _node_1265;
    MUX_UNSIGNED #(.width(2)) u_mux_1405 (
        .y(_node_1265),
        .sel(_node_1264),
        .a(_T_1441_1),
        .b(_node_1263)
    );
    wire _node_1266;
    EQ_UNSIGNED #(.width(4)) u_eq_1406 (
        .y(_node_1266),
        .a(4'd2),
        .b(_T_1462)
    );
    wire [1:0] _node_1267;
    MUX_UNSIGNED #(.width(2)) u_mux_1407 (
        .y(_node_1267),
        .sel(_node_1266),
        .a(_T_1441_2),
        .b(_node_1265)
    );
    wire _node_1268;
    EQ_UNSIGNED #(.width(4)) u_eq_1408 (
        .y(_node_1268),
        .a(4'd3),
        .b(_T_1462)
    );
    wire [1:0] _node_1269;
    MUX_UNSIGNED #(.width(2)) u_mux_1409 (
        .y(_node_1269),
        .sel(_node_1268),
        .a(_T_1441_3),
        .b(_node_1267)
    );
    wire _node_1270;
    EQ_UNSIGNED #(.width(4)) u_eq_1410 (
        .y(_node_1270),
        .a(4'd4),
        .b(_T_1462)
    );
    wire [1:0] _node_1271;
    MUX_UNSIGNED #(.width(2)) u_mux_1411 (
        .y(_node_1271),
        .sel(_node_1270),
        .a(_T_1441_4),
        .b(_node_1269)
    );
    wire _node_1272;
    EQ_UNSIGNED #(.width(4)) u_eq_1412 (
        .y(_node_1272),
        .a(4'd5),
        .b(_T_1462)
    );
    wire [1:0] _node_1273;
    MUX_UNSIGNED #(.width(2)) u_mux_1413 (
        .y(_node_1273),
        .sel(_node_1272),
        .a(_T_1441_5),
        .b(_node_1271)
    );
    wire _node_1274;
    EQ_UNSIGNED #(.width(4)) u_eq_1414 (
        .y(_node_1274),
        .a(4'd6),
        .b(_T_1462)
    );
    wire [1:0] _node_1275;
    MUX_UNSIGNED #(.width(2)) u_mux_1415 (
        .y(_node_1275),
        .sel(_node_1274),
        .a(_T_1441_6),
        .b(_node_1273)
    );
    wire _node_1276;
    EQ_UNSIGNED #(.width(4)) u_eq_1416 (
        .y(_node_1276),
        .a(4'd7),
        .b(_T_1462)
    );
    wire [1:0] _node_1277;
    MUX_UNSIGNED #(.width(2)) u_mux_1417 (
        .y(_node_1277),
        .sel(_node_1276),
        .a(_T_1441_7),
        .b(_node_1275)
    );
    wire _node_1278;
    EQ_UNSIGNED #(.width(4)) u_eq_1418 (
        .y(_node_1278),
        .a(4'd8),
        .b(_T_1462)
    );
    wire [1:0] _node_1279;
    MUX_UNSIGNED #(.width(2)) u_mux_1419 (
        .y(_node_1279),
        .sel(_node_1278),
        .a(_T_1441_8),
        .b(_node_1277)
    );
    wire _node_1280;
    EQ_UNSIGNED #(.width(4)) u_eq_1420 (
        .y(_node_1280),
        .a(4'd9),
        .b(_T_1462)
    );
    wire [1:0] _node_1281;
    MUX_UNSIGNED #(.width(2)) u_mux_1421 (
        .y(_node_1281),
        .sel(_node_1280),
        .a(_T_1441_9),
        .b(_node_1279)
    );
    wire _T_1463;
    wire [31:0] _WTEMP_50;
    PAD_UNSIGNED #(.width(2), .n(32)) u_pad_1422 (
        .y(_WTEMP_50),
        .in(_node_1281)
    );
    NEQ_UNSIGNED #(.width(32)) u_neq_1423 (
        .y(_T_1463),
        .a(_c__io_read_routing_table_response_bits),
        .b(_WTEMP_50)
    );
    wire [3:0] _T_1465;
    BITS #(.width(6), .high(3), .low(0)) bits_1424 (
        .y(_T_1465),
        .in(_value_7__q)
    );
    wire _T_1467;
    EQ_UNSIGNED #(.width(1)) u_eq_1425 (
        .y(_T_1467),
        .a(reset),
        .b(1'h0)
    );
    wire _T_1469;
    BITWISEOR #(.width(1)) bitwiseor_1426 (
        .y(_T_1469),
        .a(1'h0),
        .b(reset)
    );
    wire _T_1471;
    EQ_UNSIGNED #(.width(1)) u_eq_1427 (
        .y(_T_1471),
        .a(_T_1469),
        .b(1'h0)
    );
    wire _T_1473;
    EQ_UNSIGNED #(.width(1)) u_eq_1428 (
        .y(_T_1473),
        .a(reset),
        .b(1'h0)
    );
    wire _T_1475;
    EQ_UNSIGNED #(.width(6)) u_eq_1429 (
        .y(_T_1475),
        .a(_value_7__q),
        .b(6'h20)
    );
    wire [6:0] _T_1477;
    wire [5:0] _WTEMP_51;
    PAD_UNSIGNED #(.width(1), .n(6)) u_pad_1430 (
        .y(_WTEMP_51),
        .in(1'h1)
    );
    ADD_UNSIGNED #(.width(6)) u_add_1431 (
        .y(_T_1477),
        .a(_value_7__q),
        .b(_WTEMP_51)
    );
    wire [5:0] _T_1478;
    TAIL #(.width(7), .n(1)) tail_1432 (
        .y(_T_1478),
        .in(_T_1477)
    );
    wire _T_1481;
    EQ_UNSIGNED #(.width(1)) u_eq_1433 (
        .y(_T_1481),
        .a(__T_13__q),
        .b(1'h0)
    );
    wire _T_1483;
    wire [7:0] _WTEMP_52;
    PAD_UNSIGNED #(.width(6), .n(8)) u_pad_1434 (
        .y(_WTEMP_52),
        .in(6'h20)
    );
    EQ_UNSIGNED #(.width(8)) u_eq_1435 (
        .y(_T_1483),
        .a(__T_10__q),
        .b(_WTEMP_52)
    );
    wire _node_1282;
    MUX_UNSIGNED #(.width(1)) u_mux_1436 (
        .y(_node_1282),
        .sel(_T_1284),
        .a(_node_1153),
        .b(_node_1154)
    );
    wire [8:0] _T_1486;
    wire [7:0] _WTEMP_53;
    PAD_UNSIGNED #(.width(1), .n(8)) u_pad_1437 (
        .y(_WTEMP_53),
        .in(1'h1)
    );
    ADD_UNSIGNED #(.width(8)) u_add_1438 (
        .y(_T_1486),
        .a(__T_10__q),
        .b(_WTEMP_53)
    );
    wire [7:0] _T_1487;
    TAIL #(.width(9), .n(1)) tail_1439 (
        .y(_T_1487),
        .in(_T_1486)
    );
    wire [7:0] _node_1283;
    MUX_UNSIGNED #(.width(8)) u_mux_1440 (
        .y(_node_1283),
        .sel(_T_1284),
        .a(_node_1151),
        .b(_node_1152)
    );
    wire _node_1284;
    MUX_UNSIGNED #(.width(1)) u_mux_1441 (
        .y(_node_1284),
        .sel(_T_1483),
        .a(1'h1),
        .b(_node_1282)
    );
    wire _node_1285;
    MUX_UNSIGNED #(.width(1)) u_mux_1442 (
        .y(_node_1285),
        .sel(_T_1284),
        .a(_node_1153),
        .b(_node_1154)
    );
    wire [7:0] _node_1286;
    MUX_UNSIGNED #(.width(8)) u_mux_1443 (
        .y(_node_1286),
        .sel(_T_1481),
        .a(_T_1487),
        .b(_node_1283)
    );
    wire [7:0] _node_1287;
    MUX_UNSIGNED #(.width(8)) u_mux_1444 (
        .y(_node_1287),
        .sel(_T_1284),
        .a(_node_1151),
        .b(_node_1152)
    );
    wire _node_1288;
    MUX_UNSIGNED #(.width(1)) u_mux_1445 (
        .y(_node_1288),
        .sel(_T_1481),
        .a(_node_1284),
        .b(_node_1285)
    );
    wire _node_1289;
    MUX_UNSIGNED #(.width(1)) u_mux_1446 (
        .y(_node_1289),
        .sel(_T_1284),
        .a(_node_1153),
        .b(_node_1154)
    );
    wire [5:0] _node_1290;
    wire [5:0] _WTEMP_54;
    PAD_UNSIGNED #(.width(1), .n(6)) u_pad_1447 (
        .y(_WTEMP_54),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(6)) u_mux_1448 (
        .y(_node_1290),
        .sel(_T_1475),
        .a(_WTEMP_54),
        .b(_T_1478)
    );
    wire _T_1489;
    EQ_UNSIGNED #(.width(1)) u_eq_1449 (
        .y(_T_1489),
        .a(reset),
        .b(1'h0)
    );
    MUX_UNSIGNED #(.width(8)) u_mux_1450 (
        .y(_WTEMP_6),
        .sel(_T_1456),
        .a(_node_1286),
        .b(_node_1287)
    );
    assign _T_1045_0 = 1'h0;
    assign _T_1045_1 = 1'h0;
    assign _T_1045_10 = 1'h0;
    assign _T_1045_11 = 1'h1;
    assign _T_1045_12 = 1'h0;
    assign _T_1045_13 = 1'h0;
    assign _T_1045_14 = 1'h1;
    assign _T_1045_15 = 1'h0;
    assign _T_1045_16 = 1'h0;
    assign _T_1045_17 = 1'h0;
    assign _T_1045_18 = 1'h0;
    assign _T_1045_19 = 1'h0;
    assign _T_1045_2 = 1'h0;
    assign _T_1045_20 = 1'h0;
    assign _T_1045_21 = 1'h0;
    assign _T_1045_22 = 1'h1;
    assign _T_1045_23 = 1'h0;
    assign _T_1045_24 = 1'h0;
    assign _T_1045_25 = 1'h0;
    assign _T_1045_26 = 1'h0;
    assign _T_1045_27 = 1'h1;
    assign _T_1045_28 = 1'h0;
    assign _T_1045_29 = 1'h1;
    assign _T_1045_3 = 1'h0;
    assign _T_1045_30 = 1'h0;
    assign _T_1045_31 = 1'h0;
    assign _T_1045_32 = 1'h0;
    assign _T_1045_33 = 1'h0;
    assign _T_1045_34 = 1'h0;
    assign _T_1045_35 = 1'h0;
    assign _T_1045_36 = 1'h0;
    assign _T_1045_37 = 1'h0;
    assign _T_1045_38 = 1'h0;
    assign _T_1045_39 = 1'h0;
    assign _T_1045_4 = 1'h0;
    assign _T_1045_40 = 1'h0;
    assign _T_1045_41 = 1'h0;
    assign _T_1045_42 = 1'h0;
    assign _T_1045_43 = 1'h0;
    assign _T_1045_44 = 1'h0;
    assign _T_1045_45 = 1'h0;
    assign _T_1045_46 = 1'h0;
    assign _T_1045_47 = 1'h0;
    assign _T_1045_48 = 1'h0;
    assign _T_1045_49 = 1'h0;
    assign _T_1045_5 = 1'h0;
    assign _T_1045_50 = 1'h0;
    assign _T_1045_51 = 1'h0;
    assign _T_1045_52 = 1'h0;
    assign _T_1045_6 = 1'h0;
    assign _T_1045_7 = 1'h0;
    assign _T_1045_8 = 1'h0;
    assign _T_1045_9 = 1'h0;
    PAD_UNSIGNED #(.width(3), .n(31)) u_pad_1451 (
        .y(_T_1111_0),
        .in(3'h6)
    );
    assign _T_1111_1 = 31'h70890D84;
    PAD_UNSIGNED #(.width(29), .n(31)) u_pad_1452 (
        .y(_T_1111_2),
        .in(29'h12C3D7CC)
    );
    PAD_UNSIGNED #(.width(25), .n(31)) u_pad_1453 (
        .y(_T_1111_3),
        .in(25'h12E47AF)
    );
    assign _T_1111_4 = 31'h480EBC3D;
    PAD_UNSIGNED #(.width(1), .n(31)) u_pad_1454 (
        .y(_T_1111_5),
        .in(1'h0)
    );
    assign _T_1209_0 = 1'h0;
    assign _T_1209_1 = 1'h0;
    assign _T_1209_10 = 1'h0;
    assign _T_1209_11 = 1'h0;
    assign _T_1209_12 = 1'h1;
    assign _T_1209_13 = 1'h0;
    assign _T_1209_14 = 1'h0;
    assign _T_1209_15 = 1'h1;
    assign _T_1209_16 = 1'h0;
    assign _T_1209_17 = 1'h0;
    assign _T_1209_18 = 1'h0;
    assign _T_1209_19 = 1'h0;
    assign _T_1209_2 = 1'h0;
    assign _T_1209_20 = 1'h1;
    assign _T_1209_21 = 1'h0;
    assign _T_1209_22 = 1'h0;
    assign _T_1209_23 = 1'h0;
    assign _T_1209_24 = 1'h0;
    assign _T_1209_25 = 1'h0;
    assign _T_1209_26 = 1'h0;
    assign _T_1209_27 = 1'h0;
    assign _T_1209_28 = 1'h0;
    assign _T_1209_29 = 1'h0;
    assign _T_1209_3 = 1'h0;
    assign _T_1209_30 = 1'h1;
    assign _T_1209_31 = 1'h0;
    assign _T_1209_32 = 1'h0;
    assign _T_1209_33 = 1'h0;
    assign _T_1209_34 = 1'h0;
    assign _T_1209_35 = 1'h0;
    assign _T_1209_36 = 1'h0;
    assign _T_1209_37 = 1'h0;
    assign _T_1209_38 = 1'h0;
    assign _T_1209_39 = 1'h0;
    assign _T_1209_4 = 1'h0;
    assign _T_1209_40 = 1'h0;
    assign _T_1209_41 = 1'h0;
    assign _T_1209_42 = 1'h0;
    assign _T_1209_43 = 1'h0;
    assign _T_1209_44 = 1'h0;
    assign _T_1209_45 = 1'h0;
    assign _T_1209_46 = 1'h0;
    assign _T_1209_47 = 1'h0;
    assign _T_1209_48 = 1'h0;
    assign _T_1209_49 = 1'h0;
    assign _T_1209_5 = 1'h0;
    assign _T_1209_50 = 1'h0;
    assign _T_1209_51 = 1'h0;
    assign _T_1209_52 = 1'h0;
    assign _T_1209_6 = 1'h0;
    assign _T_1209_7 = 1'h0;
    assign _T_1209_8 = 1'h0;
    assign _T_1209_9 = 1'h0;
    PAD_UNSIGNED #(.width(4), .n(29)) u_pad_1455 (
        .y(_T_1274_0),
        .in(4'h9)
    );
    PAD_UNSIGNED #(.width(26), .n(29)) u_pad_1456 (
        .y(_T_1274_1),
        .in(26'h2F45883)
    );
    assign _T_1274_2 = 29'h107FB3AC;
    PAD_UNSIGNED #(.width(28), .n(29)) u_pad_1457 (
        .y(_T_1274_3),
        .in(28'hD5FF365)
    );
    PAD_UNSIGNED #(.width(1), .n(29)) u_pad_1458 (
        .y(_T_1274_4),
        .in(1'h0)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_1459 (
        .y(_WTEMP_7),
        .sel(_T_1456),
        .a(_node_1288),
        .b(_node_1289)
    );
    assign _T_1371_0 = 1'h1;
    assign _T_1371_1 = 1'h1;
    assign _T_1371_10 = 1'h0;
    assign _T_1371_11 = 1'h0;
    assign _T_1371_12 = 1'h0;
    assign _T_1371_13 = 1'h0;
    assign _T_1371_14 = 1'h0;
    assign _T_1371_15 = 1'h0;
    assign _T_1371_16 = 1'h0;
    assign _T_1371_17 = 1'h0;
    assign _T_1371_18 = 1'h0;
    assign _T_1371_19 = 1'h0;
    assign _T_1371_2 = 1'h1;
    assign _T_1371_20 = 1'h0;
    assign _T_1371_21 = 1'h0;
    assign _T_1371_22 = 1'h0;
    assign _T_1371_23 = 1'h0;
    assign _T_1371_24 = 1'h0;
    assign _T_1371_25 = 1'h0;
    assign _T_1371_26 = 1'h0;
    assign _T_1371_27 = 1'h0;
    assign _T_1371_28 = 1'h0;
    assign _T_1371_29 = 1'h0;
    assign _T_1371_3 = 1'h1;
    assign _T_1371_30 = 1'h0;
    assign _T_1371_31 = 1'h0;
    assign _T_1371_32 = 1'h0;
    assign _T_1371_33 = 1'h0;
    assign _T_1371_34 = 1'h0;
    assign _T_1371_35 = 1'h0;
    assign _T_1371_36 = 1'h0;
    assign _T_1371_37 = 1'h0;
    assign _T_1371_38 = 1'h0;
    assign _T_1371_39 = 1'h0;
    assign _T_1371_4 = 1'h1;
    assign _T_1371_40 = 1'h0;
    assign _T_1371_41 = 1'h0;
    assign _T_1371_42 = 1'h0;
    assign _T_1371_43 = 1'h0;
    assign _T_1371_44 = 1'h0;
    assign _T_1371_45 = 1'h0;
    assign _T_1371_46 = 1'h0;
    assign _T_1371_47 = 1'h0;
    assign _T_1371_48 = 1'h0;
    assign _T_1371_49 = 1'h0;
    assign _T_1371_5 = 1'h1;
    assign _T_1371_50 = 1'h0;
    assign _T_1371_51 = 1'h0;
    assign _T_1371_52 = 1'h0;
    assign _T_1371_6 = 1'h1;
    assign _T_1371_7 = 1'h1;
    assign _T_1371_8 = 1'h1;
    assign _T_1371_9 = 1'h0;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_1460 (
        .y(_T_1441_0),
        .in(1'h0)
    );
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_1461 (
        .y(_T_1441_1),
        .in(1'h1)
    );
    assign _T_1441_2 = 2'h2;
    assign _T_1441_3 = 2'h3;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_1462 (
        .y(_T_1441_4),
        .in(1'h0)
    );
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_1463 (
        .y(_T_1441_5),
        .in(1'h0)
    );
    assign _T_1441_6 = 2'h3;
    assign _T_1441_7 = 2'h2;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_1464 (
        .y(_T_1441_8),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_1465 (
        .y(_T_1441_9),
        .in(1'h0)
    );
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_1466 (
        .y(_T_157_0),
        .in(1'h0)
    );
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_1467 (
        .y(_T_157_1),
        .in(1'h0)
    );
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_1468 (
        .y(_T_157_2),
        .in(1'h1)
    );
    assign _T_157_3 = 2'h2;
    assign _T_157_4 = 2'h3;
    assign _T_157_5 = 2'h3;
    assign _T_157_6 = 2'h2;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_1469 (
        .y(_T_157_7),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_1470 (
        .y(_T_157_8),
        .in(1'h0)
    );
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_1471 (
        .y(_T_157_9),
        .in(1'h0)
    );
    assign _WTEMP_8 = _T_24;
    assign _T_243_0 = 1'h0;
    assign _T_243_1 = 1'h0;
    assign _T_243_10 = 1'h0;
    assign _T_243_11 = 1'h0;
    assign _T_243_12 = 1'h0;
    assign _T_243_13 = 1'h1;
    assign _T_243_14 = 1'h1;
    assign _T_243_15 = 1'h1;
    assign _T_243_16 = 1'h1;
    assign _T_243_17 = 1'h0;
    assign _T_243_18 = 1'h0;
    assign _T_243_19 = 1'h0;
    assign _T_243_2 = 1'h0;
    assign _T_243_20 = 1'h0;
    assign _T_243_21 = 1'h0;
    assign _T_243_22 = 1'h0;
    assign _T_243_23 = 1'h0;
    assign _T_243_24 = 1'h0;
    assign _T_243_25 = 1'h0;
    assign _T_243_26 = 1'h0;
    assign _T_243_27 = 1'h0;
    assign _T_243_28 = 1'h0;
    assign _T_243_29 = 1'h0;
    assign _T_243_3 = 1'h0;
    assign _T_243_30 = 1'h0;
    assign _T_243_31 = 1'h0;
    assign _T_243_32 = 1'h1;
    assign _T_243_33 = 1'h1;
    assign _T_243_34 = 1'h1;
    assign _T_243_35 = 1'h1;
    assign _T_243_36 = 1'h1;
    assign _T_243_37 = 1'h1;
    assign _T_243_38 = 1'h1;
    assign _T_243_39 = 1'h1;
    assign _T_243_4 = 1'h0;
    assign _T_243_40 = 1'h1;
    assign _T_243_41 = 1'h1;
    assign _T_243_42 = 1'h1;
    assign _T_243_43 = 1'h1;
    assign _T_243_44 = 1'h1;
    assign _T_243_45 = 1'h1;
    assign _T_243_46 = 1'h1;
    assign _T_243_47 = 1'h1;
    assign _T_243_48 = 1'h1;
    assign _T_243_49 = 1'h1;
    assign _T_243_5 = 1'h0;
    assign _T_243_50 = 1'h1;
    assign _T_243_51 = 1'h1;
    assign _T_243_52 = 1'h0;
    assign _T_243_6 = 1'h0;
    assign _T_243_7 = 1'h0;
    assign _T_243_8 = 1'h0;
    assign _T_243_9 = 1'h0;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1472 (
        .y(_T_328_0),
        .in(1'h0)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1473 (
        .y(_T_328_1),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1474 (
        .y(_T_328_10),
        .in(3'h6)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1475 (
        .y(_T_328_11),
        .in(3'h7)
    );
    assign _T_328_12 = 4'h8;
    assign _T_328_13 = 4'h9;
    assign _T_328_14 = 4'hA;
    assign _T_328_15 = 4'hB;
    assign _T_328_16 = 4'hC;
    assign _T_328_17 = 4'hD;
    assign _T_328_18 = 4'hE;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1476 (
        .y(_T_328_19),
        .in(1'h0)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1477 (
        .y(_T_328_2),
        .in(2'h2)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1478 (
        .y(_T_328_20),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1479 (
        .y(_T_328_21),
        .in(2'h2)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1480 (
        .y(_T_328_22),
        .in(2'h3)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1481 (
        .y(_T_328_23),
        .in(3'h4)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1482 (
        .y(_T_328_24),
        .in(1'h0)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1483 (
        .y(_T_328_3),
        .in(2'h3)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1484 (
        .y(_T_328_4),
        .in(1'h0)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1485 (
        .y(_T_328_5),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1486 (
        .y(_T_328_6),
        .in(2'h2)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1487 (
        .y(_T_328_7),
        .in(2'h3)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1488 (
        .y(_T_328_8),
        .in(3'h4)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1489 (
        .y(_T_328_9),
        .in(3'h5)
    );
    PAD_UNSIGNED #(.width(1), .n(31)) u_pad_1490 (
        .y(_T_383_0),
        .in(1'h0)
    );
    PAD_UNSIGNED #(.width(2), .n(31)) u_pad_1491 (
        .y(_T_383_1),
        .in(2'h3)
    );
    PAD_UNSIGNED #(.width(30), .n(31)) u_pad_1492 (
        .y(_T_383_10),
        .in(30'h280E4938)
    );
    PAD_UNSIGNED #(.width(29), .n(31)) u_pad_1493 (
        .y(_T_383_11),
        .in(29'h107FB3AC)
    );
    PAD_UNSIGNED #(.width(30), .n(31)) u_pad_1494 (
        .y(_T_383_12),
        .in(30'h2F19D47B)
    );
    PAD_UNSIGNED #(.width(29), .n(31)) u_pad_1495 (
        .y(_T_383_13),
        .in(29'h12C3D7CC)
    );
    assign _T_383_14 = 31'h5A432A9C;
    PAD_UNSIGNED #(.width(26), .n(31)) u_pad_1496 (
        .y(_T_383_15),
        .in(26'h2F9778F)
    );
    PAD_UNSIGNED #(.width(22), .n(31)) u_pad_1497 (
        .y(_T_383_16),
        .in(22'h2D705A)
    );
    assign _T_383_17 = 31'h45FB9184;
    PAD_UNSIGNED #(.width(25), .n(31)) u_pad_1498 (
        .y(_T_383_18),
        .in(25'h12E47AF)
    );
    assign _T_383_19 = 31'h7B744E21;
    PAD_UNSIGNED #(.width(3), .n(31)) u_pad_1499 (
        .y(_T_383_2),
        .in(3'h6)
    );
    assign _T_383_20 = 31'h480EBC3D;
    PAD_UNSIGNED #(.width(28), .n(31)) u_pad_1500 (
        .y(_T_383_21),
        .in(28'hD5FF365)
    );
    PAD_UNSIGNED #(.width(30), .n(31)) u_pad_1501 (
        .y(_T_383_22),
        .in(30'h205E7973)
    );
    assign _T_383_23 = 31'h5004CBD2;
    PAD_UNSIGNED #(.width(1), .n(31)) u_pad_1502 (
        .y(_T_383_24),
        .in(1'h0)
    );
    PAD_UNSIGNED #(.width(4), .n(31)) u_pad_1503 (
        .y(_T_383_3),
        .in(4'h9)
    );
    assign _T_383_4 = 31'h7DCD07AC;
    assign _T_383_5 = 31'h70890D84;
    PAD_UNSIGNED #(.width(26), .n(31)) u_pad_1504 (
        .y(_T_383_6),
        .in(26'h2F45883)
    );
    assign _T_383_7 = 31'h787ADA79;
    PAD_UNSIGNED #(.width(29), .n(31)) u_pad_1505 (
        .y(_T_383_8),
        .in(29'h16866878)
    );
    PAD_UNSIGNED #(.width(30), .n(31)) u_pad_1506 (
        .y(_T_383_9),
        .in(30'h2331B107)
    );
    MUX_UNSIGNED #(.width(8)) u_mux_1507 (
        .y(_WTEMP_4),
        .sel(_T_637),
        .a(_node_640),
        .b(_node_641)
    );
    assign _T_485_0 = 1'h0;
    assign _T_485_1 = 1'h1;
    assign _T_485_10 = 1'h0;
    assign _T_485_11 = 1'h0;
    assign _T_485_12 = 1'h0;
    assign _T_485_13 = 1'h0;
    assign _T_485_14 = 1'h0;
    assign _T_485_15 = 1'h0;
    assign _T_485_16 = 1'h0;
    assign _T_485_17 = 1'h1;
    assign _T_485_18 = 1'h1;
    assign _T_485_19 = 1'h1;
    assign _T_485_2 = 1'h0;
    assign _T_485_20 = 1'h1;
    assign _T_485_21 = 1'h1;
    assign _T_485_22 = 1'h1;
    assign _T_485_23 = 1'h1;
    assign _T_485_24 = 1'h1;
    assign _T_485_25 = 1'h1;
    assign _T_485_26 = 1'h1;
    assign _T_485_27 = 1'h1;
    assign _T_485_28 = 1'h1;
    assign _T_485_29 = 1'h1;
    assign _T_485_3 = 1'h1;
    assign _T_485_30 = 1'h1;
    assign _T_485_31 = 1'h1;
    assign _T_485_32 = 1'h0;
    assign _T_485_33 = 1'h0;
    assign _T_485_34 = 1'h0;
    assign _T_485_35 = 1'h0;
    assign _T_485_36 = 1'h0;
    assign _T_485_37 = 1'h0;
    assign _T_485_38 = 1'h0;
    assign _T_485_39 = 1'h0;
    assign _T_485_4 = 1'h0;
    assign _T_485_40 = 1'h0;
    assign _T_485_41 = 1'h0;
    assign _T_485_42 = 1'h0;
    assign _T_485_43 = 1'h0;
    assign _T_485_44 = 1'h0;
    assign _T_485_45 = 1'h0;
    assign _T_485_46 = 1'h0;
    assign _T_485_47 = 1'h0;
    assign _T_485_48 = 1'h0;
    assign _T_485_49 = 1'h0;
    assign _T_485_5 = 1'h1;
    assign _T_485_50 = 1'h0;
    assign _T_485_51 = 1'h0;
    assign _T_485_52 = 1'h0;
    assign _T_485_6 = 1'h0;
    assign _T_485_7 = 1'h1;
    assign _T_485_8 = 1'h0;
    assign _T_485_9 = 1'h0;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1508 (
        .y(_T_565_0),
        .in(1'h0)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1509 (
        .y(_T_565_1),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1510 (
        .y(_T_565_10),
        .in(3'h6)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1511 (
        .y(_T_565_11),
        .in(3'h7)
    );
    assign _T_565_12 = 4'h8;
    assign _T_565_13 = 4'h9;
    assign _T_565_14 = 4'hA;
    assign _T_565_15 = 4'hB;
    assign _T_565_16 = 4'hC;
    assign _T_565_17 = 4'hD;
    assign _T_565_18 = 4'hE;
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1512 (
        .y(_T_565_19),
        .in(1'h0)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1513 (
        .y(_T_565_2),
        .in(2'h2)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1514 (
        .y(_T_565_3),
        .in(2'h3)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1515 (
        .y(_T_565_4),
        .in(1'h0)
    );
    PAD_UNSIGNED #(.width(1), .n(4)) u_pad_1516 (
        .y(_T_565_5),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1517 (
        .y(_T_565_6),
        .in(2'h2)
    );
    PAD_UNSIGNED #(.width(2), .n(4)) u_pad_1518 (
        .y(_T_565_7),
        .in(2'h3)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1519 (
        .y(_T_565_8),
        .in(3'h4)
    );
    PAD_UNSIGNED #(.width(3), .n(4)) u_pad_1520 (
        .y(_T_565_9),
        .in(3'h5)
    );
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_1521 (
        .y(_T_610_0),
        .in(1'h1)
    );
    assign _T_610_1 = 2'h2;
    assign _T_610_10 = 2'h2;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_1522 (
        .y(_T_610_11),
        .in(1'h0)
    );
    assign _T_610_12 = 2'h2;
    assign _T_610_13 = 2'h3;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_1523 (
        .y(_T_610_14),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_1524 (
        .y(_T_610_15),
        .in(1'h1)
    );
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_1525 (
        .y(_T_610_16),
        .in(1'h1)
    );
    assign _T_610_17 = 2'h2;
    assign _T_610_18 = 2'h3;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_1526 (
        .y(_T_610_19),
        .in(1'h0)
    );
    assign _T_610_2 = 2'h3;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_1527 (
        .y(_T_610_3),
        .in(1'h0)
    );
    assign _T_610_4 = 2'h2;
    assign _T_610_5 = 2'h3;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_1528 (
        .y(_T_610_6),
        .in(1'h0)
    );
    assign _T_610_7 = 2'h2;
    assign _T_610_8 = 2'h2;
    PAD_UNSIGNED #(.width(1), .n(2)) u_pad_1529 (
        .y(_T_610_9),
        .in(1'h1)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_1530 (
        .y(_WTEMP_5),
        .sel(_T_637),
        .a(_node_642),
        .b(_node_643)
    );
    assign _T_707_0 = 1'h0;
    assign _T_707_1 = 1'h0;
    assign _T_707_10 = 1'h0;
    assign _T_707_11 = 1'h0;
    assign _T_707_12 = 1'h0;
    assign _T_707_13 = 1'h0;
    assign _T_707_14 = 1'h0;
    assign _T_707_15 = 1'h0;
    assign _T_707_16 = 1'h0;
    assign _T_707_17 = 1'h0;
    assign _T_707_18 = 1'h1;
    assign _T_707_19 = 1'h0;
    assign _T_707_2 = 1'h0;
    assign _T_707_20 = 1'h0;
    assign _T_707_21 = 1'h0;
    assign _T_707_22 = 1'h0;
    assign _T_707_23 = 1'h1;
    assign _T_707_24 = 1'h1;
    assign _T_707_25 = 1'h1;
    assign _T_707_26 = 1'h0;
    assign _T_707_27 = 1'h0;
    assign _T_707_28 = 1'h0;
    assign _T_707_29 = 1'h0;
    assign _T_707_3 = 1'h0;
    assign _T_707_30 = 1'h0;
    assign _T_707_31 = 1'h0;
    assign _T_707_32 = 1'h0;
    assign _T_707_33 = 1'h0;
    assign _T_707_34 = 1'h0;
    assign _T_707_35 = 1'h0;
    assign _T_707_36 = 1'h0;
    assign _T_707_37 = 1'h0;
    assign _T_707_38 = 1'h0;
    assign _T_707_39 = 1'h0;
    assign _T_707_4 = 1'h0;
    assign _T_707_40 = 1'h0;
    assign _T_707_41 = 1'h0;
    assign _T_707_42 = 1'h0;
    assign _T_707_43 = 1'h0;
    assign _T_707_44 = 1'h0;
    assign _T_707_45 = 1'h0;
    assign _T_707_46 = 1'h0;
    assign _T_707_47 = 1'h0;
    assign _T_707_48 = 1'h0;
    assign _T_707_49 = 1'h0;
    assign _T_707_5 = 1'h0;
    assign _T_707_50 = 1'h0;
    assign _T_707_51 = 1'h0;
    assign _T_707_52 = 1'h0;
    assign _T_707_6 = 1'h0;
    assign _T_707_7 = 1'h0;
    assign _T_707_8 = 1'h0;
    assign _T_707_9 = 1'h1;
    PAD_UNSIGNED #(.width(1), .n(31)) u_pad_1531 (
        .y(_T_773_0),
        .in(1'h0)
    );
    PAD_UNSIGNED #(.width(30), .n(31)) u_pad_1532 (
        .y(_T_773_1),
        .in(30'h2331B107)
    );
    assign _T_773_2 = 31'h5A432A9C;
    PAD_UNSIGNED #(.width(26), .n(31)) u_pad_1533 (
        .y(_T_773_3),
        .in(26'h2F9778F)
    );
    PAD_UNSIGNED #(.width(22), .n(31)) u_pad_1534 (
        .y(_T_773_4),
        .in(22'h2D705A)
    );
    PAD_UNSIGNED #(.width(1), .n(31)) u_pad_1535 (
        .y(_T_773_5),
        .in(1'h0)
    );
    assign _T_87_0 = 1'h1;
    assign _T_87_1 = 1'h0;
    assign _T_87_10 = 1'h1;
    assign _T_87_11 = 1'h1;
    assign _T_87_12 = 1'h1;
    assign _T_87_13 = 1'h0;
    assign _T_87_14 = 1'h0;
    assign _T_87_15 = 1'h0;
    assign _T_87_16 = 1'h0;
    assign _T_87_17 = 1'h0;
    assign _T_87_18 = 1'h0;
    assign _T_87_19 = 1'h0;
    assign _T_87_2 = 1'h1;
    assign _T_87_20 = 1'h0;
    assign _T_87_21 = 1'h0;
    assign _T_87_22 = 1'h0;
    assign _T_87_23 = 1'h0;
    assign _T_87_24 = 1'h0;
    assign _T_87_25 = 1'h0;
    assign _T_87_26 = 1'h0;
    assign _T_87_27 = 1'h0;
    assign _T_87_28 = 1'h0;
    assign _T_87_29 = 1'h0;
    assign _T_87_3 = 1'h0;
    assign _T_87_30 = 1'h0;
    assign _T_87_31 = 1'h0;
    assign _T_87_32 = 1'h0;
    assign _T_87_33 = 1'h0;
    assign _T_87_34 = 1'h0;
    assign _T_87_35 = 1'h0;
    assign _T_87_36 = 1'h0;
    assign _T_87_37 = 1'h0;
    assign _T_87_38 = 1'h0;
    assign _T_87_39 = 1'h0;
    assign _T_87_4 = 1'h1;
    assign _T_87_40 = 1'h0;
    assign _T_87_41 = 1'h0;
    assign _T_87_42 = 1'h0;
    assign _T_87_43 = 1'h0;
    assign _T_87_44 = 1'h0;
    assign _T_87_45 = 1'h0;
    assign _T_87_46 = 1'h0;
    assign _T_87_47 = 1'h0;
    assign _T_87_48 = 1'h0;
    assign _T_87_49 = 1'h0;
    assign _T_87_5 = 1'h0;
    assign _T_87_50 = 1'h0;
    assign _T_87_51 = 1'h0;
    assign _T_87_52 = 1'h0;
    assign _T_87_6 = 1'h1;
    assign _T_87_7 = 1'h0;
    assign _T_87_8 = 1'h1;
    assign _T_87_9 = 1'h1;
    assign _T_871_0 = 1'h0;
    assign _T_871_1 = 1'h0;
    assign _T_871_10 = 1'h1;
    assign _T_871_11 = 1'h0;
    assign _T_871_12 = 1'h0;
    assign _T_871_13 = 1'h1;
    assign _T_871_14 = 1'h0;
    assign _T_871_15 = 1'h0;
    assign _T_871_16 = 1'h1;
    assign _T_871_17 = 1'h1;
    assign _T_871_18 = 1'h0;
    assign _T_871_19 = 1'h1;
    assign _T_871_2 = 1'h0;
    assign _T_871_20 = 1'h0;
    assign _T_871_21 = 1'h1;
    assign _T_871_22 = 1'h0;
    assign _T_871_23 = 1'h0;
    assign _T_871_24 = 1'h0;
    assign _T_871_25 = 1'h0;
    assign _T_871_26 = 1'h1;
    assign _T_871_27 = 1'h0;
    assign _T_871_28 = 1'h1;
    assign _T_871_29 = 1'h0;
    assign _T_871_3 = 1'h0;
    assign _T_871_30 = 1'h0;
    assign _T_871_31 = 1'h1;
    assign _T_871_32 = 1'h1;
    assign _T_871_33 = 1'h0;
    assign _T_871_34 = 1'h0;
    assign _T_871_35 = 1'h0;
    assign _T_871_36 = 1'h0;
    assign _T_871_37 = 1'h0;
    assign _T_871_38 = 1'h0;
    assign _T_871_39 = 1'h0;
    assign _T_871_4 = 1'h0;
    assign _T_871_40 = 1'h0;
    assign _T_871_41 = 1'h0;
    assign _T_871_42 = 1'h0;
    assign _T_871_43 = 1'h0;
    assign _T_871_44 = 1'h0;
    assign _T_871_45 = 1'h0;
    assign _T_871_46 = 1'h0;
    assign _T_871_47 = 1'h0;
    assign _T_871_48 = 1'h0;
    assign _T_871_49 = 1'h0;
    assign _T_871_5 = 1'h0;
    assign _T_871_50 = 1'h0;
    assign _T_871_51 = 1'h0;
    assign _T_871_52 = 1'h0;
    assign _T_871_6 = 1'h0;
    assign _T_871_7 = 1'h0;
    assign _T_871_8 = 1'h0;
    assign _T_871_9 = 1'h0;
    PAD_UNSIGNED #(.width(2), .n(31)) u_pad_1536 (
        .y(_T_942_0),
        .in(2'h3)
    );
    assign _T_942_1 = 31'h7DCD07AC;
    PAD_UNSIGNED #(.width(1), .n(31)) u_pad_1537 (
        .y(_T_942_10),
        .in(1'h0)
    );
    assign _T_942_2 = 31'h787ADA79;
    PAD_UNSIGNED #(.width(29), .n(31)) u_pad_1538 (
        .y(_T_942_3),
        .in(29'h16866878)
    );
    PAD_UNSIGNED #(.width(30), .n(31)) u_pad_1539 (
        .y(_T_942_4),
        .in(30'h280E4938)
    );
    PAD_UNSIGNED #(.width(30), .n(31)) u_pad_1540 (
        .y(_T_942_5),
        .in(30'h2F19D47B)
    );
    assign _T_942_6 = 31'h45FB9184;
    assign _T_942_7 = 31'h7B744E21;
    PAD_UNSIGNED #(.width(30), .n(31)) u_pad_1541 (
        .y(_T_942_8),
        .in(30'h205E7973)
    );
    assign _T_942_9 = 31'h5004CBD2;
    assign _c__clock = clock;
    PAD_UNSIGNED #(.width(31), .n(64)) u_pad_1542 (
        .y(_c__io_in_bits_body),
        .in(_node_334)
    );
    PAD_UNSIGNED #(.width(4), .n(8)) u_pad_1543 (
        .y(_c__io_in_bits_header),
        .in(_node_284)
    );
    assign _c__io_in_valid = _node_440;
    PAD_UNSIGNED #(.width(4), .n(32)) u_pad_1544 (
        .y(_c__io_load_routing_table_request_bits_addr),
        .in(_node_489)
    );
    PAD_UNSIGNED #(.width(2), .n(32)) u_pad_1545 (
        .y(_c__io_load_routing_table_request_bits_data),
        .in(_node_529)
    );
    assign _c__io_load_routing_table_request_valid = _node_635;
    assign _c__io_outs_0_ready = _node_1136;
    assign _c__io_outs_1_ready = _node_750;
    assign _c__io_outs_2_ready = _node_872;
    assign _c__io_outs_3_ready = _node_1009;
    PAD_UNSIGNED #(.width(2), .n(32)) u_pad_1546 (
        .y(_c__io_read_routing_table_request_bits_addr),
        .in(_node_124)
    );
    assign _c__io_read_routing_table_request_valid = _node_230;
    assign _c__io_read_routing_table_response_ready = _node_1261;
    assign _c__reset = reset;
    MUX_UNSIGNED #(.width(4)) u_mux_1547 (
        .y(_WTEMP_10),
        .sel(_T_173),
        .a(_node_234),
        .b(_value__q)
    );
    MUX_UNSIGNED #(.width(5)) u_mux_1548 (
        .y(_WTEMP_15),
        .sel(_T_415),
        .a(_node_449),
        .b(_value_1__q)
    );
    MUX_UNSIGNED #(.width(5)) u_mux_1549 (
        .y(_WTEMP_20),
        .sel(_T_637),
        .a(_node_644),
        .b(_value_2__q)
    );
    MUX_UNSIGNED #(.width(6)) u_mux_1550 (
        .y(_WTEMP_25),
        .sel(_T_784),
        .a(_node_766),
        .b(_value_3__q)
    );
    MUX_UNSIGNED #(.width(6)) u_mux_1551 (
        .y(_WTEMP_31),
        .sel(_T_958),
        .a(_node_903),
        .b(_value_4__q)
    );
    MUX_UNSIGNED #(.width(6)) u_mux_1552 (
        .y(_WTEMP_37),
        .sel(_T_1122),
        .a(_node_1030),
        .b(_value_5__q)
    );
    MUX_UNSIGNED #(.width(6)) u_mux_1553 (
        .y(_WTEMP_43),
        .sel(_T_1284),
        .a(_node_1155),
        .b(_value_6__q)
    );
    MUX_UNSIGNED #(.width(6)) u_mux_1554 (
        .y(_WTEMP_49),
        .sel(_T_1456),
        .a(_node_1290),
        .b(_value_7__q)
    );
endmodule //RouterUnitTester
module Router(
    input clock,
    input reset,
    output io_read_routing_table_request_ready,
    input io_read_routing_table_request_valid,
    input [31:0] io_read_routing_table_request_bits_addr,
    input io_read_routing_table_response_ready,
    output io_read_routing_table_response_valid,
    output [31:0] io_read_routing_table_response_bits,
    output io_load_routing_table_request_ready,
    input io_load_routing_table_request_valid,
    input [31:0] io_load_routing_table_request_bits_addr,
    input [31:0] io_load_routing_table_request_bits_data,
    output io_in_ready,
    input io_in_valid,
    input [7:0] io_in_bits_header,
    input [63:0] io_in_bits_body,
    input io_outs_0_ready,
    output io_outs_0_valid,
    output [7:0] io_outs_0_bits_header,
    output [63:0] io_outs_0_bits_body,
    input io_outs_1_ready,
    output io_outs_1_valid,
    output [7:0] io_outs_1_bits_header,
    output [63:0] io_outs_1_bits_body,
    input io_outs_2_ready,
    output io_outs_2_valid,
    output [7:0] io_outs_2_bits_header,
    output [63:0] io_outs_2_bits_body,
    input io_outs_3_ready,
    output io_outs_3_valid,
    output [7:0] io_outs_3_bits_header,
    output [63:0] io_outs_3_bits_body
);
    wire [2:0] tbl__T_74_data;
    wire tbl__T_74_clk;
    wire tbl__T_74_en;
    wire [3:0] tbl__T_74_addr;
    wire tbl__T_81_clk;
    wire tbl__T_81_en;
    wire tbl__T_81_mask;
    wire [3:0] tbl__T_81_addr;
    wire [2:0] tbl__T_81_data;
    wire [2:0] tbl__T_92_data;
    wire tbl__T_92_clk;
    wire tbl__T_92_en;
    wire [3:0] tbl__T_92_addr;
    wire [2:0] tbl__T_104_data;
    wire tbl__T_104_clk;
    wire tbl__T_104_en;
    wire [3:0] tbl__T_104_addr;
    wire [8:0] tbl_read_datas;
    wire [2:0] tbl_read_clks;
    wire [2:0] tbl_read_ens;
    wire [11:0] tbl_read_addrs;
    wire tbl_write_clks;
    wire tbl_write_ens;
    wire tbl_write_masks;
    wire [3:0] tbl_write_addrs;
    wire [2:0] tbl_write_datas;
    BITS #(.width(9), .high(2), .low(0)) bits_1 (
        .y(tbl__T_74_data),
        .in(tbl_read_datas)
    );
    BITS #(.width(9), .high(5), .low(3)) bits_2 (
        .y(tbl__T_92_data),
        .in(tbl_read_datas)
    );
    BITS #(.width(9), .high(8), .low(6)) bits_3 (
        .y(tbl__T_104_data),
        .in(tbl_read_datas)
    );
    wire [1:0] _WTEMP_0;
    CAT #(.width_a(1), .width_b(1)) cat_4 (
        .y(_WTEMP_0),
        .a(tbl__T_104_clk),
        .b(tbl__T_92_clk)
    );
    CAT #(.width_a(2), .width_b(1)) cat_5 (
        .y(tbl_read_clks),
        .a(_WTEMP_0),
        .b(tbl__T_74_clk)
    );
    wire [1:0] _WTEMP_1;
    CAT #(.width_a(1), .width_b(1)) cat_6 (
        .y(_WTEMP_1),
        .a(tbl__T_104_en),
        .b(tbl__T_92_en)
    );
    CAT #(.width_a(2), .width_b(1)) cat_7 (
        .y(tbl_read_ens),
        .a(_WTEMP_1),
        .b(tbl__T_74_en)
    );
    wire [7:0] _WTEMP_2;
    CAT #(.width_a(4), .width_b(4)) cat_8 (
        .y(_WTEMP_2),
        .a(tbl__T_104_addr),
        .b(tbl__T_92_addr)
    );
    CAT #(.width_a(8), .width_b(4)) cat_9 (
        .y(tbl_read_addrs),
        .a(_WTEMP_2),
        .b(tbl__T_74_addr)
    );
    assign tbl_write_datas = tbl__T_81_data;
    assign tbl_write_clks = tbl__T_81_clk;
    assign tbl_write_ens = tbl__T_81_en;
    assign tbl_write_addrs = tbl__T_81_addr;
    assign tbl_write_masks = tbl__T_81_mask;
    MRMWMEM #(.depth(15), .addrbits(4), .width(3), .readernum(3), .writernum(1), .isSyncRead(0)) tbl (
        .read_datas(tbl_read_datas),
        .read_clks(tbl_read_clks),
        .read_ens(tbl_read_ens),
        .read_addrs(tbl_read_addrs),
        .write_clks(tbl_write_clks),
        .write_ens(tbl_write_ens),
        .write_masks(tbl_write_masks),
        .write_addrs(tbl_write_addrs),
        .write_datas(tbl_write_datas)
    );
    wire [31:0] _T_57;
    wire [7:0] _T_61_header;
    wire [63:0] _T_61_body;
    wire [7:0] _T_64_header;
    wire [63:0] _T_64_body;
    wire [7:0] _T_67_header;
    wire [63:0] _T_67_body;
    wire [7:0] _T_70_header;
    wire [63:0] _T_70_body;
    wire _T_71;
    BITWISEAND #(.width(1)) bitwiseand_10 (
        .y(_T_71),
        .a(io_read_routing_table_request_valid),
        .b(io_read_routing_table_response_ready)
    );
    wire [3:0] _T_73;
    BITS #(.width(32), .high(3), .low(0)) bits_11 (
        .y(_T_73),
        .in(io_read_routing_table_request_bits_addr)
    );
    assign tbl__T_74_addr = _T_73;
    assign tbl__T_74_en = _T_71;
    assign tbl__T_74_clk = clock;
    wire _node_0;
    assign _node_0 = 1'h0;
    wire [31:0] _node_1;
    assign _node_1 = _T_57;
    wire _node_2;
    assign _node_2 = 1'h0;
    wire _T_77;
    EQ_UNSIGNED #(.width(1)) u_eq_12 (
        .y(_T_77),
        .a(_T_71),
        .b(1'h0)
    );
    wire _T_78;
    BITWISEAND #(.width(1)) bitwiseand_13 (
        .y(_T_78),
        .a(_T_77),
        .b(io_load_routing_table_request_valid)
    );
    wire [3:0] _T_80;
    BITS #(.width(32), .high(3), .low(0)) bits_14 (
        .y(_T_80),
        .in(io_load_routing_table_request_bits_addr)
    );
    assign tbl__T_81_addr = _T_80;
    assign tbl__T_81_en = _T_78;
    assign tbl__T_81_clk = clock;
    assign tbl__T_81_mask = 1'h1;
    wire _T_83;
    EQ_UNSIGNED #(.width(1)) u_eq_15 (
        .y(_T_83),
        .a(reset),
        .b(1'h0)
    );
    wire _node_3;
    assign _node_3 = 1'h0;
    wire _T_85;
    EQ_UNSIGNED #(.width(1)) u_eq_16 (
        .y(_T_85),
        .a(_T_71),
        .b(1'h0)
    );
    wire _T_87;
    EQ_UNSIGNED #(.width(1)) u_eq_17 (
        .y(_T_87),
        .a(io_load_routing_table_request_valid),
        .b(1'h0)
    );
    wire _T_88;
    BITWISEAND #(.width(1)) bitwiseand_18 (
        .y(_T_88),
        .a(_T_85),
        .b(_T_87)
    );
    wire _T_89;
    BITWISEAND #(.width(1)) bitwiseand_19 (
        .y(_T_89),
        .a(_T_88),
        .b(io_in_valid)
    );
    wire [4:0] _T_90;
    BITS #(.width(8), .high(4), .low(0)) bits_20 (
        .y(_T_90),
        .in(io_in_bits_header)
    );
    wire [3:0] _T_91;
    BITS #(.width(5), .high(3), .low(0)) bits_21 (
        .y(_T_91),
        .in(_T_90)
    );
    assign tbl__T_92_addr = _T_91;
    assign tbl__T_92_en = _T_89;
    assign tbl__T_92_clk = clock;
    wire [1:0] _T_96;
    BITS #(.width(3), .high(1), .low(0)) bits_22 (
        .y(_T_96),
        .in(tbl__T_92_data)
    );
    wire [1:0] _T_101;
    BITS #(.width(3), .high(1), .low(0)) bits_23 (
        .y(_T_101),
        .in(tbl__T_92_data)
    );
    wire _node_4;
    EQ_UNSIGNED #(.width(2)) u_eq_24 (
        .y(_node_4),
        .a(_T_101),
        .b(2'd0)
    );
    wire _node_5;
    assign _node_5 = 1'h0;
    wire _node_6;
    EQ_UNSIGNED #(.width(2)) u_eq_25 (
        .y(_node_6),
        .a(_T_101),
        .b(2'd1)
    );
    wire _node_7;
    assign _node_7 = 1'h0;
    wire _node_8;
    EQ_UNSIGNED #(.width(2)) u_eq_26 (
        .y(_node_8),
        .a(_T_101),
        .b(2'd2)
    );
    wire _node_9;
    assign _node_9 = 1'h0;
    wire _node_10;
    EQ_UNSIGNED #(.width(2)) u_eq_27 (
        .y(_node_10),
        .a(_T_101),
        .b(2'd3)
    );
    wire _node_11;
    assign _node_11 = 1'h0;
    wire _node_12;
    EQ_UNSIGNED #(.width(2)) u_eq_28 (
        .y(_node_12),
        .a(_T_101),
        .b(2'd0)
    );
    wire [63:0] _node_13;
    assign _node_13 = _T_61_body;
    wire _node_14;
    EQ_UNSIGNED #(.width(2)) u_eq_29 (
        .y(_node_14),
        .a(_T_101),
        .b(2'd1)
    );
    wire [63:0] _node_15;
    assign _node_15 = _T_64_body;
    wire _node_16;
    EQ_UNSIGNED #(.width(2)) u_eq_30 (
        .y(_node_16),
        .a(_T_101),
        .b(2'd2)
    );
    wire [63:0] _node_17;
    assign _node_17 = _T_67_body;
    wire _node_18;
    EQ_UNSIGNED #(.width(2)) u_eq_31 (
        .y(_node_18),
        .a(_T_101),
        .b(2'd3)
    );
    wire [63:0] _node_19;
    assign _node_19 = _T_70_body;
    wire _node_20;
    EQ_UNSIGNED #(.width(2)) u_eq_32 (
        .y(_node_20),
        .a(_T_101),
        .b(2'd0)
    );
    wire [7:0] _node_21;
    assign _node_21 = _T_61_header;
    wire _node_22;
    EQ_UNSIGNED #(.width(2)) u_eq_33 (
        .y(_node_22),
        .a(_T_101),
        .b(2'd1)
    );
    wire [7:0] _node_23;
    assign _node_23 = _T_64_header;
    wire _node_24;
    EQ_UNSIGNED #(.width(2)) u_eq_34 (
        .y(_node_24),
        .a(_T_101),
        .b(2'd2)
    );
    wire [7:0] _node_25;
    assign _node_25 = _T_67_header;
    wire _node_26;
    EQ_UNSIGNED #(.width(2)) u_eq_35 (
        .y(_node_26),
        .a(_T_101),
        .b(2'd3)
    );
    wire [7:0] _node_27;
    assign _node_27 = _T_70_header;
    wire [3:0] _T_103;
    BITS #(.width(8), .high(3), .low(0)) bits_36 (
        .y(_T_103),
        .in(io_in_bits_header)
    );
    wire _node_28;
    EQ_UNSIGNED #(.width(2)) u_eq_37 (
        .y(_node_28),
        .a(2'd0),
        .b(_T_96)
    );
    wire _node_29;
    assign _node_29 = io_outs_0_ready;
    wire _node_30;
    EQ_UNSIGNED #(.width(2)) u_eq_38 (
        .y(_node_30),
        .a(2'd1),
        .b(_T_96)
    );
    wire _node_31;
    MUX_UNSIGNED #(.width(1)) u_mux_39 (
        .y(_node_31),
        .sel(_node_30),
        .a(io_outs_1_ready),
        .b(_node_29)
    );
    wire _node_32;
    EQ_UNSIGNED #(.width(2)) u_eq_40 (
        .y(_node_32),
        .a(2'd2),
        .b(_T_96)
    );
    wire _node_33;
    MUX_UNSIGNED #(.width(1)) u_mux_41 (
        .y(_node_33),
        .sel(_node_32),
        .a(io_outs_2_ready),
        .b(_node_31)
    );
    wire _node_34;
    EQ_UNSIGNED #(.width(2)) u_eq_42 (
        .y(_node_34),
        .a(2'd3),
        .b(_T_96)
    );
    wire _node_35;
    MUX_UNSIGNED #(.width(1)) u_mux_43 (
        .y(_node_35),
        .sel(_node_34),
        .a(io_outs_3_ready),
        .b(_node_33)
    );
    wire _node_36;
    BITWISEAND #(.width(1)) bitwiseand_44 (
        .y(_node_36),
        .a(_node_35),
        .b(_T_89)
    );
    wire _node_37;
    EQ_UNSIGNED #(.width(2)) u_eq_45 (
        .y(_node_37),
        .a(2'd0),
        .b(_T_96)
    );
    wire _node_38;
    assign _node_38 = io_outs_0_ready;
    wire _node_39;
    EQ_UNSIGNED #(.width(2)) u_eq_46 (
        .y(_node_39),
        .a(2'd1),
        .b(_T_96)
    );
    wire _node_40;
    MUX_UNSIGNED #(.width(1)) u_mux_47 (
        .y(_node_40),
        .sel(_node_39),
        .a(io_outs_1_ready),
        .b(_node_38)
    );
    wire _node_41;
    EQ_UNSIGNED #(.width(2)) u_eq_48 (
        .y(_node_41),
        .a(2'd2),
        .b(_T_96)
    );
    wire _node_42;
    MUX_UNSIGNED #(.width(1)) u_mux_49 (
        .y(_node_42),
        .sel(_node_41),
        .a(io_outs_2_ready),
        .b(_node_40)
    );
    wire _node_43;
    EQ_UNSIGNED #(.width(2)) u_eq_50 (
        .y(_node_43),
        .a(2'd3),
        .b(_T_96)
    );
    wire _node_44;
    MUX_UNSIGNED #(.width(1)) u_mux_51 (
        .y(_node_44),
        .sel(_node_43),
        .a(io_outs_3_ready),
        .b(_node_42)
    );
    wire _node_45;
    BITWISEAND #(.width(1)) bitwiseand_52 (
        .y(_node_45),
        .a(_node_44),
        .b(_T_89)
    );
    assign tbl__T_104_addr = _T_103;
    assign tbl__T_104_en = _node_45;
    assign tbl__T_104_clk = clock;
    wire _T_106;
    EQ_UNSIGNED #(.width(1)) u_eq_53 (
        .y(_T_106),
        .a(reset),
        .b(1'h0)
    );
    wire _node_46;
    EQ_UNSIGNED #(.width(2)) u_eq_54 (
        .y(_node_46),
        .a(2'd0),
        .b(_T_96)
    );
    wire _node_47;
    assign _node_47 = io_outs_0_ready;
    wire _node_48;
    EQ_UNSIGNED #(.width(2)) u_eq_55 (
        .y(_node_48),
        .a(2'd1),
        .b(_T_96)
    );
    wire _node_49;
    MUX_UNSIGNED #(.width(1)) u_mux_56 (
        .y(_node_49),
        .sel(_node_48),
        .a(io_outs_1_ready),
        .b(_node_47)
    );
    wire _node_50;
    EQ_UNSIGNED #(.width(2)) u_eq_57 (
        .y(_node_50),
        .a(2'd2),
        .b(_T_96)
    );
    wire _node_51;
    MUX_UNSIGNED #(.width(1)) u_mux_58 (
        .y(_node_51),
        .sel(_node_50),
        .a(io_outs_2_ready),
        .b(_node_49)
    );
    wire _node_52;
    EQ_UNSIGNED #(.width(2)) u_eq_59 (
        .y(_node_52),
        .a(2'd3),
        .b(_T_96)
    );
    wire _node_53;
    MUX_UNSIGNED #(.width(1)) u_mux_60 (
        .y(_node_53),
        .sel(_node_52),
        .a(io_outs_3_ready),
        .b(_node_51)
    );
    wire _node_54;
    assign _node_54 = 1'h0;
    wire [63:0] _node_55;
    MUX_UNSIGNED #(.width(64)) u_mux_61 (
        .y(_node_55),
        .sel(_node_12),
        .a(io_in_bits_body),
        .b(_node_13)
    );
    wire [63:0] _node_56;
    assign _node_56 = _T_61_body;
    wire [7:0] _node_57;
    MUX_UNSIGNED #(.width(8)) u_mux_62 (
        .y(_node_57),
        .sel(_node_20),
        .a(io_in_bits_header),
        .b(_node_21)
    );
    wire [7:0] _node_58;
    assign _node_58 = _T_61_header;
    wire _node_59;
    MUX_UNSIGNED #(.width(1)) u_mux_63 (
        .y(_node_59),
        .sel(_node_4),
        .a(1'h1),
        .b(_node_5)
    );
    wire _node_60;
    assign _node_60 = 1'h0;
    wire [63:0] _node_61;
    MUX_UNSIGNED #(.width(64)) u_mux_64 (
        .y(_node_61),
        .sel(_node_14),
        .a(io_in_bits_body),
        .b(_node_15)
    );
    wire [63:0] _node_62;
    assign _node_62 = _T_64_body;
    wire [7:0] _node_63;
    MUX_UNSIGNED #(.width(8)) u_mux_65 (
        .y(_node_63),
        .sel(_node_22),
        .a(io_in_bits_header),
        .b(_node_23)
    );
    wire [7:0] _node_64;
    assign _node_64 = _T_64_header;
    wire _node_65;
    MUX_UNSIGNED #(.width(1)) u_mux_66 (
        .y(_node_65),
        .sel(_node_6),
        .a(1'h1),
        .b(_node_7)
    );
    wire _node_66;
    assign _node_66 = 1'h0;
    wire [63:0] _node_67;
    MUX_UNSIGNED #(.width(64)) u_mux_67 (
        .y(_node_67),
        .sel(_node_16),
        .a(io_in_bits_body),
        .b(_node_17)
    );
    wire [63:0] _node_68;
    assign _node_68 = _T_67_body;
    wire [7:0] _node_69;
    MUX_UNSIGNED #(.width(8)) u_mux_68 (
        .y(_node_69),
        .sel(_node_24),
        .a(io_in_bits_header),
        .b(_node_25)
    );
    wire [7:0] _node_70;
    assign _node_70 = _T_67_header;
    wire _node_71;
    MUX_UNSIGNED #(.width(1)) u_mux_69 (
        .y(_node_71),
        .sel(_node_8),
        .a(1'h1),
        .b(_node_9)
    );
    wire _node_72;
    assign _node_72 = 1'h0;
    wire [63:0] _node_73;
    MUX_UNSIGNED #(.width(64)) u_mux_70 (
        .y(_node_73),
        .sel(_node_18),
        .a(io_in_bits_body),
        .b(_node_19)
    );
    wire [63:0] _node_74;
    assign _node_74 = _T_70_body;
    wire [7:0] _node_75;
    MUX_UNSIGNED #(.width(8)) u_mux_71 (
        .y(_node_75),
        .sel(_node_26),
        .a(io_in_bits_header),
        .b(_node_27)
    );
    wire [7:0] _node_76;
    assign _node_76 = _T_70_header;
    wire _node_77;
    MUX_UNSIGNED #(.width(1)) u_mux_72 (
        .y(_node_77),
        .sel(_node_10),
        .a(1'h1),
        .b(_node_11)
    );
    wire _node_78;
    assign _node_78 = 1'h0;
    wire _node_79;
    MUX_UNSIGNED #(.width(1)) u_mux_73 (
        .y(_node_79),
        .sel(_node_53),
        .a(1'h1),
        .b(_node_54)
    );
    wire _node_80;
    assign _node_80 = 1'h0;
    wire [63:0] _node_81;
    MUX_UNSIGNED #(.width(64)) u_mux_74 (
        .y(_node_81),
        .sel(_node_53),
        .a(_node_55),
        .b(_node_56)
    );
    wire [63:0] _node_82;
    assign _node_82 = _T_61_body;
    wire [7:0] _node_83;
    MUX_UNSIGNED #(.width(8)) u_mux_75 (
        .y(_node_83),
        .sel(_node_53),
        .a(_node_57),
        .b(_node_58)
    );
    wire [7:0] _node_84;
    assign _node_84 = _T_61_header;
    wire _node_85;
    MUX_UNSIGNED #(.width(1)) u_mux_76 (
        .y(_node_85),
        .sel(_node_53),
        .a(_node_59),
        .b(_node_60)
    );
    wire _node_86;
    assign _node_86 = 1'h0;
    wire [63:0] _node_87;
    MUX_UNSIGNED #(.width(64)) u_mux_77 (
        .y(_node_87),
        .sel(_node_53),
        .a(_node_61),
        .b(_node_62)
    );
    wire [63:0] _node_88;
    assign _node_88 = _T_64_body;
    wire [7:0] _node_89;
    MUX_UNSIGNED #(.width(8)) u_mux_78 (
        .y(_node_89),
        .sel(_node_53),
        .a(_node_63),
        .b(_node_64)
    );
    wire [7:0] _node_90;
    assign _node_90 = _T_64_header;
    wire _node_91;
    MUX_UNSIGNED #(.width(1)) u_mux_79 (
        .y(_node_91),
        .sel(_node_53),
        .a(_node_65),
        .b(_node_66)
    );
    wire _node_92;
    assign _node_92 = 1'h0;
    wire [63:0] _node_93;
    MUX_UNSIGNED #(.width(64)) u_mux_80 (
        .y(_node_93),
        .sel(_node_53),
        .a(_node_67),
        .b(_node_68)
    );
    wire [63:0] _node_94;
    assign _node_94 = _T_67_body;
    wire [7:0] _node_95;
    MUX_UNSIGNED #(.width(8)) u_mux_81 (
        .y(_node_95),
        .sel(_node_53),
        .a(_node_69),
        .b(_node_70)
    );
    wire [7:0] _node_96;
    assign _node_96 = _T_67_header;
    wire _node_97;
    MUX_UNSIGNED #(.width(1)) u_mux_82 (
        .y(_node_97),
        .sel(_node_53),
        .a(_node_71),
        .b(_node_72)
    );
    wire _node_98;
    assign _node_98 = 1'h0;
    wire [63:0] _node_99;
    MUX_UNSIGNED #(.width(64)) u_mux_83 (
        .y(_node_99),
        .sel(_node_53),
        .a(_node_73),
        .b(_node_74)
    );
    wire [63:0] _node_100;
    assign _node_100 = _T_70_body;
    wire [7:0] _node_101;
    MUX_UNSIGNED #(.width(8)) u_mux_84 (
        .y(_node_101),
        .sel(_node_53),
        .a(_node_75),
        .b(_node_76)
    );
    wire [7:0] _node_102;
    assign _node_102 = _T_70_header;
    wire _node_103;
    MUX_UNSIGNED #(.width(1)) u_mux_85 (
        .y(_node_103),
        .sel(_node_53),
        .a(_node_77),
        .b(_node_78)
    );
    wire _node_104;
    assign _node_104 = 1'h0;
    MUX_UNSIGNED #(.width(1)) u_mux_86 (
        .y(io_in_ready),
        .sel(_T_89),
        .a(_node_79),
        .b(_node_80)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_87 (
        .y(io_load_routing_table_request_ready),
        .sel(_T_78),
        .a(1'h1),
        .b(_node_3)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_88 (
        .y(io_outs_0_bits_body),
        .sel(_T_89),
        .a(_node_81),
        .b(_node_82)
    );
    MUX_UNSIGNED #(.width(8)) u_mux_89 (
        .y(io_outs_0_bits_header),
        .sel(_T_89),
        .a(_node_83),
        .b(_node_84)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_90 (
        .y(io_outs_0_valid),
        .sel(_T_89),
        .a(_node_85),
        .b(_node_86)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_91 (
        .y(io_outs_1_bits_body),
        .sel(_T_89),
        .a(_node_87),
        .b(_node_88)
    );
    MUX_UNSIGNED #(.width(8)) u_mux_92 (
        .y(io_outs_1_bits_header),
        .sel(_T_89),
        .a(_node_89),
        .b(_node_90)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_93 (
        .y(io_outs_1_valid),
        .sel(_T_89),
        .a(_node_91),
        .b(_node_92)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_94 (
        .y(io_outs_2_bits_body),
        .sel(_T_89),
        .a(_node_93),
        .b(_node_94)
    );
    MUX_UNSIGNED #(.width(8)) u_mux_95 (
        .y(io_outs_2_bits_header),
        .sel(_T_89),
        .a(_node_95),
        .b(_node_96)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_96 (
        .y(io_outs_2_valid),
        .sel(_T_89),
        .a(_node_97),
        .b(_node_98)
    );
    MUX_UNSIGNED #(.width(64)) u_mux_97 (
        .y(io_outs_3_bits_body),
        .sel(_T_89),
        .a(_node_99),
        .b(_node_100)
    );
    MUX_UNSIGNED #(.width(8)) u_mux_98 (
        .y(io_outs_3_bits_header),
        .sel(_T_89),
        .a(_node_101),
        .b(_node_102)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_99 (
        .y(io_outs_3_valid),
        .sel(_T_89),
        .a(_node_103),
        .b(_node_104)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_100 (
        .y(io_read_routing_table_request_ready),
        .sel(_T_71),
        .a(1'h1),
        .b(_node_0)
    );
    wire [31:0] _WTEMP_3;
    PAD_UNSIGNED #(.width(3), .n(32)) u_pad_101 (
        .y(_WTEMP_3),
        .in(tbl__T_74_data)
    );
    MUX_UNSIGNED #(.width(32)) u_mux_102 (
        .y(io_read_routing_table_response_bits),
        .sel(_T_71),
        .a(_WTEMP_3),
        .b(_node_1)
    );
    MUX_UNSIGNED #(.width(1)) u_mux_103 (
        .y(io_read_routing_table_response_valid),
        .sel(_T_71),
        .a(1'h1),
        .b(_node_2)
    );
    BITS #(.width(32), .high(2), .low(0)) bits_104 (
        .y(tbl__T_81_data),
        .in(io_load_routing_table_request_bits_data)
    );
endmodule //Router
module BITS(y, in);
    parameter width = 4;
    parameter high = 2;
    parameter low = 0;
    output [high-low:0] y;
    input [width-1:0] in;
    assign y = in[high:low];
endmodule // BITS
module CAT(y, a, b);
    parameter width_a = 4;
    parameter width_b = 4;
    output [width_a+width_b-1:0] y;
    input [width_a-1:0] a;
    input [width_b-1:0] b;
    assign y = {a, b};
endmodule // CAT
module MRMWMEM(read_datas, read_clks, read_ens, read_addrs, write_clks, write_ens, write_masks, write_addrs, write_datas);
    parameter depth = 16;
    parameter addrbits = 4;
    parameter width = 32;
    parameter readernum = 2;
    parameter writernum = 2;
    parameter isSyncRead = 0;
    output [(width*readernum-1):0] read_datas;
    input [(1*readernum-1):0] read_clks;
    input [(1*readernum-1):0] read_ens;
    input [(addrbits*readernum-1):0] read_addrs;
    input [1*writernum-1:0] write_clks;
    input [1*writernum-1:0] write_ens;
    input [1*writernum-1:0] write_masks;
    input [(addrbits*writernum-1):0] write_addrs;
    input [(width*writernum-1):0] write_datas;
    reg [width-1:0] memcore [0:depth-1];
    wire [(addrbits*readernum-1):0] final_read_addrs;
    genvar gv_n;
    generate
        for (gv_n = 0; gv_n < readernum; gv_n = gv_n + 1) begin: get_final_raddrs
            if (isSyncRead) begin: raddr_processor
                reg [addrbits-1:0] read_addr_pipe_0;
                always @(posedge read_clks[gv_n]) begin
                    if (read_ens[gv_n]) begin
                        read_addr_pipe_0 <= read_addrs[gv_n*addrbits +: addrbits];
                    end
                end
                assign final_read_addrs[gv_n*addrbits +: addrbits] = read_addr_pipe_0;
            end else begin: raddr_processor
                assign final_read_addrs[gv_n*addrbits +: addrbits] = read_addrs[gv_n*addrbits +: addrbits];
            end
        end
    endgenerate
    genvar gv_k;
    generate
        for (gv_k = 0; gv_k < readernum; gv_k = gv_k + 1) begin: form_read_datas
            assign read_datas[gv_k*width +: width] = memcore[final_read_addrs[gv_k*addrbits +: addrbits]];
        end
    endgenerate
    integer i;
    always @(posedge write_clks[0]) begin
        for (i = 0; i < writernum; i = i + 1) begin
            if (write_ens[i] & write_masks[i]) begin
                memcore[write_addrs[i*addrbits +: addrbits]] <= write_datas[i*width +: width];
            end
        end
    end
endmodule // MRMWMEM
module BITWISEAND(y, a, b);
    parameter width = 4;
    output [width-1:0] y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a & b;
endmodule // BITWISEAND
module EQ_UNSIGNED(y, a, b);
    parameter width = 4;
    output y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a == b;
endmodule // EQ_UNSIGNED
module MUX_UNSIGNED(y, sel, a, b);
    parameter width = 4;
    output [width-1:0] y;
    input sel;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = sel ? a : b;
endmodule // MUX_UNSIGNED
module PAD_UNSIGNED(y, in);
    parameter width = 4;
    parameter n = 4;
    output [(n > width ? n : width)-1:0] y;
    input [width-1:0] in;
    assign y = (n > width) ? {{(n - width){1'b0}}, in} : in;
endmodule // PAD_UNSIGNED
module DFF_POSCLK(q, d, clk);
    parameter width = 4;
    output reg [width-1:0] q;
    input [width-1:0] d;
    input clk;
    always @(posedge clk) begin
        q <= d;
    end
endmodule // DFF_POSCLK
module ADD_UNSIGNED(y, a, b);
    parameter width = 4;
    output [width:0] y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a + b;
endmodule // ADD_UNSIGNED
module TAIL(y, in);
    parameter width = 4;
    parameter n = 2;
    output [width-n-1:0] y;
    input [width-1:0] in;
    assign y = in[width-n-1:0];
endmodule // TAIL
module GT_UNSIGNED(y, a, b);
    parameter width = 4;
    output y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a > b;
endmodule // GT_UNSIGNED
module NEQ_UNSIGNED(y, a, b);
    parameter width = 4;
    output y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a != b;
endmodule // NEQ_UNSIGNED
module BITWISEOR(y, a, b);
    parameter width = 4;
    output [width-1:0] y;
    input [width-1:0] a;
    input [width-1:0] b;
    assign y = a | b;
endmodule // BITWISEOR
