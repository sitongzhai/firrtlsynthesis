module TestMem(
    input clock,
    input reset
);
endmodule //TestMem
